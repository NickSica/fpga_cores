`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 160960)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5LViCV63n3qWjbWsRE22/y3hmn2EOYmqR9ZBIZuVn/yajH0YuWh2jJSx
LS8cTrCrJG9a0HW5H9DuXzZVlpkoEQiHLEQWceJuKOAezrBpz9XVZedASPpN4NFYbPSrByrSH/zw
BQENwQqwE+ME4OLOzZMgWgdyM+HKQB5HR3jLPQTKkLUSXDssHwJoicaFKz6E1Px4YWiEWUgGtEzh
lw8xSwVLzk+rhrO9LcgytMUfbTe+JmycUg7FU8XFssFu9wcwogHqDnJOiUDqteSHO+oYszuE421Y
HOaljtlR2TZCdTBhB0RAXk6Fo9fAFZre58ToxaJz++885n2cbFdAOi79k5I4zZbpq3S6Wp0p73f6
UxsMN27ixPgyzTZnnSQLKzUVIJMXr35Pw3PX5Xg7q9j0vnRlBWoriR0iUWLRPNuT+LsGartygSFs
fADEctDh5UPW0ePnrMUCSdLprLnPsGicBqNvnHlqqpPVmVKJ/EBTCbyL3PJB25A8Te1uImiDTRTU
tiv+PUnmrV4Iv31A/cQ3/5oYJ+YtvZdNK+O3Ik3J6AXzAC7xuYKBkAp7Ychyg7JIABgUJWfoorlk
xASKUSoxbroyX0GsZAzDBJMAWMV/LDuKf2bdOyLwwNwcQhhN/OgOD+dCAMSJe/Z466bLdR4xZtTg
9PjWNEUfKR1vLIpXGGbwPqR3IhIHWWEEMgoxam9a0Ipzzp7pdrK4lvjP0CdZlaTpgKgWkFoz7AWH
eEDEU3KQFN4B2oVOOQ77j2V0RPFmvGQOvq2IAShW3WfIpxdAgFDimQvO/gZZcOJ3/5CYYB+lqc9u
FMJqy5NpBfsL/7XotbyuFGxR6XsA+RYUZz+n7Ab7kuO63NLqyUxtEM4a9pLkoYuDjzVGWu0/E9RN
t/SrUG+bgQJMLa2HHbusv5UrmloSIXFmf5umjLFWzEJXHMBJ+xhTE97QaYIStbgLUIeed+ShCoY7
Lx3w8a0P0s47kHwRojyAM90cJ+a+Arjeqir/9I8zxurjWCptofc4l4E26yp+N/PqfgYyffrHA6CT
+h3TrBDJ7+bdJ5X9YspBxY/TqVq7eG9gMBz4xDkxS+BoiRauK5G0jd93GVDZkFcozctoW09RJqdF
r/XvDjgHN0bhFQCYdJpQeQGuAMZkWjjzN5JeDfiHmZL8FNzDmkQHPy0iYU0OBR3InVdTBhEdk4en
6IGDiw1fkRTBbIzOH1UoUzbDZfaJ3JX3wuYXUnkUXWgvs0Twa/0sSpbCG0dqZc0jzGhzqDtyDFft
qIh6Ik0k2GMbfkPtA83abb9GUqlhIr9oZ2d7uSG/o6oE3kvgDuSCh7EPZ4gMOp14s1N+EfBG0H6h
5M0FCnWdKDyakFLxyiXB11IjC3PDqVQBgbmjbN8o53C+MxlKwSvapEVcwksU9wzSDfmoG5eANFU9
oH2BmtYybs9CbbXoTUjo2Rgnns6qp2fSsKSLU3RAHIyAg41UWFTL9JoZ/UJTvFycG3/RipvqOMX1
FfUoWrYeQwatek5lng0FQneF4NWuzTSiuUhzhkUybmiHKrfSkabD2JDoCBbqL7dSjMhfcodv40X0
YHuvy7Giaz89pyuRml1HoeKZdclvZhI/Vd3ozDKEtxk4QKbtt+XtYIfU2g0cesqRGKr9Oy19Ywe0
/AnDeUY7D3oNFFjNfI59ext9OxLRC+28OCeOv+Jusi7zq5odVaugNjcWHbmJVXGhN6uCmD5E3jmn
M3H6bHRX918A1AIUicVK9ECGnGfNCwL5h9Ly4PXnCJuwx1tPwpeADsRjQg5mEPFa2EinY4Wb/nuw
jKmW4ywuV7lnNFwmtwXn4+/A5EDj1o8+ZNJ5LIcFZegoC3nNsejzB2dRzBOWpSjxuzIyCQChwZed
Lr49vKFyLnp302Z/UTWcpEMoXiCHksjheIky0vE8MSG8QVGVRbry0VCXPay0b/gHH2yMp8bZBAKw
+EGy4rtG2D9tuBdySkc/i6AuyO8EVlcu4f4OT/UQL+ILPGCd2sdlCy0xUunNDu5wLiysqSOR/M9x
ELMvYIK2TTVbq6zR4Sek95iXGmF0mjEtQq12OgIQ+oHMu8DrISOjSeuXWiI+sCmaCcsbZMxp+PmR
8G0OjfZHf3xQmKd8VlOo+ydTbZOd1mNf0zIRp++unQdTwyH0alyYJZ1TDgQFaP8Cz/5ctpKp2VZI
DDczU2AubI/PILhZr1+4n+xGxlX5/TX2aQN1g54Im+ER8xPUvoDyUpvltd3ZVj+QH9FkxWhDaMs3
skiILEpcQ8LpdrV3IIZ9u19ZiqcueQ0sroubXYmLz54bH9v50igVuq2kZLL1bWd++pEh+WA9keEJ
Z7AgUMl/aExQ8wIky7puWBHE4R47pLKZAv9LxkxtLk6ZPtsIkGgDIY8zzIBox0TeApqHp0aLJ3jB
4D08Uu+3fTIbMNVZq67UcRZiIlnd8ZhY8egf4TNZYVjjtmkrnfMXcogvzVvG3basN8Fpo1xeix9E
cLHUm/2XUpo3sG32x5tjYStqQNePgZggr0+K0eytNWx9v5yWWCUBoSns5UfX1wla4Cmh4mwsB08M
dHE8zFTPb7ebk3/jgxJlGgaRS3c04r09q2Sipvcbj27BBfjc8JiITxcNOd3vgPKi80Q6YuzUF1RP
kysf++8sD9NH+3ikZfIaIMIydj+Hp639M+t+wYdlVzwhNVxKUjdHtbXidRRDU5dgg/XSsswm/Om7
smZ86wZY/sOCVcgmrEAfb0+s+wviGbNz1mgomJHZZfCHKKBSEq67bYljS0Ddq+XH3EIvijmcUKgG
e9N7Dri6L5DPOTaPs09HtRhMUe4Qn5EouSwMWxIQRTFo6Li+YTSeb8W0P3Qk2ljWlVLCKvLkQs3r
dbp/lmT71UIzMXOJIKYBrtA9e5hRvQzeO3aRsLLjAVCQp/wLEpldyvP+kqc5NZdKzaiIKbv6HqO8
u+3mAEIMXhiTrANp8b3XGPuQ4ZXQNcaUJ2OCPtKH6tUCNUazDWpb+LcSdNyMdFCzyGqCSjoNF6ee
le0nkMKTO3PwRkCIbYMgCz8apV19QY+RDrQRDmPBKrZHmSuVlBgGH8x6ytntW6qihEQNpZUIpM2z
N/6aEcQgS8fM66Dif8s5DYfmhtYt9tnMIunxJZJ1JAfUNwihRlZ6ZLBjfT7YDwdoW3m+C5TUdCLX
9lDCbWobg6XYYGENG8HFyQY2GuwKmJv3tK6ttBtbRyYB/zi/mQ/TT2O5engYgVh1Udf8e37X4mqt
eeS2umF/6lS4/LZsc+AyO7MoDTnBQbqY/+rDsvPZlns0qDE39QMKnrG21fwBpcMSv7sYeqqyPe5Y
RxRergwS2U2dlSkax5VvDy8qOMt4aG0IXJL4LvVrfOzHp/F4tn6UbWLL3Nxv4yctkmjsavXzZFfr
yixG+tfWDxkEVvQ/cS6nyWuwvdne/M8mKpknfGrQssrB06bzsZbuGsYYlhFK5NG1P9WP2eVDwMNV
G7boFMef0SRfq3t9JOSqCvaQFZzYoNSxYFY0SoaUZvXYaSagQPkGepPU+3bJelrnrwkaotRGnBOA
QNSCfLDW3tqhVjbuvXWabPjdrFChou9bVMbwLEj7UnW4S9sc8iJ5qcDBg08JxJf4U3jLys7q3Phx
0jz2riBZnSn7rXE/pgEd2KqMYQFJFSWx1pEUStTJ9KxKIC8DO1sR/AYikdGcj3ZEkbg4eXXl3UWD
2N+6o+gwTdapBtQY3sSEbdWW9mzcFNnDNftF/ebukKsxc7RfAhcQjAxjkD5a/myoSxUm3+vjfT4r
aAo18B1jcOroUsgbRP0NeBTkI62ul2t2xoEVGS6p3jvtq/dN5tjlOssBRymw77DW7hdu73EGUb75
whJ7MnFvVRvk/aTzctFYzVxdubBhiiOFwc8gfC2N+lu8KXWJXFrVPhZ+TnI561KIznTustdfcHiz
wyknjbjpyJjA0XDR5/WD2LZQVsewKtMT4YCPeDb4W/+fPfzhFje5mA+sOo9FSmSaP1umByd3SPlr
hchtUbXcNOWbYhHA+vsYGUs0cb2E0KOf+Uy2yQ+6UY0SNloCED5vmAawNezkjJ2Rtee0x1U4Flfj
VgJf1zyAd8O0uiW98p6aD87JaNQFI5r3PO7r8WaPSmqz2/yPXEA7NCLPjthpo/F9wx+KarNi9trL
PdAbDm1EyNwGUsDxmCxmWzJaYx5g9gsEVwLkCBYESK5su6abb+mNqQECsCeKuZTvFnZueW9V44AH
ZSqvkOXmZKutnHRIePdzDwbvP4Oia4prIIJ6XT3ceq9q34fN9I8SJScvgpRLjk3uKbhJt0tCSyjI
M/nDJaBJociejM3WbJXVasRPu8jeCbQ3C8pF6KbJJ7RuMaB82jOjibiX0sGaX05Zw6O33kgGyLQF
/kIj7FXdXf5d8WpgqYaCxSNpNn1fGnkpv3Tx2qip6rOL5fNJsXZn+gHXdXNVAGbyV9xctNOt1k6+
dvxb7het3dF5I47rDMd7Hcyd3o5qdoJneeSfEqmkAffwrG4QNu8DffxnHu3lw8Am4vw1xa8m3dIY
121q2XMv9AZzaIrf1xXChmDcJZkLHiVCIEWJqLYrPWTKdHkeOR9TXOdeK+GNWdickR1SeVNBCgpt
4uRa+zEUm9cDxSyZQE8h2HzPCVqAQH7WPSoNY7rkEwdMzLMkI/b/wJd7lAEIcMEPy6NB0MaHnk7C
tKLZ4soWY0wYzw1yvbANzNlVBJKbouH0YLhr7Jjo2Q3aXSLp3Sx2kPZ9oksyhCY+GUPfkAhV7KKZ
7UmQRN1mh2lIg1H0e1TXjIljUjKj0pHeJ42JEV39UuAPd1Z5jIQRw1SaFQugcDQHapaanA4qNgQz
xaW7D3DGWFFuqMd9Du/zLBXZF5I3EAjzQAb5oMiasvjpG8sy63JZ6P32fu1JlJGWEd+5WvB+wSXV
Y/MbsqEmlYuihzraROCdz25FjmoSyBiE+tAjmk+3MGiY/BjY0LmkKWlt75S3/etpHNWI/SKe64S+
75FXqVTcoOM3lfK49KGo63IQPqnNsVvgKKJXSw7tUhY1afQlH2WCiVzYt96hsAdr9fjPGt5yOoAy
DazUyTrzd4sEb8+2ZWb6B42zlLUEEshqc8MPkdkPoXuYKGSW00xiHIErOINHpPvuyg3WOstc4ie2
0qTQm6NGOlbE30DWI6jAgeKIsVoW/uzjyeMIEtH8Alk7p18+ZR8VIW86i7xv4KjiQxanN0TwpgpU
guw9MWwmWTMXRW4yiNatuv5bD21xSE115TtxAtzxrLcsMvUaISDBOtCrXzhjOe/q9hMNYAZvVvTt
WF7rgF4jGq4qBNcRWoJTqNYrPnt/cpVMJTx0oWhutqCXlYAf4JjnMmPTwDQ9gpBuRPexhW+hf0Ih
Mj1u61KCT79roiu192iRlKlAyA5bNXPoCxJk2J9fwcGGtyWRKK3RZtslqq2f6N2/Z5wR0GOMYiSg
L+tkSNEk3e9kp5RvgidCZ8K+C+ioqHnxDDX9Rk2hTeZnNtkovzMNthmaUOKlTgHXz6L8FjAil8K6
uIfGNEWyOIUIfuf/5EoHZ/MMH99YUF94HyFlb49EIfT2LlbHcsk9mLwTYiSfKhTr483kExxOuth3
VDIpLDEbzxpQZw0uealLHhJKBiAFZ0SP8+4ZSm8p1RR6ibcD//TEo99q9fFSxcJ9wE8avu08TXcd
sfxBcuDKzy3MsFYXlFn/gGfoRU/ZhE9St7FMHZAhR8CRnQOQFRg3wlHWgzSsUtMrfZSOw+hK2966
yln89zfne3wu+zaGs6Dqgac7pdH0NIRUXlNmfhHEYwkj/4fs+IEHV1hAOK24aYAY/6dOiIuq3iuM
JBlVvCmFgpGWPmKHxP/Pvciwd7a8JhTaas6FxxmoLDAzgyDgb7gVXhaVkHGUlxv3YZq+BxtJ8ssO
/6hOLIZH0IcH0Mer0wbw9kRc5DfyAHWC1sciuZxaeGmoj4wpQenf40L+JQF5HtSO9E1dEeWm3Daz
/GiZpUrQ4ndg2WV3Q4IYonKxRiF1oESUk+GMAmtHlA+LdkUcMUeCx/ptk17HdxiIPGlU65aOdtao
U6YpHdBQeq1YBbWV/5MUZvXrGt594cNdYK3PGReQInEWkmxbEnGtLSHvnk9lIgTSA9jVHJQqXng/
pMob8OuxzAOj2qqn8KYYHOGM/OKiRO0IDbqmU9iT0AtV8OZGgsMQzBT3xChAMSlip+1WbpquCjwT
V4eYCTCcEBpyTRcnbcVNl/KRMJJ+UzvboHK4FqqvwEh1cmBdwiu24QuZ7nsGwQAKm8ipL6qQ0kSU
GWb+AkvD33FjdeaphVRs6G2Q3uiDvIA4+ljx2hqklAe+vKdGi8/PJ4QJDPTOmyywqAbAOYavmhaH
vggZlU1BMgmSgu2dSX/w1b4+r4Jjs+lEHXyYZTQKjHy74+Y5H6CwtbtToPUyATPhURIwhy5BGJwP
T4HRWwRwsW0XFnnuzOZIorjKt/GpnreMO/VdtZAhacMwi7zmwZivQBNwUl9AUZ/ZVFDF9YMmJYZa
3Po0UReM7onMZlMGS+t+FM7c+J6FcFWx0OVYdb6J3tQX4isyvXuPyNzS+wyHfJNfImMqsx9VjBYt
coP32uVIk0+RmPBufNS3vk1aoRxX1Ldm36yZVYgJZCkCCvXQg7c6sBIzioFpVaQQXDk8Oqtw8tTl
AOdK3t7ZvJ3EIuqFp0ofcse6BHX14n5ZibjyThbcTsRd/jHAFF3YB7MvO5dVCWTK1gCO2RmVAj+P
K1gMx6aQoETeyx6QVtVkEZw2JB4PYkiF8O5ZZDyXcmOQbi/TDblRjGlOchVxIs/+fndKQrerhCIB
AjYEcQRrkv6hxSMRjdpAV1zR9/gy65BHq2xMmzdhjvC1OUOS/YjExWsdWFRPHAhesUhsr6q6YPJW
I6/BasJ+1bTNXu+h94sFI64B21NvBOP5X0/4AMyssgTobJn8ok8a/8s8EkpdrPI/XYXo/Adpar2i
ZIAlqv82qU7HLMMHGQaMkDxChYnCnE7sGBzTXgmgmOBCzdW7iCq5kcPmlDXFim7o2eRiEHcd/pcV
KOiNUD0KG86r0EbZj5Af3Afd8SdZuVPkbk8tnGzmQbc0Po9Uiyf/aRkCsgoiQ5hWh4cPYcTat+6U
IoFY7+gpoyMHxqVjTCE8ruLMSp+AAf23VwLnRRmylMQ3jhC4k9+Y6iG5219EXefFdWprdoQ+bPE9
CuxEcYs2s0PmsR75oNyKs4s8SjUUaGMfvuVFfLdI3MJJEpaCqmHQhhwixI0qk0CZArDVwJOZl3yu
CiuUQXq0htRyDA0FJditnL56g3gJ49Dlpcva2W7/onF2OSYykEe6vKPy++v9i1mH1Md0VGG4hag4
0Y+RBtgFYNl4xA5ejxLKvU9xCgteuK8rtxYxsNcWkUxv+Jc7/6jIqYQ+XLT6ZwYvf0+m0wB6zBeR
UNf9WL1fdkBlQuNkpZjs3+gFE/SpMAGw/dEq8ofVHr1228cxXuxUZjjwIbYduD+4SeJBawjXg/64
OMCXf4etHeD4qro2tZ8c5aLq4sCPOAM+FfsgnLkOJQJO2aVkEydUzjQZCy3g+qF+WTbSoM0FUukL
ipShDmB52Wsmu9O098bUN86syLVsfycY/vX4lZdIqfmKfK442L/cNJlS9Ss7uWO4xyyyuT8l6XAB
GMljopIzMoRokZUJbOanJd7EDr84l91anb5gHXIbZ4yOAirMHc5l+OjhEzNLE2T16+GMCL4BQoEM
tv2drVAFQhFq8r+NdvLTakj6IsC5sP7MegMFiiLhYQB+osGTcQSawIVVlJyK6lBVfmcSzh6NlVOz
Dcd9dFSjo0yd3LIhSx0X2lTmy5Sss7lWm1giyp8uXx66/ZBXTy4ZHBkz1oWlkJWpoPXTtCEu9tez
/nFWS1KsxSS7Us/K/RfZh01b802p8N/091nx7if0OMEBBj1iJSTqt87LNGBaKpYvd7JkAy3fgH9H
QZYg0w2V/CHuuJSZjeohb41fpxFzaUH2E2PzOUqwg6sF1bJ5OQkCfMT+mwQYNp7M99OvQ0YDkWC8
sjEQElu3kazBYIW2G568/qiS0HN6NPI8TSOzVNlXuhGnVXvmLvAzpEEpJuib0oVhc/jlO99aEFC4
At5qsWTqpdnxftOnRVSX3/0nLbFv91+gKASEJ4ruzT1moouzuQq8xclbX/6ITAqSMb1NWyNzUDna
wo5Gvam3ObGWPmk9V/mcjpq1j0WJSTCWFu9+VGK3Mgyk2FkZOPJYDxQdlTi5okEhO+54dI+7hSVR
QxBeUcZQbmSLbCKAdOuI+16tq5I+7O14kuyjc9BxjiICQjnpfj1k5SJJWZ2LbC3HftI7NooJ4RLi
txlm+rlypmf9Sf1dJ1RR8lm3S9kXc/H2PDKFVYGc/d9HxJgydBIffR3lwgMCrok8hHfaUWiC8azy
YxTT8DkIGDC2EW+cLfppon0Ztf9anMwOYm7ntTHjOJDaXg+KRr8ikSsUVd90cpn5dfXzGJu8TE0L
jSMFNgtOWKkYOEdTVlPjga7vjA876hQOLLrWSEPvi8d2rYJ1DmXYssrk9b9yTx4lVxHSlwrJzoV/
PUqqM/mBFuYN7RRZ4vLPC0JjSALpqX2YQCHMlUvbL+pcSVy4XnyMy/eWCho1ile9IvEUFp9fKSUo
+sXSSGWwDRL2FqfoNGBBGVf8g/vPWY/tOOdHZYwhRF+HD+9EKehek4kB3mTLgyS4h28MMCDJaPFS
CpStx1hs2/dPcFpUafCMZzfUbGJymf4v8LqA1lcc9ZIAqCgy1euTVVshOysUgN4pzIN153OiTbcM
BssdJwqSoZb557yUAhBfO27urJAJiayhKYa8wY6fTEXB/HWs1vOq7XoXTxQwPK0QWvgNi1Oilkw5
YkECByUAjZtB8oJRRnrBgydzLHrFbOQTXXoeJnd5HkBN+WPlWRsl+yrI3Ibyw7ZiYKNZAmPdvX15
XxoKNrcb2gvm1e3XKToms6xR5WOkCXk2f68xq+CVGnJzAw9s29DxkH6SVFFUHWDFX/pOcTxjtlji
OpPkvjFWaV2lFbFBwkQRqdjdM2iWsXDz54pzWzMA6oFN3UFRuFVFUv8HA8qdlB/nwXqY+PpmhnP2
wEAB+kSuLXnx05W0KysW15wGnY4UR38MV9hz1KGvjVoFPoUihTSkSQTCXLQwhiB/OOausD0C9KU9
AdzwBwGXAjWuVZUVROEAvvfX9kSm+ox5t1dmGXJPYjDkmR48tgNmynx7RZSK0HifaR7xuOF2EY7J
x39gJq5p1Sdwu+nsLiiCIbrhjQaySz5vnfkW1QKvbH0XOafpGo3vRdk5bHbJbKa2MNIR/zqVP1kE
5qTZf6R6ud1Nklw3tsIL8g8WS/BKPGxTtZyHpzG1TVBGTSjdHAHy30kgLdFy6ZKgvXxfqvL0bsLR
WJxrzN0HKYFWzeWZDV+xeRDTjRGKRCWe6VwuZB6FHzDiTPYksPEO91gU/5cu8R+S9qrvO8PcD+2y
Tws2haLtpnFswf5zPQ2OMzbMEuD9lZQijT6gabTR8Yv/ZWvY7PrMYKnFopYQylvO2utJNHHZwbzm
l6UZqhbUDqDO8s0Wk4aLZFVHMrauUsKuQS2S5lx26P0SJgJFNW6uMMBikusC+ysl5AE0SfQZI4bL
TneLBSQCYpnaoEnTlh+EMAN/4r2/eOOoeeXUcZWQ1SIL0KRM2wxA6R28uT2oW45cIG34ZjZrkJF9
g0gLGxq5+8NWe7i/KR8nNoPFwlfVuWyCedrPXSIHNkiy1w+wgvSarIii31sRejhv/xHzeeLItQO5
7DYSeuTIntdfb2LNy/tKlZPOADKo+MBYMjBB7D+6d3wiFwpn09/EbTyHCxYmWCfa0Gao5UDFNxLW
eWYab2iNvflYVrwkISLrF1aATcgLkdPPDXqcCvk9OtwsD4w3baIayEvl62Ru8Wy7TGyBS4oHnHOJ
qxZSGkgvVSew9717/ly4dWBcyxKmZ1Gr2k8Sl6ZHyzwAQ2DlNQLI39fvBP4Otf5Dj+pWE7kbjcTh
5YhbHshG1D4AFDb9Wx9KIj6UJSQ/zdPjuOPt9bULGEzIbwoN+BYheuqXqZlG5FsiWLET8CFuyuLF
9pD2RrR0WCQH4Ojg5aOG+MLaxv4RShGHI1IMdsNwu6cfQ505aubmPRu2Jv6W9Ud2Ev8NfbamFEFd
yvpduC+VAaRoa4Wi9UpT8Gkp9hwD/7b7bFwZOFMYnWgu5Se7T0wS9C96ODrKygM4Sq7qBmQJETFg
tG2FZs/amK0sxAjXWDmhBztdF1tmNcCwxOud9aVXLFXTLw91a6lBY7rT0g8JkMpdUfoHNrbFGWWd
TysvBb33cwIIN+ICmq9xkPYltfiuO/FC9Des4LL3hk0ELH+tgZR0GtvcU6Q/H8vSk08PhLm9KoGo
EfKzAE4AtDPG8DLgrJwup82F0jOLPdU4DpOMmqTXTOZ9ceWRQ3q+DlEo2NgF8C0wtJL0h+nRyJps
P8fjQQ0h59EkX0cKpVqamjUzYchHAiz1R7J4oxA1AOFWwcau6qwCJ+7PnrnRkgXU8dixYBerE/+x
sieRnw8nbrxAWGSLx+5C3ptSckH/6tvPZBxZyICssQUSrWmyVEKiuqnfUR0FfzlQ9mFHLw4O9yqB
Xm0vc6hTD9eBRMCOP/zOHnQGpAC/iz+V716kdmhB+nIuDL2KFFC8hWVgA2f7ZC+3GUZ6VYobX1/1
0BGLB0LzQuntY8w0rTScwHFOqs9KBQ7u7SXS78ym/gva8n/AJ3K1SmS5b1NtEzFtfXpDpAQJNhkY
gi5kAm1fB27+JMO8dFYt80vVQRjkuGsnNNjKtTOxlU3SNYYPyB+02SCYEdhgUt9SLdfolO57NENz
bnWKKIL9TsJyFtVdu1DHzuuSCd62D8EgsCnPZxB/HL+g260251F3hiR8jwmUDjLC0BrHV1AfCZE0
8byBEiDWdWFlnrT0YXJv6HkPd5vSnEKfS4wB1mjBh9rYsdO+j7U5pVCPXAZ7Wy1yE5bb8FKmOpC/
yO1qTEorfh6Yf6f1W1YAmQsqm1OO6KXXFVTik1bpGh+nrm/FSr9K7zmpaUS6jOrDGzS3WugGfYzC
D5jxD/YkUO2O8q5YQKHXflHYhoaL+CVAS6g+Zq+TdvMzYkw4BnkUwrWqfmFwgsobnNby3uXWp3Ga
GzDw6LUuyLQNDf5c/7l1o0Fm3J6m3QxmitZ/J3hq/PT1OaJ/CUzpe6PRC9oDGG7ba3WHeg9bNaMG
kSQFaKIPoxze4F8R7aUNtWtJ3kQ+ydqQT42Ipa6giBbzmEv5PfcCsdT3t9uC6VlDQQuhtVkjZ4/3
qNEKezosertxXwNMaYKl1mAxC0n3Ze2qaCxv3zvHT9zqMYhrPPqOgwwUsnE9rqpzfitM5aVQ+1Ig
fkn/cDHQXqT5LGuYiu/Pq4Y8Rr1XNtMZ0Eo76lIT+4Lv1CYHekFqu3Lm748Lrd8qGXAWmPenzPQr
iwHop9w5C0bMQYIk81o8qz3BRp4O5XkXBH9psDQrzdi5K7xmx7h6UjX1zoXFL6NVEwTg0G7wZyHN
WlZvKhTXUIOt3PBIixjw1wmSHg7c6oPaN2qP7xxljaDlOAepCGKqbJ9qIEbtFeHyuOv+4ZRxyNFF
ksRBPmBdjwVdUBqdHgBRnxEt0hVCEl5TarjI604sEMY2KrmmVVu8sZzWIAr08VtbSb2gsJtxYJC/
hDUBfLR/8sIDT/AyHm/1p3VejNKPZ9E5wbX3gbew+iHZrQJeHNWnyExCDOT/jBHcCj+AapEdYYSf
cfdL/0486KPBTF8D0WXrEoiUiNAe0sDqpO7r2jYFPsG77bZoCbV0J46mcEsQG4ny9CwoJ2sTv3SI
WeYo5qlC/djlHNcDahBCQxeOpADcGXtFbA7tjwYjV2b+kxJeTB6fcYrZubEuGTJNrXksHQt2oiZI
WelJENRP9RFGRMevxWhgKeu3nWyKs2SxWOh3wNmPvPm8Mx141Q5SAUfQhAKqtBFrj7mVbIdPPE2D
FTWUpQ/3yZHxxnsd2cy+wWKNn3QL9/n7ZD0yFF2yHrnecGbLfEywm0QsmaOh/ZCJW+UoJSXKW/+N
sBmQmlBxDzY4CCGPsX8wOgH2a5bSTZhYhC5rc/M+Z02DjwvF3C2L4f4U5X/BKX9Y7qVxN9jUKOBi
KR52UsPdZ2bqQNEcUviObiNbyy03EAxAt3v6zmmKv/mqQuD57VSFKn7G5zoDh5honqpV+3KN/465
Bg0pd0lrnoFEniFnadqVA+TSFIjIslxeu3s2/KsDYMCu2vqjJR/JtAvxSuk7/dR/nH8lD6EbnBhB
xkd7lQ6BzxST6KEnXtvAu18M9NP5hyhNZUd1OyIgblcn0btoUnX0q/0c9zLc9K2cTFYJ85iaPaZK
9kvIi+U63mTaeOcLTfN0xCOSmUG2vI8D7/frc7tdKvR/26+YKWpeVsquJZKQkn8ZEW5Q6w4Mwaja
1bscRfR1YD/wKOGgx6RtQ6B36rfFEzaAvkDl5tzHvmYEme4/TmfEe99QTspkh7m6rHg91yqmDmZZ
3MEGUrpio1HAWOFoHlsH+M04Qyqffyho8QBEBFeBTPs8kMxi5YIZfn7qEKedyBXwQzbxinIGfE6Z
Yp8CK0KZaJKGpi81URONQ5+mlabRdDv7vUVgQ6Gqdz0sWrC9NZOdxKNoD0zo0qa6yVgTZKw1Chj0
OPmPmB0/G9Ub0tRlrTurM42fCckzyi/MWrWtBoekZsmexNMetoBCEOAl58dvvzpXKm0aFYGlj383
3/r2bpdsEIxouDS300H2tNK+wKmZHOxgzfMOjgv2KHvUNg1htWbiSAGKlKc7BOrS80/0npuRrJVS
2gL5lTvZkqueoF/moigC2jDJFmID1/tNZQh9nVkpFMpGgIy1U16ke0Zw3XMVh3cNoIXv7fPBofLs
SJoopwKkTrtDnP+YmZ1o8FG0JFi5xI4OlMs4O8YALxGKyUttDD3Jm9k8CpYhfAPrOyD+sn9PK5ng
xGciuBsxUohemjKqvRLWk+wWewAEqsBmzS5Uk3tU79xi3isnFzuyl6hx+ho0H31+GD5rbOJby0K/
sOjkokSnqGZXfMSBhzM8vr8oYD34aDW1TQeegVxHm+Bo4g7rGNW9oPE1KEo6kog4XJ8aoLYlJfoD
0Ek8/CZ6mNrdT2VSzj7Dv6K70BAJXct6z96MEUm1hhiZDmMl/zvs67rpLu6TxcICyl04TDwg2QgT
NWlp6zmzNWg1Q6HpngFKrTKkt2VX+Hnj8604J7LTLWEjyz+rKyjZSfKVkUokFR7KUJQCRN3OR4Rr
L+pcB0qDIsjiNAISd2BT52YHF8a3v98pMMlsJkHKwqbwHzDqxENmT4/IMY5y8JfigKV9c03uV4/s
aSkbYikeaBkryDfakpr3jQtbu0KamPWSpDezDr10Zo4Mw+2rDsbrCqLg9HntZI5jeUFluuJ9tUDg
sinyEIwcfS8D6fKjA5NlqyW30AZNe9gAQAOpjKQQAzCqXoPdi763wrecq4bXpHPUmVlcSk6dvHgu
XN3EbSQcdDBp0BgpE1xJblRQxVHGwvABGujWOa6p9degGfSNdCrJxDsEGvAl1y4kqCjKcPMUDsVG
geMyNF0x0PH24Ufcu8v/FHA7jkKVW2+kZdq8zJnk1xgwAYO2t+OcdJmdralitmcPe00CCbiTg/Cz
j5u3IOwqgxN5EcK6m8hsUYmZ38ECF27oVIoOMZvhVIjMh1MJ0Uv6tas04miGojHJdib4kuNeX3Hj
mULec5PR0JEYsvYGxWOx6tQkz9xzwpYIrzkimMTyKLdUknO2Gzfnzdg7gPriW5cMtgM+4iEDr9l/
htDggc7mhhP2gtrmAD1g/NSwwg7JhEnImKkzmFt04hAeYPkHbTBPRr8/6I7HggfcpxxrFFfEXc0Z
ESOK+t73P3AW96yRAsfozLGQTCqBAf9o99zJzGaCwb2Y5iBStgDD5fkGEKc4UZj6e8H2GAJVylh7
3T9v6BMi/1M1t+XlX7Kjp74gO0rD2fAofLdlPl1U+ti5V++Ha4lTa9z7qT7i7t7nqYV3FWgHRfjV
GADy3qxNQyKKEOJGXJd4vlkuPFGOFRjlCt1/UsHp/N0FehVCRNM4vYj67KKXFE1fggZL8TGNETUy
lD+8G1S9BwIkgP6PHWSbSLdIYXvYwrJ6TURPP+FQeuJcqFrgY5LeIi1S7vybYRuCWxLV3pWfn9cs
QOS4n+vnHPs/SKCR/L2guSthYqPIA1pOTMRASmouxu+9WzG4KjOoSsQHQLKQDpFPociCDHS3X7Kc
WQEB8+E/VEvANsgeYeS6zBTjXjhErJ5iEX0ZP+DAqG+bZkHXA0ZFSs0fXqDrvoMoPCgGVAAfWiw9
kHVHWNpNaLIjN5hCdikFVjs5grUqGXdOAJ1uBGceKVatlD684C1wBHsW4MICVPP0SAr2+jggu1pw
dCXIbkQ8G7NqcCTUCC1YFFegA9I8qkrInq0l0L0GpO5P4/38/DMJPki2hm5tZXRAnUCSETAY5+Fh
LYWCLYFDj459LTYUVIYmMRNUOgKRpC0fOrc+hyR4HuEN1YrZJqkT1kbV96UEx5MNwJohjaXms2fs
FeM77uxprbP2uZDCy1+Zx/AgE6fsJVAdJ+BUCqZyT6YK1/6dU+dT+q9H/298tleVNP7IESfIeDFc
ajWjwShn6mRi9IXuLXR92dd+EWeH36tYoZMaa4hrw7ssVge6Z2ETzrg5xj5bK3LI0SuyMQkSTEJC
gZBCY1Awmz0CysSdqQVDTxjpLl+WcZBn0ZrDo18FYw4hdpmcYX8/3CkYzxjKo8aD+hPz9lNRtxO7
CFwKDHBzj09HWbcJ0PUZ96Uswd5L4ShGBpukqivxPViaPXYD/yKhWIPXnC6y/RTb8aSQ+Zqbde+N
jFC1J/Nd/qc5otb7l6ecJhI1tKqdPMRC7kCrRA7wCt/UXlJshsvLZ3OFTWj+gqt/C7cAUBEJ5bf7
SSfUUrW00oZQOq8RT9UqOaklfy3hsx2jcwofNSluCekIBHEIXiDfRldEFCKUzADM4G6dfGb6OrPh
JhTn3KiSTFnVbqun6BpujiLfPfxDx0K8dBnAFXFL1p+diWLjcUdp39WufGiRsbnBhmUqTLMcSmjZ
7QkBVExXK8bV6cmOxyaAfWlOvTASsjNN4gJOUOmnkR2xngmacKExDBv+Z2oaSS45bmRLf81mqrXa
OoemGr2yvAxEKKOHCoHZpWqKiVI4VH5RNqU02OO2huxDJgcVi8sf/nyx8sNcqUoPh/XNRT2WnGkk
zNQiFZrHzNDbXBWZnjESSoPDvwHzoapD/YMa7K+hMI443O4ESbyBylN1h2EcfrzN6cH7o4g/ubFR
qQme9mAK/cF/epzdxRnjPQZ8ffj74NwfBPewUAgpTM3mf3GLgXb6XxvmAVtzs/iKJzWQH8V/QJly
uqp33sYEX0uESq1jIRzZ7wBMy4msVGVqsn0AMWvnL8wjr3AvMA/8dE1xXmjbOiicjvXIIUv0jguq
dYgoPn+1XcKewKJmlW3ql+Q59RXich3Q+x7/SjQybfsWyFHS9Uw/vXB+pCZHPMe844uDxwg5mn9I
Zms9hqZM4/CPtwI069mdIPRQsVjmCfWtG7aNYD2SMynAyfJSSGbNS+1I0MwRaRZqN4QXvYx1s5UY
lI/yWuyLEvry/G1Muye046hUYmUg22litavMeKZTTebBtV66RYatalvepxXYY9DX+2b2MICuZs2g
yuO2T17TsTGIYtPrEauqJ8ThBk1UogdDL+x5PPp1yGi9A3h+dchXYU9PbQ3kpqrtT42iCCRg22QQ
B9QIYHaq1NOawOyhMaH4qqQbmkI1R08FYJNnEIv7d2IS6374q1TanSOoxzPrBkblBgY2zDoCUWh8
akZZ7ecwtLImV1GL1gfZKu3QVm2pLdoIogqVP1qhxiF01XAKl6wWW1E5lKng+hYOvGG20Qgt3UmG
fo3gtVmhLxuSHTZWIZR/HlkZYy0L6iytMbAbqU7B/nbs7E+4/GIxDit66SwRTrbR9H6WQcVaFOrF
qqmww3EVGadCr7d9ODUSF3PBWZOyFzryOkmx4ZgN85SORZhAA3e4z2tG1hGRIJJWnmneiNgpBJG5
0WVb4Pa94nxjFrWyVivTNOHRsuc82CLb+vgdjplh32E/bEYXFelynjmwQDUABLn/JXTMqJKD7V6M
zxgukxGVdM7iMWYR4NxwxIDmoyO7j1dlggtxg27EcHhgCvFabkV4wExYbYfyDXM3r6OhJL+OtJ4R
g8HcfLIzrip9h/k4NsEKAZ5FwOyiG5yazy+5SsH7keLOloxXU16vdDv6lcUWe88AFl9Db3MsgJRK
kTP1o+pj08RXTdZ/Or1Rovso1dEJbXx7RwfNZLNb8jifOwcidGC7w+/JCQZ7Dhik53ExF5RKtomO
zQF5IbqyUPiFObxffhLi6SR+C4XVkWLgWa/PgNJOg+cVC/sh+fd8deRGIcqDEPpVXrR2sOV1st7r
H6kfC5CuudqY0cJkqKETxXVZX3RJt9gp7zInDD4Eje/7dZSwWdQJ8MfwbQ6iDVtcMJDVFEAZHlNZ
pSQVwkutzl1RIKQOEA4CRSWH9DSlDUkW+IvNkZnicz55BA6qbxKa2yW3IRGw4ZINLSgr2Vg7Wlco
S8QL83gJoQFXNVBdrwdtjGTYMyvOvBbVyDUEgPcF4/ikzWYVNdg4bOI5gMRL5FzjfRa0tGX3ltI5
DP5c4tfuDJjOZ/CBCEmnngmk3um5K1o0Bj7UWwWpTT5xnpb9yZ+Wo60h3NiuHBSjVQuA+PoU2BdB
sEg/D/ugS8CyvpZ0UUI1cZFAGGqIBpfkx9j/muji6jlDidhCjQTBTt0WtB5+2MmoRzRpLYpBnGQo
6kb7zMGY/IUZMMx0QUU3J8oGBBtTGfxy0H08HrPzPi4dQlwvcJ2gyHveGUunZ+Ta9+INK3Yf6XjC
HdhZGgmwkR1+itgKjNWbe+S54cD296T/pnbo5RYDuuQF8IkoSApN892Z+FwI4sS1XNxvCfi1BQP5
kZiF8HMBJZ/Q0FmZl+oTOXQACDt6AMND2Y3BQgMOeWRCqE5pKUuJpoDIa3hjm+v1Y8NrgGoZxa97
NcqyzhqTYAfc7Lef9yDDpvBl5k3a+ULDnkWBDUDmJC0hnu85r+go1btz8PAeOc2LYBd/zdYXsJsU
YyVgzkKjE9I1MT8ugsEpNmHhuYSMKEZghj0fhezbQwOsnMCNYfi2o/6fPiVAsPyVrSpqnU8wzlVZ
onlkX9HrWchAJIm04gZRmlJul1VGq6777kELUmDEu8vH7uo5a8NluRo/Ni1pOTk9kShPjjFQ5txK
Be28m/URwv9p+lUlGGkTJ//WE7njGK56Roi9gNbzveG8DhXSqRnWIcmK2uNp0yn5KZQmRdPN1GNp
nwRqcafgHedVMEpGqh8vG63VdVhcH5QlBa9DJdRcaZmRCkyAvSz6hnvpuVyreWCWgLb7ugDVjFdx
+HwkC/QOJmLUHKwxRY2rE2mdQtU3BkGXwKtPmOSK9ra6W/Z/lPviYrf5pczSZnZQRDJ7etIEyGKH
kfcvn3eluwpZDNuSTS03Ve5dwKHk3dGsne+4Y5sBFzFbl8oSIqfN5NNqTh1W+kAt5I975KKD4i7C
WFYKUKqsHoyt9KoqUv/DEipADAJklPybI176n0shZX6Rlx5F4oeqIdItfetqjwCeSwExE+YEWg0b
HVaM3lz1g97vQ9rso+OmnN1jSo5fN5Clmtkr/r6B3QzYK/jug+a+hs2w/I0PS8cW753QC01Jbvv4
U+5IQsBuzb8aGiJGCwwoqrV1SfuqE3v3VTHwYq8vuZPYzKWp+mQyni9dlc0foZ5jf602Jy77ouO+
E2iqHigNmI+nbyEh4eFjAVzYAB7aXhAhHhg0TO1KwtckPnbqrBtOhGuzIRra2QTdIevWCQHjbBh+
I0p3zHO/jIHZFL20BCtjxPEVrEtGacOwjcdMpqNkD2ffwMGTTUfXtfvksKi6ENH6ZhFOqU10EAlf
CQSbdCUDoWISqdwgBZmoj+Rf6gZVj9neYmRVoX6+daMQ73V6JgcienvpunWvUMw/b4wabyCXchTR
AyGi9GH5TwkUjwJpABS0UuXuQ2P8lKtgHcOd0U4lVFD9ovdnct8dJbBpBwi5VkkdPfiCTFXcxZ4w
ylFbH69EkikEys0wCfEhLDLtDIZqh0usg5LAqwRmMExzdj390ylLGae7TyVuC3RfMMHUHLnb4+Xj
4oWEaPCZHWXtOY7vpMV4918BztNCIpdgLxbkfEkKFVjk8pIzysxN3W9bkLLPN11r0CTS/kCm6oWB
NNv02BOs7OMKIBqQXlxdIur0nYqkleNWIGTBs5pOAvR/qEDj+1iBSuuF3saqMc6MOm3uDhvKCb/N
jWHNUVI+WoJAT97eUJTy768LaVqWIBOsKIbb3x6fybwbm6gUdiKVhAFhjRWy29j4/qSiLIk0gxJM
IMnm00l6+hwVCaR5bC8NvZR65ZbscygoUIm3vLjNhsgXsmAib9QRE0ZmOMTOw3YO2SUx15OoYj2z
CUcxtGyPw23ygnVSJMWc6hNRzGKWgY/zczhaKjzlzjI6icentN+b1HKPNWNkAY7wbXTeNabyOncI
bKxecOmyzwn+8j/nrapd0sIjpxXUE4nJe13ujB4OrNuJXJ3YK5XY1GCY7nU7L2983wPRUPbCkv2w
0mZ/EATPqQcqDTZ1JUTftTVqzxcKB5HQscqegLop4lvKS09iDfzzpFOI3FqCiHelpFgsiwi4+BQT
0Hq+/g4M7KczypKnZx5Ir6+0NX5v3DAlGyXMFZV2vKcuoXc/q2zyTl4ElIflwaPHfBk6fobmUb9i
4wiPbJdYHZURH1DN/YKBcclU5a/7eHyMaA9I3+SPNbd+Hk2DNLxwlu1qsNw+/Fe1qkC8W5BmtNQf
6hlxVZfKEpvoGyRpJwA/95vhrDyUdqXKLGMcrBk6VTu+BgsNVhTMxGavEqih1A/hMp8bXqEdyKY0
HGnnHogcg3UhrfaPh/oMjsWr8CERgj2PCkKGtfGXly123B74UkxBxpZGwpw9gJEy3sKXR/WsYfdZ
PckquqYxy5CyskYVlqoqpoBYUtljPirDmC1y1Gt+rayc51fRtGG8s+EysZDIkII4xZ+ODePmDPgw
HcqjJA2oGEhBPMrr7EMbR4rl/YO9HxW+360YFyD8ULTRvQ8Lv15wmqha6U/KEYMddGEM2a73eokp
xniF/K6L+1eEF4x4u3lx0eaPOHRpxPRTcHp7aGYeOsYmQTdWpXN0J2KdnHbJTAHDyLau11NEdMXc
8tkqRt8gIkM6vR9Rwf9NX124YC02nLm3TRT0cEQS8MfnJuyN8yKrW5zX9AzMG0kylWNT2/q7m47p
I3BZlG4DqhZYG1ti5bbmUmhRos8cT0GSlaYVuwwhTyOm7y+B74qVoTWaIeGCyAzSQDGfuht+lUzn
kF1RQ5o7LZKCqDM5XOaKQs8gErYPNPWNUlzLBwCWPTMCFwAu+WCZM5/MSPe5oLRd1OyfTX2b8pGJ
MjelDFA8sK62srX6SkcjxLn7ZfghwVGVNPnxuwf8ph8eD+FdLcoRVyjfn9FcTKh3oukwQoKUpFvG
7GGOllw9gT2E6gfCZ+OD8o4ZYZNPJlFiooml7cw+Lbj4evvBfBNoA8jCJZ0+2lJvUU6rB7DinXTe
lL0hUc76uLoHeVKmzovWDI9xIXFihpzTCUxUf6JB7p8S7xMgYSw9kHnH2D8cYBpUB027wJuFQ6cK
OLagETOgG1kIJl5Koc2KxAICa6qpY0YPkI8V62YrTfSqheq3P1J09I+P/QmhaMh6APU7ARRezyax
OFcI05VGefu8qQBsd+iwnsgFFyXm0fgwafmfMQ2LEerau7SlAMA1vTmP7wgSk87n/Q4rcL+fCFzZ
N11HYjt8a/grqxiJXUeyAShhfs0kujmP0q2wodooJqhK2YYkbekzZVui+03pBw19LeYug514EtcS
4253k+lGnbyU2+KJF+IKKVcIQjwErkxAewKqPTzRot6/M1eOcRgHtpD+h2hbovjDM3TfNSYzKyFp
SmMCkizMA2c2HagpOzvTPGD9XWUFg2mFX+51TjkYm4+EALGjQL/hQcuow0ovgxjYy8qGbgu1rthN
bNCjgMnpZGq+tTshbaF2pCxgKazpP8+aOdR0ioyNGtdFM33Ee4tBxfcaeUdC6oaA44+3tdoGD7l2
PcZ9pEdi3Ys8L/AfZfMKuKZ50TMa8oF1WTYIwVsKXHkJ8jf4mvBrMWdqkifvj6jLukZBnLbXZr7W
LsnmwiOsuO87zcLBsmUS1VPqBd+FAClMhUYF8OeSQbGNB5/GnONLqQ1lNbgtRtdtNLK9FClN00bX
FPNyqTGsQUCMeDpdOJJ2bR6z1R65RuauOhGuJZWGqd9YOJTTs+PoHhz1wmqo5kInioQ0t/OdFrah
M5tljcc65DM5TVZwcmhqDa6FnIzbkcEKlQ1YYgM2BNVAm4MnUruZCZlv3t9UtiN3PQ904yhXG5WX
orblLjCWePDWZLxSD7RN1kSrbOHQSf3rjgN6KCbwLy4SpB/qzHABmkuHZhPMpDmoNC3HMCX7r0xP
MAlEKoBhGV/6cNYnu2uN6dX5xcSla4K/GupNR8NqErvdOd7jbVHcWYKupfUKFZBKk200U9jbGoA0
NKtvRB4XOwUJh1pqXy4xDzUCRybI5UbLQRmFy1E0ZLEftYao5Rb0PkcjZHXUvglZ/GUyO72MXCTY
B9i+Nc1s6FnJiQ6+kF5pfhNtlrM9xl45xVrsVxdy6m4rV3XPc5JF25Zpd17BZVSXToZeIy8wMwuQ
Rca7D/z1tP09SIbWYq7BI9TmGvaZn+XNMFBQeRncuT+IPam+tf8KyeVxuBN9arxweom4dh6VS6X1
zwddwMvjZT1BwbL4cp68fnRu1fCCjMrb2OjIJddfheiCgEkd5gaG0K+7KGpBXTxF8uo5xYSlYnec
naW4qsBPN4SvKNBDRMPxv4k2V6O/ZDSE9LpBIHjHY2QDutTI0j5DjvQzqetKY/PTNAYbiEvcx2n0
KhixMSl4m7WPIWkAVt2Z6+m/vnq8Wq7vhqeGijsc1eP87Iq3byRmnCqjsLqsAI6HzZ/Dt+vxyc21
DKXUYKYYVPl20sEttTqcHshxOI9AJVWP6qWzQIVx8vVRmgLaHxIsvBogx+WKnL9wx2WjudN+ViYY
EadeqDsgpdl/Tjh0yf93Afroijelg5itvtazooymO40grayRjUBSzMyXtT3zXu8FFROSqbkuxkYO
5hgAMiP5xrFNZ/VoYVy3dKJ9MglTED5igXUDzG4hQPnTeElR/m6+3+sqRePOwRhDBFBQBGMb8hFI
lOQVvEVJ9r5f6uSZ2U/YlPRXF9NXflW/4ivhAyg9j9UQxqJkSvP3T138ABXSQsTDMtm4rlDw9L1k
32kaczeXC63NzVJeFV1Qn1z16JwtLKQlroIsLHgdnQVQnZLL8oxRbA9l4EM9riO3nPEGSrBa30Xh
NuIpEcZqYx7e6vrLq8NcaDzN2FH7jTAX2ZFh5uMzEBEYWhlxBofSliYRC9laJ9wxIElYl8zuk+tq
eLt3i2sVR0laSYlRqOUgotOVhhcf5LlAM3vcOaALjPSJ87QiGA8TAF4P5zdugCdyj1c8bpjnzzWi
3heh7BYeIbTfuw4fmmIpL8RO8MY+H7sr4yKM0e0bSBUWA9iSm5amAFJJU8066Pi8KIzal1OHYG/q
60OrgT4IZofES3NZH6sqfHaXcVttdqJbz4bOKJgnEYrT6/EwrBcV1C6i7J3hPT95+4JGJl6aAut6
KEcKTHkTXW97xXLbCyRz52zP9QG5hboVImqeNrvpFLvy9cZmz8ff9EBs74lcj0j/voQHsIY33rMb
+8hO9B00ZVc19hH1usMfZW15Jl+FJvkNPyt6us5uPCDjrMHfOGL89CPDKTgObCXWVVO6N0lHVQv9
/3i312iq1D0Oh315BH43/aRebMrlbpAX79mkXX7IigWu9w2jZA1TpGk8q61fyT6CI2RdafOh59v9
zZ+P3zmZKza8roKHOgXGXOmmeO1YI3THwFg4OO7MCM/rejIkpDcmVGWnTjP8CfLXqZm1TH3B2wmP
q0a8HDm5IB02FHVrMU/y7PKi7xNAWBoloF9i/BsrAnrDhLNuaH/otsCvEplP7jW/Tjl2J4I1Tz3q
HJSaUedmsu3GYB/y0BZoK2Vdc/1zzwe1VgVlwRNhJEWedj9k3NtLPLCNvcM6KhInKKHNQxONfoVX
nClKYX5gZEHY52oMW0RkniTYn1fHC/J8mA76RCFeDUUod+HerTUv4VGTEuS0B1SXOpAzv2r67XB7
z1olIFd8wGL+QJrCuKJjLHfPZ7C88TtPtn5hKn1elQUheNxhz9VT2qu9LDTssNhg4vVdPjODb/8a
gVdUcZdKMooEW6JoxRehnQR3nU8xJGg46lpjtHfH0cXb2LIMTFq1L/En4Lume4IBK2fZ1h6N7rIp
k7JlncmyGPRFeNUm+Eek3GOfJIEfTyMpV3NXDsnJMcxswtXWq8gd7sinDT3FS+2cnq3gHfp7pziK
UANQ/FtWAoQPWr5H0HzoiowE4pijDnk2Lt/BGAPKJMsEhPjQbmW63Fu6yKvhYgM193Yc+OajCkkO
K3xwIA/WKZp2JKCbmcMSIoaj6v8pK5vcjszdZFfOOF/zlY/9dathfIoYf0oJ5z88Um0afalCfQoB
9/QLXODnraccE1fEViKS2Ix+k+tMndQtXOK7UMxohWh21WJJbi9pyNOO8eMbMi/lwR3myNhN0rQi
t18POCz8eRp6CDKnuCmduqNBU6uC74M4loMr55kI1QXtkixz1O0PVlT/C30PycqpZIuwuBDxH5aN
HtmIRjJagpgxS7lySlFQ+E8BZbstsaC0kKmo9ooa2WVRAuQ5B9DVOIUlfAW6V3k3GNNLjMsW17OL
duMI3Md5U/PBeUcl9IRKfpJx3YUAueHSRY5ge3If9ClrP/pCD/jXpBdARLh2S6Lszvhg/9UMMtTJ
267g0NB+6YeeZgRuyN51FeIFgVUTvEeonOKCdWY7/7VEh4IaK+YqLhzSeGzt5DNfe5tGi4QVCvUt
oFLyImmPioutmf5iqlE9M2O8dJ4YyftZmtzbJPFwGt46gM5CB438oBY+nDWj5YtclG15rT8qlVv/
hDE/ddcelM9X5CQTMYdL150AoANyJltrUk4shwSh/gQDt5pMCsjVfab2mzuu9V9EKr+NLj+zGWSx
htxWmL+VlVV1BO2Rc0lfFpioOlnbmWs4sbK4OSzdW1W29u2usQMbXWIDtEINUeKnb792S7nekvPh
I7tGcJ6uif+c7PbxBfv8vO7qybiIuMaSqttjGp3KxLsM4genU8fUND41xnlDOfBuLEK5X6zdQTK6
WWXasqadRsrrFxYodT5yNs55Zhu4hTyt+9icA0d1HWB/DoBbEKwnwgcHpqJm3poCLp3DmO7akhdS
2ZAjaIJ1MuPWntoT0kXdLPBNYvF0N00WGGsRYcYKCBqSKQnqiJ+XUd47ns4MFuBUAP+TfEdDdg9R
Fc/oMF70YcW5IrQiI+xg0J7GK1PBu7j8PqYZTRqEpLENwqg13hoC7ItKZqWj4+yHQCQJsnJDwCTD
UcGLAQU5csB0D4io/MlO6b1adcUBmS9AqSXkLgZy+UiYn6kxq1nmrK5RDZS80+Ol+PGmPfRYQgZx
HQi0zzynDXCXQESW5j6iCSg1pquMapVWpIEe5WJVYTpPUcd7SxNR8fA6PVJcyM8dd5YtE8Fn4EVO
dPJHArxUWsDeU0/4WaoZGAcUWKxqUrY9c030fo8hjoA+NxrKawILusQBzEElz4MZb1hK6ldyI7yK
n4AJr8mgY+K9eWk1MiU0TqXv/AHJzld64WWZTuEO4fNmsNW3W+qEv7YxavZ+wEdrV2CENKnuMx0r
HH/JA4oPZJWGur+NFqO0iJdQFwoff67JXmFzfCgCFqPDw6pyfLvW3rSvwVhvhkrK3n8Ocw3zzXdD
0PeyCZAjgCPzL3bCnCkocbrigfqmbcT2uqoSJxrsvT7U3KG4Iv0lkyjdWrb43Y7yqEVrdqrQnY/A
nM8CA7sdpu30wpDKbFKD240XgmN5wwmiRNqO0XJgeu3+jhDgPX8C7ioT/yCcyvd4aMiQqRRJ+6Bq
9xHqUZNGSABzQcVEbWr9ihjsTB4oL1pRGQm1MDxy1mLoLlA7VSJozrj84xGQEqDl0jiUckA5eKmw
Uy+5aTufkIPWxhIJSVljRzwmhcSc3kRYbJctFJ+ZPxW17jUnPZGgWCrTdtUESrfSAlzM4IQgoT0u
rhAK147CPQDhKlFnLaKC/5IBZ7MukdoehnEd1XZr4p/6uQGMzQa10qFyRVbmz4AWR5E6haTf1mAF
7GAVIebCPeuFQZ1BdpJD9ZTnNHFQ+bSbAO3DHIHMjs9E4W2bhbYnuevCyraDrMkGX4ALQ3ceBPib
10J0MkYhIVI/btE5j8BcT7OSeyzRhbmLa2E7u9IPLuI7lc8wQpR1tQRBfu12TsazlDbcWiIm0JGp
1NrqttYCS91ucIuOOJudsEo2ySAHYeTxh7vGaYutsKK2N00izKuc7IJsmp1KlJzaz2PuPcoaxrxe
fGhp6auf73y1FGgUKakqOcWBcpO6oZhjVu38s0HgJDiLMnncXsvukOXKE0+kVqRdODKRczTG/a28
h7XdeChAveY8qRvYeNf6TFIz2yjdvISa40wk+c4ojqOLxRWr5oue7djZS4CJNwSrzTEKv4Hk6nKl
MwsivUebqywlF2Fk1Z8vglVhofaitgavBbUbyXSjXrpRvXTeIoLA666y780Y3PJyiElZoDUD2Qcr
qpoJ084jluUSf8UrMl9n82DTfLF7jVQIRSMgUrNcWwPMuaUyToF30LiU0yTJqiYOkE4EMj1vMvnU
2E+DaEf9f39Me4WpxXK5/v1ItnXbysRl8bl31pAc1X8mhZXBDXetkSfEKTdFRU71vstqMjhVdzC7
L+9DqiDFycNAGpUtq7V4oiWStTlEGeK6g9ppEcS3jLKT9X4LgsGyZMCLb18Nyn+BBTPX8giLdQiB
7VYip03c6DIvXMWALKuR60WNO3178fGZll1NcgSDqDCSjyaZicjTEUgYBfvWauaVsJhGhKiirunX
v9kSGcIB4TfqsmYcCKiQZa7Rm7N3yg7hbN+ByheVC2a0KTEtypeWY++OV9Wqub77E5f9q5OfttOK
yBH0/4jGrPEpvzynt0pE2KERYEsVp0sOB8I7J78qWpYftFqTJ/7/SwubkqMXBL66UH/+tn/gliZh
oX30I1k3fpDEWuQE2osejkkqx1ZULbaKJk8VqqAi314kXe7ROLWa0+yNT8rfaNUY1Wj2E3JqtryK
gqQHZZO1cgLGwZU68Tz/S/AvKDsGid51OUNzt4FWDTigNmgHvSabob8jShgHw5Wxj5DXvtqoZpan
Oci4Hu6n6mFV5y1pigPQhJ36VHufgJeSgECNwBWTLGjkDX9wFPM8teM4QU5AOnWD3/E/Bue5MHs3
XtHbe35g5xOzP6gGa7BswuNWIYflxEUKRjJxLxKeBKPadzziIVFRPGVHI7zYk6NqZsErf8gHw+uQ
qstZ83OQjKJ4QY4n4dtw3c/NuoLT0fksB85vI1iETlyBJbFUapCGuhoL5r4cCgLSXuDW/pBDW/Zo
QYTnF0YapYW4rsoVqF7PRPxAQ10cJ3E+ylz42fhsjytH48FQiOUp1AOjwDMqhGlkHH7rayUXk9bm
r4t4lTW9xjQHUdZ82N+QwpesGD+NCnX8Rp3LA3UsOORxzt/e/+rAucWEyDHVfeW6fV82RDG5qD11
9s5++bzZcEB5fcsOYa3RHa8FzEskkAmIiy1AC2y+xjJUt/NqEEXyJ5yw20NtF/sgPRN2zqI5XTk7
kEvkHK3ghVuZRkODKWPjGm+qcDsege+zK/UqwwZMANvhPZAu0jpnWcfmR1N9vrN/auRVb8Xdg0ML
M78em8RbcbiAOpo49qlBFaMO+WVW2IrHvtJHvvMBJrEmSeQDIM0F4sXclyHRbVIe4poZpbvJf1U8
3JpUcJgeA5zPVgLVnQavp2LEJ5dJy2rMbi0aJZ0asbsvsMFuttu1QZG7c8Ut+fzGJHbZrHHBFbks
QhKsh36JS4Dhzb4HbLgsvGDP9RY5gLs+cJpAf/0hC66oklFOu+cG/C96OlfdNgiNV2tayeRqNeob
sbgCbxX6HILkgiIDWfgjkh6mhdCP5+X+AHyEVX4NX4tLZ9BrLNO0lYVCsbYsDHiUJUIfs3yeYIz6
gFN71a6t7r6Dplau4JmI1kmMszWYSy81efIdKy06aGc6ySE4sIBoNwM6MDIM+hikvaXoAfZpjOqj
1tMFI+mwqgw60J/HkPX19qRN3XOouAGT+uX4RH9dbO6uGm/Tizri4KIfVD3SZv2OXydsIDMkALKh
MZvCXeOhU0HFwqJScBkt1GVYWxrnaZufLCBokDwtYq1o6uTXwbL9dCTo3o6it8i5yI+LnFzvCXKG
6cAoBwnk/iFYibcSa16mRwOvCFBhkSk2iRE/L78+iklcD0GM1x/nkOJVFhn7yTDHCjNqPvBQZ4lj
HKaxnaZlExSkurMRKaotNc5jgofd3wpdu4Ctxn5nzPA4+0dqoIqj4CKwKGpeaR2XeafzHd0AyOrh
3zeNM8lf+Ew1ZzmswUwVybgs76e42DStu/Wn2+yp69qfOyZ8nXsSk3Jz3Jv/J7pb1YW7bqAgF7Rq
rIFow9rxciGd+3jcRHK5eaJAq/bWjxpMyEicwfeulYnJwx8hllB/hFVaw+/uCElWnfknTk2rkBPL
qqedeQVc9Z62W6JHCD25UGidkIi1uKkZyQIGS/ZYxu/o5PC7MWjZMr2F83mZnELd76LRNvgWIfTJ
KsfuDYNOcyfR7vKQLfoLjx3THh+DG80djT+uHyRoipl9kB5pU9GoMUjXisizzZjPQIwWBoqHQA/q
p6v++Jg40FpPTs0OxkafxhPK0zASInUavH2921s/+zu5pE7rfXeuWQGtBb9/+sqDV/CYG+Ob9Dp0
SS67TdQumvEHvyW89OmmzYiRfqsbYk4wgQEO2BewSIgr/hUMKbyZ1ZQlmtAJDgRMZCSTSJGaAKwz
bcxkvbH9KE94WLHgxSqtdo4W+7vJrhH3I4EBIJbLpAyd430oTiRqkXnxEgo4YLXDG7QV8R7HDuw3
A9938NGG2WM1KhuLwmD/oDmzN/JQJQ0++Z5aUGO73of6jB/oXgXxL73gDxuWLvVstVcL94H9GOKA
KzJ/TjGoNr6ej716PaxozAmwNePXtQNmZ4U0ACn8ZA3OK2l+nswOXUOSEOZhzi8RbPUzFMNJuuQi
x8ZMZXcI5De37CqPsN5P9IElIqISWSiE1djD5lRs7j44tXwZ19bo5GHvNvnVOICEZth9C44CRnlC
T83AqFd+VSEs2u/Q35n7MBEEwAnqk03pOQAgtO2hz6lCBZZjWVc6pzUBp3ajrePH8O0udToHykdO
6bIyC6cGbvH4CMfxuUdlUxI74ZsJr0WHJ3RiHx9ut9BGjU2KrJNyqWxwYnDN6ZXICy2+NFzT8wwK
qjogKGVAOojQSg47wfUsS6jsHYVByAHYpJ2UBAFUNrilVH/fp6Qm2zOydtYaf9Ia9xFs+6qLv0W3
KqoVKoOLskaKHKcsl5kd3Op2urxzjjjpC46LPC8rf14xPSrujTw9Eg0lIOoxZvFGY8YVCNMisSoo
D4EZ9OeK9I2Jzu2RPe8j8pfNiK3DKE89TiEZr20hvpb8xGuiSt5G+DI6Qt5VCX/bMaHx7I6Txwc9
sVGVuY+T+eWUyBoqRuquBrb2hLCWmpeTk/us7KPAB2oI8heTfHPDF/0gXCwXbAHiUT9DDv4NnVj8
HUYPqU9aG42jItOL5bEyQcfPU713VmKrflwhVbUTHjX4Rf6FQKEU484/ms1ndq3bp6fmhOX6dItM
E3kHbJpatqbpOApzvIIDyyTlUfqw4m6LWVgmCzh8Gsai8MrRnqOKMe915ud+lJbZV8ixEQIS3Uhh
asjimXbbG5DjCq6BRVkahi3iDFcFWHwsgJxK4jUGKX5tfEqVM7xP4pKRGJTPp+X6dBQ/cfjOEkc3
VtB1eYgybUlUsbxgznJNRuLtJ8vqqkuBalJT8tmth98vcqIYKf50DwMsKXUwZZ1GVh+p2yx6SDjb
rmSlDCnRhn9EJVCiSp4QmJlSIjcT5HmEezcSSZ2CS1F5N+W8vDn1yvoOVOfcIHAek5RjQ+WRTqJO
ezQP5RTYC7eiWFdqQEiRo4sQBviNZbwXYw5rXLZE3FFSwi7/UsrkSkhuys+XELhtQJUcQ+YxeVGW
6PiARScZ40x1+AmMpgo/e1pUF2k67C6QpUIGd/7P8q3x7qKhjIhIrnzco/iLF11geG3Lkc7XANlI
pStuMDgORB+yIWHbRIGbVzJQuIW6L8kDaqEzrZM8y/sVh3pgPcZbllx+AwiFbzmZGJ5GMJhaXPCY
uJWONdx4IViIcQ+m959AFp3IrewzgVC3iXNcEGY1f02N7YL5M0TPDo6tly1ynhA2m6hTh6KOUYHw
MHa0j6nBglApQV+MuDPYW0kmfaPxUq3yNf/8xATUMmyAigYJ37y3g+gX71JdWXcV8D6d7nMSHk8m
m4kSFLJ48OdxJbtO3pHWSABWe8Pm7EmczBnctIFk99F38Bm7XDpGY4xV916AVbKURnwVST0az4p9
5ANZq21b0D9kP6Z9jipqqNfn4QO2+jDFiDMeBvm2Lxpg5Grt8msWuGJcxnkNQAVlKOBP6Tf/Ldrj
FuhNBtWmL8ZaT/bGrS+HeqynmNu8LU78RL5Nv2tf39wrx9Ba5523sd8jCdE2pfw0GEyOXxIIBpiJ
+H7w/iYibK8eO4SiFFzGu+O/MWoH4Dy+j8ziil2XnzCZD2w3uvszzo81XfdLIXWUbM8u6GZpx8R2
Y4DZZkSvh0pbKTY1rjqh1du6jfGAl+FNmFgp8q6cUURzdzlbGFtuhziyJuZusTRXO3gBE0h0oCHF
hXviwn2gj0QGXSLnhrHsKu5Gj5eo/hIrygx6h0wx2ki98UI6y7UYywOOL0dY4WjvpqEuOkQyGI1o
VxTG74LM+nF75F46IRS2TqalifB3ZvsmzDD9oCHtBEt3Qhh4KICqlG/9qt0gscFsuARtL2/C4j6U
ocs1MsmWOYlHjd1Iybn+w/It5XFIdbaWcmuYvdkzX8LHwqnBuBcWOmzg6CBUjOYGsKf883IvCTMQ
knzWUZT/n67LLX+Qj8dxSFbrG7ZCK9Hc4J0m0VimQ6Tm5W0g1SpNNpRPcGWtGzpiCzdWv/OkPOV0
VX4HIqeg45nYApfY08J4QadcnQLahWXH1KmMn5tsLhfCDeGULtAbImY/8rhGHlkrgOaJ9ufg9SgR
/xeRZez4U1/DRyEZIKz/qTEAYwX2X2ci432wt5UPfSCmeYydn5+gY9V6kpPG75A7N8nPHFXq+A78
omlVcC0FSdvr8ZN6Uc4IfqQqc+E3zw1pHT/v8YBLqXY2m855uDH494MFVVlxGaNjQ5sUMUDrAdgD
a0TE1ltpQ/ySnxM2gHyK/2OhrhBeZEfrOCYL2n/1v8wLc8iAsaNqbaSLUfqYIB1bTVMbFkAhmu2A
79LXypdBgS6eKT10ZDGJFWrj+tkBWDwubzB1QzUqD0IGxQrFD0VxF34H67imz0mLYwfK82En3E2l
J3Jh74eXpuy2P8c3a525iv4QTLDRzrFMq2WJOeMpfIv8Rie/caALnMxuPZxJciPKPE01cpd9PbYB
lvNILSEFA6BLgy4P8aYegV0izvSdVY/F8v187c+ep3bz1I6MimPJPh5UbajfY0JHKw1dYWOJpSx9
DgKkfAM73f85Ga1Gmj6S9JZpE1BeFmHWCuQyAZklfHMXBBuvjQJNU+GSkZfVrletdudHvH3pMA7c
XyxtvIUtGgYscBj6ngEt7du6TVQyEJrQoFZpMkQ4ICcf69yhB7UYQLI2CglPlhB/YWJJ79xIJ9Lx
B/6SKX6bYNjC2O6ouA3y/S9bNwWYPi+8DNHD4vlR9/ZHYmf3YFSksEDjjt7ONNqGjWCJT3byHI5O
TwNvn1CHof7yoX1qtr8ZG17RyDRt+WQIKF7XZr7QCIQaBhc3p+0KIcNWkUjiqceOKc1n7JDIq+o5
mHTAMAAZ948sXBH+T9ga/9tCMd8U2eDR4ZzMJEiBn0lKf/1o5eUpkEaplaV1t1t61pHCtd7iJu05
n4DyIDvF2T3cB9IgWQKhcYMuizdvOIOkkqJfJdea4tp/KHxZG96tRA3Yal1gsalTXMtyQdM+2YkH
PmiIslNRdTvDHaFsrinUMdh8k9LnM4USVg1VssowD+7l/rT/WavvTd+n7wMgj5yzrIR75DWBH1pS
h7W2g0OS052XZ/WbxGKMGf2i6vYCVb2wOtZ4WVC3YoyZd6gBPcBwGSjYOX6iNXXrUI6jt8qfeb4E
LGAgW3I5q3LX2KvjVPd8DaY4Yd5lBhWwjzF53ZKGjRi/gVJZZ50bI9TjOyM+5janbdJjM0nkrcvl
tife6VXBXpQ4aGc4WTq6SuUwbQgDLzDFOw9DUptLaCnYxsQrMFSxtCZLKcmNJwcDcMwQdyK7pF2L
kFU8Hbk4I8DWmbiRF5ZxOHKvxSu+Bqgj73F7BXNMJammAcQRUl//4WcztNRap2gqU0TlcOOcljth
cc+MwsPrViE4F8ctHv6wIkMEa1mJd/ZZgmNoBgMeXL3Rl+mvcVfkAKedxJUy6vJYU9HOnlWfJgu4
OPdQFACZ2J8ZP9QBz9TzjdN5YCDmkcJSLL7bufP+78o72oSLqvVuSSrXvC6f/sXRO18vrukw65n3
hXfvhZuIUBdQLC8nJHY02XNTx5m5p7W3atNTNPoz4VBBOrLxiWUUEjUkeU2vgTl6Zo7n18CViVe+
RrEjHVgTGOleUru+zXgKQFFFj4/z1o9yrQWMA/DyBqhJSrn+UHvGKMnB2ujIu5Y7fmLTfrV528aw
bJrkEE8tvePoudGr30KqHhXo3y4FVwm9nDa/BE9RzrcGZpfoxYRQidN2mNGI39UV3VPSKmuD0Xll
0QSpIpUW4b/noQi4HPiMJ6xTPrdSNTkPpw75akghIIHcbl2/8JK0TJgvGPpSM+SuVksL+Y/bQs/u
VicmzCZ+cfd4aSA7XHeFDjexZGjIUyMLXXfzWlaXwHPXOtWdekQGnzVpglrmFhGbisVfxpLruI57
6i+der6k73pI+g2V60O+7pzTI5AondWWIjC4aCPZiXoTgpeeH0htyDPUHm+9q1k7tE/zpYmLQs07
OrJnYVRXRlCrLgdMW2VsWIBpkf9Co6N1C0gToCLrvRTiUK7fGRmI4+6JgJVd92Bw6cXdqh8q6eOR
cMePWYy+7WDw0cRRQtCanMedRGRBLNreRIAq+VRuwKnzUxdbrrrhGgIhmN6LkctEVOEyI/cnR1Nw
XkdiDQMibC6+lBYuPzDdXdKSWSpSDTQknerXWx6H9Rm2iXk2IWsCM3xxW+ztVQLDrBsenC3Wjbvw
lS0OVOS1yRn7FzmZG5xo/+4aIDgglLzaF94RPyRiSuKkVaCfUf/gwzV9U0g42JWy5dS5itVu3fJX
urpvosLFZ09y7kFiwmHo8JnPftmn3FCJQ6/ENcFUJsg1qKDPxcCdPf2vNkWQaPC9ICc4HZjcA0Fm
bFVLVC2yRTQVyRE9/mgM6PRlYTd5Pyhm1KLTa/GMuJ6H5Nt9WwSKYnSN5N9oOzW/f72UO+QPStWz
LnzD1zQMXpdr2Leyq70lhzLXraOczTdM4nsMnVf0L9LNTzl8NNUKefdToY0YEBmgxvZDA3ouNvd+
6rhOEoIvPqyT+0q+oVd6J8a+uEUg97cE6hWhrhUHCul2IwS7AosS+RU1kBD/Yw6Q8JchJSN3E+Wd
8GhAFoEl8zDINdVZBA7UjSxeQ3ZW05Cws22dNHR1xaFGx5M/d1n2xfg1I7Jenjs8KxaGj6Tq/azl
LsA/clKh8p+AUvJZFXRVtl8ux8ATUZV6L3ZlpwNh7JTUhFJIkpIAD6TPjvexQjOirBbRP7cOplDY
utjwasZjzIR4ezl3nGAFXYBVoq1dZwTTAhSubNcN+cD+ScRg8oVATpC/7a1IeYoo9aY06LRP3TBs
rXWk6bdtZQPt181eRd+D01ZCu6EIZJPPggCPrdMjD+CzqBgAXWk0OKsPGnwZ9OSEhrqDNNM+zzIc
nkFaIdq0zie6l///YkvJSa0flbRn4qqjZvaM8lrsoClsaNYS/cMohBPG1qYmRXSj4p60cSMFVu43
4pqI/bABrb5MJR6BQxcEmr2w8CxwL+XYpEDHjWwabmPVQA5pfCMN6psRA2mkjgUTVVjKY/q2wJRH
uJdy1DRqywJq+XTfgaZgKhUC0rHhxL9LJfUCE6Ax6j6c0wAB3ra05p1HwBAlfb/eY5uCFDHJWIrc
+0KVXOm3oSkR+HWSXPiqQJS1S8cbcGDZK4fa5fwfL7JtqVQuFiT9GDRdv5UgfBFii8mxW4flk9J1
1TVfYn1CluFxTF8qswtv8bqJNc/iPatMN7bl8AGd6Ei/rM/peGt1d5vlO5SmUtYTeddIO4xbR3It
Qk5VMe8LZHbVTSAviWfYkrunJXipmxkkeShA+Fxy/16TNAnHvt4aXrO6oYqR3T+OeVRFr/Emt0Ry
8cFRTidGwCng838WiAHyyP7f50DiJby2icRvigd8NwqyOMgmcwlsqOPdW78P4T03DwsXveShEO9+
5e6QANi4WiEZvrS3dYjPydOslTSYdOTzaVDR2/T6nK+g9FmybOD8+nBgoOYQVF7U3xSaH6XZ/a3C
P98qat/q+38Lq+jP6+x/tvTuVpOCjLk9UlH3rb6/U5QkomQGMSvCyqFFUMwb9r6QoagnlaSiE4mf
WjR05OJmRIhya4DgDlX+gQy70B4Qg8ZE9vPvdqagHDJVwL7jQeYMAIdgu/kZ6FL0n/pCDnAz6ofC
0KduO2LExrLJ9SEp/2WHXFC1ODS+CrmTZ8mtkZxGWj1WXzW93QEY7ppBGenF2qsdVsFXzv9xg6Ue
EvLO06eB+MovhF0HN8Jhdb4OxSZLNxhMnFIeA2gAzm6Lo7W+v4rEgMVgJ3PAqPI/oOKPfD7gK8Kr
bSRJiETScVdcX6e8yjnPFjuMceqnCHDs1aC1aU1zabAmgNC+/O/9kk0n9mhWngkVnr9ab4rG1+AN
xCoXtzqM216Ab2FxI/OV33mMj6YmXgsuwmlgD04Nsu+PGHuEJXut1HZErTNm0s41IAm/fwNqPgOq
yLZ5Lh/5H5cI0lHtV4CjaB/o2w+k/yxn7veUR/x80Gt+cph+qNAj5atYGelQkQHmGFofpuZvInLx
DARbtp/gsqUl5B1Iu4gSYLvrf5qXEJfYwFkE7u8OYBoLPE59vKIJ4fu5/GR5VmvpSVWkQkK5jmHi
+ieYS962iI8uFWh208ULRFu8F+DMBs4mZsvwQR5zUHlUsjl9ODYDayd4pFr+n/7F8NK3YKk1iTdb
ao7WCHsZWuywRjtxEMNfkUgf6z/2v/Vi4cgoN0zxjjDO+F0g+s99X4JEOOsQlH9Q6FO8KL35IIrt
ERicmE/DRRm4dSgdZM86x2W3h1fnwvtkM0n4/6c5EqEJrhWirXWXXG9NardyuJoWS+aVBn12uKJ/
l5Q9dRnG4mOvRRFvOyd7Ble21Zcq2QAWovaddi9Un8GvNu1TzCfonLb4B3UekWpeuE5q0nwQWNo+
Po1OK8fp2OU5ErxDfCFrJLzrZyZVKkVpMyLw7zgCYCcjojhBu5nR8xDMinT1F51QITGjjt4Pctni
OasbDbWbLT27NBE7tkipx2IvOYjCaTSFFu1y/wdjBiCGhhAS1mboSoiHf8zQAh6JiJGrjzm8c4iF
uyAY7/23RQZKUtm/S4AyPZ1HSpNJKTLV0y9cGcRafAOrW0uCYglcCaBFZDhM2B5PWJ/La2b0cVM4
MW/tteE9j9rfjlvzaMMlEwA0tWI62rJswm/QwmlptWQnOv0JX/EVQ7DwvAvBRzXLfnISViCJrIsL
boyjS0234phSORQVbTM3i1nU39YVjcj1oihEN8CzD+nI8VNEiLwRHuGpGFcehxK/JAt2x+CZuGlz
FuK1Ch5UHHqre5N4Sw69wFm3ZLwR7YKl0CphUBIIr1tofAmcu6JS1UbmNXRVBAQT/+3ZlGrypJrb
8fD0G/BWgoDm/gNdxtAQoQGSVTodPlxlJDSb0QiiNoHP9nw5jv10ou2E2D3URZgKGDRQNwmK2dRF
l9EIfHFGRqL08YknOGQSbphAb3FjNlYIyM6WTWI+HoR4Nkq0K/u+BIK+qS10cIBkH6xsZFSmwSvg
SAZ+FdrW6LcLyxnf6MxUhrdu5H+v6I21Rq/vdSdgtnFElajcNHABU+rmCcI8pUEhJn04pIk3bDtM
8oWi6Fw8guZnAgkuztoCRpNq1Mxj9htJ/wyWfjCCvyZE6J4GCgUxCSo32yPXesWpwVMUOJJQkpOZ
D5S2QYcwdewlN9LttlwJUEY4GR8pcfF1LfUHykZF7R5+vdNJJnY6xuJa9sWB7nCOlTvWieEI8Sz1
3vN7XndE/H4QQXpeCIC7s94aUw5tyyxx6dtNWvyP7MLtPmrbEX0E8A8otQ/zLqANPIcygwqS1fm3
97zZkNDpLjBZ2/b1/I7OTXy1y5hHYWNdcljbLHgzA/TPcykRoCq4msWjDTLPEdBJtAIJBqZZKFX4
XDd4wO+Xnyl7ogaGYIK1BwIWUroviLJg6jRjBDbGQGCDDPKaDup9N2jJwXfwV7zrAeqquIDH3TDp
/Ye/UgR09na9TwzfmGaSuCgUyhWJ5tdfh0XOFkv8TetZSuYEKEkHcwjBsv0B6ollq6AGUsb91jSj
ASRmlRTyTmmxFv+ahy/5NFSSpkItdz+qzhoMZA4Mnvh4J8YBKV8sRjiF+lnQLN3YccHeFtN8PEST
tL3qJ6zl+ger+9qNWCF+e4rz30ntOfxzNLJpEr8JOh5etHixsuEWjRGkCcHv+n9wnEhMWsKP51b3
wtBU2hBUDqlh/d3IfZCDZLhbN9sXBqtDvJaxUM6tNh9IbD+2rB5+g5SYRmAARRf64j62xl3ra/ve
0OAX2OTEQBxWoTO1TkDLUgpbfV0kjHE3wHQCxgiqTgD6LnrmpgOggRLql78oc2+vp9RTj2OE5NPv
koFeRw2R8lPRHv9ALnO1/QhhgPDoZ8dv+JQPr7tc1fPuMHENA547x8CSJAFvp2PwJtPCnn/vKifJ
eP++7UBpBb4QgGUMN1JhphjeolZnp31ejwpRNvf6TCwwy8mGQXN/mM1HiA3fcsaC+PE3fZzvVjft
pd/mRt/ZH14XN2tWZMUjHw9NcK0GK2lzgXnvTCZqKVdiOKmPVdD/h2HAyvlgoMpeg3LcHXekTDkb
yH86P+Zu2rcBxabb14xLnL/Der7g+g9sUtNREVhPODyTBlvwXihAgUznUCt+kO88z+SYmjtcM1oJ
skwJ9UySlW/i1WK3KPb+CQIg5o7o3qkReACMqzEcIR/kg7NvKgUOGFUntd+dT7jpzqE1fM2uFrR0
UePyxPiVy9g2x39IwwaiOAnB7nvhUN4va7Ywvu9ZWsEQghyldVg4qIFqzbJLKMjp1aj1f3fZc+jz
ZUseoniG/VtkYNXBvtOcPSB5GOSv84lPy0JvPQI5xlAG8/tYUcu+S1ftoJJ8aP47WT4S2v+a6LQY
Pwc0N5BNUQOGGPvMM+585nW+m7fQem+Q15tswWT5o6yklC1HAOyvLg2/7OBIYeyEMiMmCbgSENHx
WbwypR8QpR3jb1c/cVWaRkPoU+jA6Prl2sNqUY1fW7pFli4vPUG1FpErUCeMmbPCDjJtbq/gRHCD
ri+qrhw46uvOlVcsNzuZj06EvS2iqCx/dCfLB1Za5vC24r67+a6AYlo3IL/Gx/Ty3ao1QQVBdspP
xIRUweGdV8LM8Z/+rpkISFjWlP9m9+tXpiDJqKog8RfBgXsUp/UcPOdoyr8ME0iSDqe/VQQ4uFX6
l0h7Xbysku4Ylk2vElfbGMc7Vh78vM5vT/Rxozx2pa4Ry6/DJsSrQMEdiPQjr4KTxyKcZ0ZQxppK
Wljwl+zOJGfNAlMAmgxbTaM9NaSoh9RFEcDdCm/pcLQ7vaYdFQqduaoz7mg1uqoRLPUv2D1jmsjT
ZoxBw170VzMQ18NBex4IXvMvk1GxcyR+2/rXP2PgU8TiX1wvXtiJ5IgL1vBlvCD35n+Js3xey4VM
Udi/jfMzRmn9Hx8TDqquC0usHjgvWwq4LkkMVUMf1IxCerfHgcBJddyhmBMOUBw5bbTWbE4EmCP6
I8fIJd8V7wSBLds9gW7DML5p5gnGpLUEcJrw4Zb058lPeScAHn8HNzX1zpY14vEmScmZ6RSiQJv4
dcUu3pT2oAHTPfziJYU2ifM4WeSU+gDEzHshyCbh7CBzMB7UVd5wJ9r7A3WHOedn305vYXWkqbQZ
4QJsNlOsyVUMMUoEo1v/5GkBlYEZ2FKM9gF/gPQclml9JbH9M1pCEVPHP+4+8NHLcMUiwIGvcExJ
qzNMUA+axZpBe1qlU0KZWRhR4UvPWn1RoWUTOMxdLX9VRiAwaJL50fX/BWy7N/G/P5AcCgdtbiNP
GHPl0GRxhQfmGdc/1qPceXb9ZC7wgc+QICGbiQrDpnwKASb32ZDNPoD75c2JR3xLubeWTzyX0066
7V0pmMJBy2DiJOE7MAkCQSJdnDva06Hmwi3sQfeeh+wVITiuKCoEq+fF6UE1ocYjV2846Uq4TroA
Zv7mmaRqAo4IZJ2HQT2ha4cfFnceOYFxPGkF/qDNB/t8036l7eBB8XK3lJsZ9W7nOr2DmuYv0hWs
92NOKtiKwdK/Q4lFHfnAbu4AzxSi5DcDMONvTxogyc447yXBr9X1Q+RfGpt7EZH0Oz04zKbK66Sc
S7Sc8Vvw5809Rs1eAKQgTHy5aEuI7Cf2DRpbafCdb1oczY5JoHcu9Q9G4tFVm65ycUzFDNqC8xQc
F8fLX28ukTLLO/1R5rfTDmcPS1MgHicMRQH0Kkeml/eeRnzq3X2yAMrU7WsTmS4woscDafy4w/Jy
jJCXTLlWje4ishP3UyiSMHxpmctevlN8cmyHJpCWWp3eDl1h8LCUZnycEsiYqCkn6k46IOxW1kus
ORI0NLjJ5TKG0oBxB2g3nhLTYuFvyoKKMTfC+jf+HhV04DpaupPUMiC8HoZIF3yoe49wTxPCdDOJ
WjBo7GBdMBDlVGsMesTyoZ/XhYCJp44GjYn6l0OX+w+k3PGoHPdXIloI9wZ1hYc29niL2KvQJwbE
xgAlPvyEzD9sgWfUbYJkjSenV60YwsnjOAtJ3wycf+wNstYzXzZGw77VBbCqnPo3zwJmXoHIFZW8
8YFGUvEVq3T5KRHkXp9Yx53vi2t5YcIFuKRXyvjNxXTwkUnGIdzTl3lbpAedSmTvwLmM0KPjrsCc
HSccqFTsiIpK4bQ+gmvdx7niDwiomTzPTucgKMQ3ajmMIny7rp9IcypajsUp6o9Mz8Jmeo+G4Dzz
FChBfkhqkNXgjjacOk5+A/vDoqIX3d3IaXc2LUFkGN7m/6Ppin9bLfllZBFuZM4SkNKOvlYtBAc3
0RlHppjRBGZMUJALoj81IO+ghNUaC/Zh2GGlNbRl3XOoeCuluSSsc57bkIdHvDhC1kJ3LRHDbZBx
yg2vW4FIh9G6OphTa7zT4KpeCl9z4Z9vvoAcoE6ShCV07VYkG+c117+Obg/Fh7u3Jgu6qPGkjLlp
+Gr3HNceHkWM8je/mR9AA3w/WetT7UCtQmR1yoOVQEfAm/BlxMndAS1M3R7EazbVmJZfhYhrWnXv
LU9ETCBh/C9LZYJUrSYEBXnfg5iEVmkBei2LsHY13b0O0SnMO+8Z+Rhh/iT2ghNheSVgqJp6FfLj
1NBIYRrgz16uXLjI5CBpDDxfkCHOmRBDMyjoJAKxaGAD35+hV/aVZj8tMjqyQcIGxW8jNQHTdCmp
EToQvPxtxGXdAzK8o06Hp4eK3UyddyUbwjJIPg3tGo8UwENZSs9sW4aNTDXe2jpRCbGb+Qq4V0v3
ksLkqRtIC5fFkG49D3pVEuFvmUdF/QFvEX5xxqkTx41gDS1XvnoM5vndniqixFK4ai0RgxM+hTz6
2oQ5vUG3Nyf4BbPmIkBXyaBbJajCXUNnKb7cInUPPx5QIBeZjjw+r7Um8bhZr8w2PHPTydPwfnda
ulwPFCmYR29I6xPVY3Iea3GuHVNKINils6MQx1CkCpaFE/fY0aD6w06a2lbLc21swBU/XaGLucBd
YMe9pi46PK4Ut7eoKYAjnbgl2g/IoO6UW0e6O+og+sILzxhXBy+6TihgImQ8oPF5pSisRpO10lRt
/P8B4qXCA66pEzPPfB/X4EfwMGXCTWlSr+Xmzc+XFmxkpSoba4woBW+2ba/ljBlIfYjTBl/ptwW9
Iygof4WaSDE2Ea1oUnMz1j2p6wVRT8t0WhPPhDzZEWacuQZjngXYE2AWvMdj6sL3f8GhkxMxy+Hs
IGVgXfFd56ef2kT8xC+SUkK8X9eg+PWKEvccRAN+6ILpo9VoNKSjaUE6GIfEMGZsXpjXSfGaTc++
Vw45DcDMuG8YgGKv64O5DuP0VG4Ampg+u2IhBVibs6MBoHVyUikedYovsVwghupfaCCzpWMVcy+q
YSrYB2ISvoXvf/1endZ1DmND6zkav8+Sb3yfcOvFAL1jaerSJa2AMhY7Npvl52bfG5KjVdJHzFx3
VwYGvX0b1Lj7KiHR9b+X9fxv13dgQCvZGJEr5YPndTMHzwaIa23pkTeAdt++9mFnLF1ou/T4hKhE
DYkJTjdmDkLq1Avsj/6Fqxxye+LeuFlbC6JQqBjA2zlzwGvsLH2gh/p8IXaA1+53MgsiUa3gwJc9
/fMWrlNjijSggpWCb58dw/CJluVaRpiO8zVliKuBz1se98n2sjJ5TFUFAZbCxAUWkS9qds1kNRNb
bU9y1cijdFluhS+D0uX5sOKpg5pZXezuhkAbN6c9h+KMP6csu4/On973RLR8O9TBi64frECDCrqD
6weLM1J2707w4kRR7B1/Y0YDMsvwqMniiynh/xkT/1hoLQSwjHGnBW7Bdvr7PsWLU+AVOsBIbOr1
O6r+1PyYRxpjSCWeftsNQbnGPIiLB0BN1OioLddtROGaKyqcxpTdTWgqXlrEln//znTLCxpkEQ8N
ndqc8/iQzJPTMhbeHkZEkGbGezxLkdAgRMao8q0R2quUFYGqkA0BdAXWEKH6mwbr+Chwgln4AF7D
3FiRu6opaQrXByEocvd6qAvc5rTVzvcXhZOr8VaoFoNjNd5syFBwo6h3wwZtFMFrdcznkNIWEqbM
1ErpjTHKg+ThaGaBq6QDsbOGqx96WuKzrOWC1TgA54J9fswg7KTFWtCFZwdEilBvLwaTE+Mlqjqz
5vkY81gLamp5gZf1ukYJ3bolzl3n4s3GBqnU95t8iN3cKZ31ZxxN41PjbvG80SoUmNH7alEQH+EB
kxOcmu5+j+Qzq4CIrq8J27j7yTf3uv3kVnCsozJW5YkKHU/AjY+xHiY2U2R9e79Os9S/ERNte2oW
2n28kj9wIY4va2ciZwdXU5fSYhCoEFfypNlNOe72DS96uvAs/t/XdExqUIpn4Ku9vOqRkd8uI3FG
NWqI/F89Fgo7AKPTrUuS5GZ+f+Tiu/PVShMIxTKGZiODIi8SHv8GC+Qt7a3qRcMEFCPqJn/EwiB+
Zj5uG2X+Cmrg5nJeemS6jkXkL9nk8b0roUtGwpntkxt9kG/mSlvjTpTDQ4YefT5PlNoQqNnQi+li
QZA7iIEK+Qi3gX+rea/6ktwbRtkBfI7d4zgigtMokE7SHg5GoUGVX6XNCgm6fhQG26YUJ4JI5WwI
YupokNbFutIpqzrvMwm2aoHcMb1D8pLA2tAN1TnNqzd7Wo18Lx4eb0K9HHkYTu1dtiytfFmKJVwg
qf0mvD5ksLuNECgqD1STzuezCzzv1QoXjbxLCKyQtSONVY37/aro+e8PrGQQGvCkUDyhdtTozx9j
0w/vjxKmkVW27+VEWkNlOIMemo+Y+ljClvrG2W3be+EyBDv4i0oAvNOngGHbJw+fX7GTeLVpOjHU
DmuUcI7X2V5AO7CAlarbUet7q2AmHTIsvLicUA+rqIq2gJvwKu9cS2Xaxc9CIFKnSiZosJVuSscd
ZVkrLNFL4MyG65uksYV0O7DNhOS2bM4tN9m0jqCE5a0AltlnECDZEQLKAyu3Gyu2aYc/rcSiK6Dz
DEqPXjjMEkqrsOuJFTbVnpdENy1L89/VImPUTtPQ7QByhoqKYMP+LqzQdojV9P36l/ng+EPqNIWp
0XCc0sGVgCSv0pbCF9+BOQeWYgiao/R29qZ4i1G42OhCTZAWOZ3D8+6jcVsMrtb3y+qS24J4/vJE
mzldMsCBQh04Y6DQwHfHtS0lKxTPHEjK6v5KaP1bB0MZB1MQoztyZXS4DdOcXE5yfeHvsjozDJw+
k+tiQYGvlzxVE/eH3SKMqnIcav2bHeL/Bsvn3PKn7ajJ6Dhet77AQfWkqSv28befuIL3rUqrtWjv
2mZ38ScFvT1KtfER8PvHMbrf6iYb31eCdGS/7SSNghL1OF3S6OIBlc2co7mqxoa9wZaAmJqovlxI
xWLieQEqOhtf81Dngcncnuhisp15UDUsS4Gvm/GNASfENkb/WK6ojSfMlg6sgd3r6o/LQEicp4tZ
p3BiudgVaDSsJpNWlBtExmZNiK2rKK8GAnwKZl2TtlmGfCsgNdc/oMPwoPDybEW3GLw0jN61ZHnY
TBRVw/tfsGjDsuC7dZ28vZ6vQ3E4RrALVxjv4EtM2ox5ktf1YdpL/9+EoYb8K9LXoFaTnbAIt0r/
GS+jaASnzH2su6A3I9BDupLRodFEoS54h/GO436Sav16+CExotofdIZz7KUb+mIOQGcfdnL/Gkz6
S1VQbMteMeYuDTF/GuoKG1uv1S+dVrRaywanaVPJebGeGhYPKOJxZnQgJPWGkZeocASwQcpQ0i89
zmgnVHxmitUu/bQKsMASae6b/fcOXYmB0OLoF8FKGZg0TxzxIEufpBSH2MUNNdX2kND/ohl4uAvK
+OW9DDcgdwb7SIfG0AszT70oDhOVIo1bkk0VcvDeqw46Ec8YQmukW3mnaisdv/SSRMzpGXrWpIfT
OhjLZzFY0mSPdySK9rkLkPFb8n0J5zW8GvO0UvfCWdfLwJWS8QZ4SYvvx+yAz1NrPZ91P6t4nOXj
LXT03PiSyMxfpfOaRS+pC3oLwZP99atNJE35XhO77qWnqE/h4DL/nuNXRidi1GKKpcG9u+KmRbge
BfFjfFuvtuiorXSnMncTuzsHamU+uNTEvr65F+Hc/s1uhOMMu26FBnNf+6zi6oZGGs6nrvr1vPBu
m4GREF69otfjmTOAJSxaM4DciG9wWDyM97HwV0AXlOp9C0OvqEZIJifGHUmfQTNZtROth9ebIfzw
6O5boI1I9dXR/6XH/cMlsBoo8jcQu2potuXA6KYhrHNmjeM2ZObvAhs9hRwLyNXaDxu/IKNTukiJ
rF523p81NZm1t2FrATbSjzD2OtEonq8Bpo47Aw1uw/iagH3PDrr7ezwQpTZTd4fR1BT2wT97A3+x
4LfcpRjHwtF+g4NSsG9/YmmlaOxsvSqv938IEPbGMsGeX/GSVC8CkEuSRY/e45wicMUG8EY5U5er
nhnrmIg43vMkwUs3V/oEWuNRLGZz16gz0j1hewKzAkoDCfj4l9/2dCo5zqKkl/oQyCeDT9X2t+a4
K87XCgswYymWDsXTq8qovPIc8HW5LyEbA16YA2wbR8TExNe6gBvBxh6z30twDyJwxNMonycQi+S8
7pACZ7tBs8ycaYnPkwQsgz7wZdjrYCkYTVfF40WpNl4s7pSE7+cQFNb0V5G4RL9Ow7UjkTOUZrIP
m314dCjWelavCPABtlwGvhQpuAsf2QxnxNsEQBX9ROxVGQ+GPXUD/R+5DHSn8NUE38qY3KgNU699
X2Q/T+p+Myyn6s/4ahjwSMF9+JIRjm5XMPBJD+UDzFHVrpfuAej/49AOo4qjcL1MkSQhuA7jvYpp
tjwR15yD09FTh4p3JyD3aJb/hEoGNsqG6GgsP7e3RDCaFluuLxNX+4yhhMVErihcNRkYH5E2lOGB
f6Hm6TVD8Sx95NRM2ppHRuO+U0lQ9TGulN0ijSAM0iawzOtCULIhFlm6fO03A1Ba6xsPzTJ0EPQD
6KKjUB9WrzhkOGuA+vca2iG7QJBdcRf/k5aCPj/HMZ9oRu0odE4iWCHw+VXpq2uGZIoX/jElyWAS
QP3ESvZxiYeg67MWskhXZAPOwI781U080Ir7TqfwxJNLOlCGaCLREONj+an4tbCUIEHOL71p1shH
Q4hIHfHoyHdlouZWmwqePV/Hs1hCdNeVVKUbPDpEQuyWwMRX32dEo4N5HtHE/XpxJU218EUT2sdF
CqacLPaDz4vM3usjiskBTN1QzIutG2xpK9PY6jyDLAFvYhMKBGeRAllEq4dL/3v9tNZahXKgxnOr
9bH+YJ4/vZDDa8+xT4cKAzqubzoa4aC0kh3mphu7gbl3B+Nh9e5vK1MqVgmnsfkPy49ErwBb21TC
LP8xIQZoksd0SHpajhYZPtbBr6fsoAWMla5pX0WYBfYBhBz/D7s9lohu+TSCjZwKA/4ypbBf64pG
kePvdaJSUV1FYpMDLvP04k+tZJSZzrebyISBbab+ThJ6tHc5BcrujWFIo8Dba5l89dVmRDxPEcTN
qv//fFPo5XNx8nbi4ChjP8L9/tA3nYHq8gC833tqj/HYkRoyhLTAGiteprz0NAAAwrosTKN697Ae
N7AIa0gto3zSze/MDzaoCwBxgvFGzP12Jf6OKUNH3rUzynvSHH9aaB4pvHybd6zzHz/3Q/wyV9Xk
Ad1eufMcr9ciUigN+jkIpQ5S2cH70SGLhnl8J5s4yDSJUFR9OiARoQc/dQkXx1QN2pUMoHmAZcy7
QulhFRd+oiftxBTIrNO2V5XGNzObC/wjWGiOd8IseiQ66fFrF2ErUR0l2LEaJ0ijqqExn3MkCKmM
W/0JIRZLUgvLxMX1vvuY/RxlW8XHNXsfCMDZfawpeYjU8DcO7ImRLoILm4YPvsvox3lPgMKO8KDX
vyjwh2XTI53a+wJU6eBNjbjnNwJPTdo+ObXzhxxCzgEj1AYvfpESmVgK4R7CVKjgKeqLDOZ6HpIC
4Ei9AWDbcr3Hrnf/ybG8OvauhJulJKHMmhE5kmvxNt5ixLmIoYKA2W9pudmHkIdiMMtsOgrPlQgu
qMdvrEWNjA3qXpvar5lodiKh4/D1TcMhMtZzC0jbxqgvIgE5Ut/HvLVy4W9izac2zZkfCQL/g1qm
GiEnQccnQryDmJupyLWBmLh3hcaoh4na4oZunLiPouGWXUhx0OgZMYgAEbllxEJ24Ee+mtQ8Nbwg
PGT4iZD5c9usAQoOC1/nZQV++9/VhCFUE/wPt+MHrHCdq+Y1GApZQohY8hSKuuNO/4KIAK/jdZUa
tnY2fKBqC+j4iz0WLueckI0ICgVAM5ifG7EvfMqnwreT1Squz72PE3CEQ+5SeQOg7QBaCItMppvN
eUFFueHyLVotpoJk4V5E23BgHTa74IZmntc3zkxdMI30qskHM1cDzARRxcu+IYEfk8j5YarNiqca
aWaBbC2c94P+Mgxf+Vnno8eJfIYHx1O3ZE/y5sF2Q2yAv3DumqSD/eBlVJCNqIeXWWJddC6DBKMo
Q6dHI83XNArCxFYG4+IRz0F1pjKxv/OqFB2Gua3VWG8oN+D5hBxDFQraREYUlv5k9RWkOsg71WcK
sUCQFYoJv8Ib1lmBR5J1IepUL0Y6Vs+jOTtTNfmnVY4bgQ5/FRGhkek7oMsGLRPWfTqmRU4VdSN2
Isd6BZeh9eYOagnL6nPbASaN+Kpn+oj1ZlvA678rE+/N3Lj3V+sxp83rMCqJTvLOOzNoVAnQ5cFF
6dJiyTUYGOS2BrPc/i8ts78OJg+gwZw11VtTPNfydi/HPN8EnuN1Ng3WWpcBGGxij8sfe9fz/luf
i5l/k0m/R4RsSq58cFobRPRtnl1odz4LVSOEjdBHWOeQa1F+1spFwXV3gtLLtgnOkaNrXZKEjavN
uV+vD07Uo4tZxh2DxicGtrrKl9yKrCW96eImc5Y1xYikNbB176XRuq4FxKNSusN/VKCokf+waXdd
ek8f8kfnMnlp2WdXAO98Yd2TbPM1yC2PwUJwBS6hqeJiUgMmy0iHcbUpZTM3b1uJ30pGVCbVoYsW
eXwdFbB4WLrFKrTCGP1lWko4ugfkHItLWBpfaxgD9w4rgp44jGDRNZ+2C4a20jqSVsBGocuJR0SO
pEooRalaVaZDGgwJDbk5REFYcpasZ7+m0fyaqIpU5EtDh1kSUAtm3x2Jz65Im/cEpqlYvIS9DpOa
6sYjV1BO9ULtqN71I9jpgfKleJ7q2W7wB/Ld5z3+r31B7uqtQ05hgy1RZg4S0z6iUhRh+tbpqZ7p
B0BeHLBh+e3xMvYf85ebbmXEVWjDTYfpGeVME5Spd8D0rL9AOJYtRPWoseWgNrxwWvQabOpX2aNd
1NAN7LaiC7YRgncLgY//KromsweT4jCEyDlnZU2k1FT+pgZfNaNptJ0f1iXrE1dKF+gwGIVQtYPp
3wk5z7x+t9q8YuxIs3XrcAuCCpT4vufgOj89+8nd24XUm11BYEptuwTTBQoGZ/JoTV7tyGdbSaY/
f4z3g47swAF/mtwlbxabDjKybgpSle+MUMhmhauetVyhLlXA0T5AfPp00M2Q/Zkiqa5hhSmUmnnP
RpHAB76bmxjc9/ZBaXs0QakSyJ4oUanz+fjysdlDl0cLBoW1fBkVFulBXvH9V3e9dHZr2m1tTjW2
/wn9BM9DWLRmzdPXUWVibEqa+xLv+zaJ+hHbp24gjuDLjACoGdDmOtX1+uTKyPoUrPNU/mYgoPGa
luQt9U3ove31ZI9vH90sRr9OQJNA/jxNbb8Nx1Z7yQH9J5rBS8y9RfRjHR2/RbIPRWIaKyUjaOAu
XMJXS7Gj3uQ46CEduvsioSsBmKR95hybmHDUgB9LG9CqMAvlaoX+v46ADTckjCCPrEVpVaPkXz27
Hh2KL60ujKEXFnL1jiyiDWR8ju1DErp6gbccmHOx1MjrEPM48QFG9jq79RFDOYFa+dr0iBfBl9Z6
EzTiBCLZYH46Uuwb+UpqlaG3RvoSBkEabijg85FFZpNBD5JLVyKZ6jsJ7GFnG6hsr6qOlAhdK1F7
hqH+0oUyY0xF5cP5eelrFLR18sGgWqblRoQTCU/dq8+mj7SzI2WLBpI1isz8WUyyu17qyRZAR9jT
a0hhm2bPQN6oBr+wDoanAdp8yCPrRhfgP8ggJhShXzor+hH7p84RdDNQVLJ0Vef8RNYV5VO7CRrC
Q4p1nK/Q/p43QUObBFbWBgyPGzPJvM+2JV1edrqk5UcpS/4r3GcJL9uxpLPVVbVi/FED6GUbC4GO
PTqyMsOJjGE+KNYTNUxK5T7w+zgaqSQSb9vSSaQvyQR49ht5KVjHt55sQLkqRExYL0qXuDUvW0Qn
xrhUCQc4voUDSUJI6lF4wxzNVP5D2iwcZGWnnT4UG7gc9WIWTayeavGs2ndMfWSUJhppxB41aBBi
IfBek4U1xwFiJl+S+dchLOuZzUVPjfdXHwxhP9MGtQKsA5rto1RyRjjhoyhatDzSQe54/Yg6V3u3
ehhdTCLK5XsgQPacGwkKe17/ax47DHOLc8BrJmouVsZh58LmQVmZNj0oq0dEZrq2+dbDGbI8BkXv
RCIgxrw+VemcVBoTy7HHwPvOVJ+FrskVJyfT2CnwraumsZuWSSkLVrwRgBRX76Fdjnmv+mSuSNqG
uesEHPj2HFk9X++MJUozazoaQfYpDPm+bbgipuyIRhaA4Ba4YrALNpHLIkwtALcswvDZ0U+nAJk+
p1rbwl+57suJwJiuJ4bsS5KbGRTAfhDJN6j03hb66ut4JIC5vL/yOsr8fHCrWIal4DCpkxoQeFbS
o8vQVUzQWJCpnzyQ4cuDe+5ErKz59VQgkWoTd6XJoEPo20nIJabMDMaJ1x7careXXF7mCoXse340
jGUtfkHbNsGbUQAGUYu0iY6tKmHjxkBuIyxtGW+C23Q7WvHNs51+l0RRz0wUWfHWmGrVAZQYpJCY
u+O++ofmDAoDEdbpjbv56l1rWzbFceN5BLuPdj26Ha87fsltIouqE+0u9SKPsbvE9bGjQK8Gn2xT
WTwHL5NLb6wjV/tJCrxDAWKSKyQdKq4cC9wMcHBtfqtXnxf83bo37mrgX5e1uILXGvdPW6Aj6/si
Zsrg3tG/zEL/Q1/KBmOMQ8OM4QK958wHd5LkY+VVXnS6ly/uR9UDWAVqLf+mIBDQGS/kW0U8Y4c7
VbpOzmJRydP7dMrQ5ufaZT6ZTFXozZxL2585omwgrcbDfAA5Xr1n0CBuhe8zT9HpTLYpyvXhGol0
z4hFtMaOUOWG/MveZ4xbDUPjUd/5F0uAuchquZPVS783kzdH7tpF68aRjv0sFpGkneXrU4hzWPP3
qaW3EL0YOPmLe8nygDpU4Py7f8XQkx0M1zplcWnHo064K2jz9TY+0a3I0UT54ufg7lo1NWu4Qj/8
OSUE3HfMAwHabH1W82ckwwMDqOzvViG7QcKsfyKsf3/kqSpslVVbXAxoG/fEZe7SPTRGOxUy3aku
/KfKbgWlIEAzAEXgRq14t1m7LhYhT4p6Ge/GnQoUjW+Bi3gzfXMdxpG6Jhrj5rC6o2TW49whl5wG
3PI92JNfMxpq+gDAwI6THeAN0z7iCT0FTvbfZ1LGJCB5l4pz7c5EIc1vbkvX0PQKIOHbRTUVOiSf
IC6Q6CAdGZ7wYNf/4mgF3Kuqx3fkM5+sBUWgLaRC0blSdt9QZJitGo57mbjdKJDDPQzyLbGFoCX4
frZDs/tf3MKnFOoN+IVkhxPco4LRgLSQsFAW9E1FAbw0XD+9V8MUtVXpqIwsY4xPKdcr9Vm+L8TE
uILSCf5MKpEkW17ywtXyIu5tJ+apVCVzb5nqBDdY3Je7DNtrZMSrg6+n/CUWGzmVpMoyjMvUWz+n
uzx15fLZ8xYlqwUgEdImI49bk/LjUXU6efp1nPvxaZOjMs023Ll8xV3v2JC/XT4i5HPGfUk9TeJ5
fhDEQCYvlTCG2bB3f3Akp3htlGuMz1bNKH/LR5kJSL99dOLYYivxxiEc91x17aruuIK1xw6MUYVy
spSfPCdgmDKuDo0ScPn1K7MDx0cGnt33kg0ohV6VQN7DpFNcFRd5KU5cj6frutwDHV4Ecm5X1Wn/
flCMx5CEnSZ4draPykxvFdloC4+PsECR8GWTfdJ5YRi2rvnADSPvGgyt5Ir142iI6VAlosBkYjVt
gXUb55VC1JC0fBhNr9aJAmeu5wsoS8Lq+tfezax25LUUA+0TnHpkQemuleC/3/1C7Qj2W3qwEFC4
iuR9lR+6n8xteT3oVFu8geLT+XuSVhgIYwXXquVvC/52WCWsMX/9rI1vnoTulVB9U6dHz4dOXM5Q
Uv7h83NDcs4saaw8ClFQLQAXgkYieebIf5vNkHTkWTSOIcPRdyZ0NdgR2WjmEeRbQOLTODabkhQu
vaeeD8QKPQEdd3H0fu5Oy3JUJJmc57Zuzn8HhC+0jaj9kfmNSKTG7eHCiLmR1QxPRWmP7cMZp3UD
0v5vYYkvphMJ6rULFFI3Si3Ieq/wT/CEVLuduNYRsWnxE+xVXuwXvz5R1xKdMb7jIaFuYdQOsqcX
siAZtK+ZPZCw6Fp/ksGTbNxtGqCtcmgErOIKkOC5a7l0L99HxAg8NPV+ifh6NEtVLCXCw0DQWb3N
lPwLFLaFrJSdmMth5jBI0ozmIC0W7bY7CeRfbtR3HusaKvhw97ABluoP09Jap/FKUeqz6todBS9v
spmombl3QDlA6ubwkMd6HKMEYDN20RfB64qi42jTq9sYUgSagFAWbVKJ1QqYzzQZcgwTdAZDkJsI
gTGTaPaxvK9N/52hu/SnXibD3v4LBGO84bHYq5PaIJ7Dp7vkHdanhnvrCz6YgDD77Cb6eiLhX53K
BFPOaRgk4d++Beif52EOKf1qJJLKHtI7xl7UENNr6V56DSA5YOJBCQ35nWCcGlx4S/3fQaBixYyt
TrupErvXfWYBlpOMX91Xs2US6oH11wP6tGeKCo8caIjGDw0F0cy5VXPThirsDPCp1yAp6FGppLFT
c+93UUg/v4r1Nq++S7V1talkt+53B96CQ1k6SWk3B0SbPq3pa9g1u3U9WcXQRgXS40IqADOFBW8d
Vb77TBhhTB/h5hPaUlgz7tW84Ff5EcVY2ZJc8tmh0+PNvU7LzNczWNlvlOyM4HOxsVobcLOrRPi8
0Kq9qjxB6Q8d7gubLvWUjsmDasIa0rZK5u7qPsc3BE2f+bY6OhrW4F++j9N11ro0+w8RShblD8L7
5deF0Ze5FM1zcvY2wjte+SDXDX0kftdubXMnQkvISsIAOeMVdh6jlMTVSCLVzptpqiyBwbgZ2i8j
R3FdN4iuUOkRqnDIeI248b3BYnNXSMIqj/UHTzct5PYxpqwFtFa5F2rWu5EbV5zSJnbaBbbZBqLL
Ywbdz9pLw92zqrLnRG09cor26Nnok+EpY8LTszx6ywfNL91H4V3vM9m34uHT9XTaTZNGbGTAQCdd
xwDzwsp0iyV5jcmAHw+gPqTj5SkGfdKYfAVzwRR4xeAect5bBC/GFSKCwu2ItPlHf/5Z1Uji86tc
oaUqChsqhI6OC8P6At9uvBwaOhf+XZaIEgiTr6IhRw1hvzVfUbaiF50CsEBP4b9CmPLz+AIU/NVp
zFDfrlpgRzvYxlC88poWWPXptm/6NizcEKUg3Qb6tTPyeuFgQ+3EAtTSlCi/KX2CSGs1BMtLCp4v
596w0GLfj/T9tHBpARihcr5628zVDO/SprNKJUHnMOdvWgg+0Nt82Fso3HmkjsZpxyYo50olN14f
TEK9RJ1D6VHB6r1jrtEGiGg6LiuFbAaia7xDK/BJcOWPMSErmu5EAPUvB9u8LlR3PNeCRjckf/Av
BjI21vJ9SzGEqlz6qGWOpzKO5L8uTMV3jQtROkcETs1KRz2m+6bbT80QAegreacAPamA7gVTgwGe
lMxYka1n6pC4k+jgZ+6t6SfoQec440/ojsNTllYsDekp6Q8OtOyVo+lr7mSEzkbo0ec5xS8whYHZ
wlVP6z/4nFRsxCp5nHudDT4rks+9Mk+8OdhgIyDrIdvsFM6Fvyg0kjMi60HNdgcWCqr8ff5VOFAN
mh9KzkBpcOAzS9nTOhi3lW4ffh9bdt+tSB2Nf+qS+X34QaVMzBnZ4MOzSW9L5QzNjkdXXts67I3w
solsh3whPpAB6o80N707NJcgAxxQdI/5Yj5D9T101lGgkpHmcbvgBi05dwGFmKa0aDA7Rf33rGyF
jmJ4pO5Xx2ZieEu6E44P8ztz6wFLfibOFJDhy5zPbD3zaX9OCpXlYCSN2A4swGQ6KoahTbZntzRg
LGNWaLqb3ODlRj8hxA4arWrfccD7oC61xYxIA1R1y4Yrwy+XTIWPpKE8SZvWztpnpaZ5IYxyJRcZ
7z3FcrfwwfZRJQdfoOIDiEvHwSLBsUbPZ3E0qEML2fKALd845qcb6BsXdigLCYSrNiHS3Kz6HlGU
3ToOgCa8Ww3c7qusXBg/7188fnqX70EaKdY0kDxA6jj/IMA4NIeMG5x04e/QSZmFZuyrDZYb+Ijb
rM7R1h02XY9Ux+nszgGOcjUg7U0YAPwu/Qd92vUggTEV73NFf7rzIUXHApXRdBbomyaYfVLRfF8G
4hpN9rWOTYdRnpbYfpRH26NUXPE0zc8ZCQPiPWQKI8HOcT/eAbR/l5rcybzD4i5ZK8KEIQXggsO9
HBWRkYe+wakCwcUfuwhJneh1ZBV6apraPGsvZ2pbpKVZ5wAZJEmqKb29BI1XS/1qurvCwb5OgsI0
0UiDMULOS5lgw/q2Wbpcs1d0qqq7mwJSLWXzAUnXJmGz9aflUtatdCboIWfsebo/svH+qNjSjWaE
iJNaV7XUVxUYo7j5b2KXVrjscvOg3ee54o5o7awExnDZV4r5+hbJKg5tcp/NR19E/Cs1/oo09gI2
wuaseN5c+W92wY4HEHKYr0WT1NjC87B3HP7LvN6KJOCBiod5GgFVLBtf/BCgnYujbWFORw4ALP4l
60qnVRVN5eKkgbPSq2JFjj5lvu0KF3Cy+VAIl/aPrH3902R4k1iPY0DXyWSLbjqzDhpkMxEmrgHR
Cixo5c9sozk5Eyc+5HcMA6wAY0tvPzBOtF5mBNQmmCEwIQnEMrn4tPtYXzkQnZ38xNDtaxY9oTyI
3pYxK4YpnW+DdThcj92ekaKMwhFJzka/aT/IQraISEQi+POKnuKK+XvemCJ246sl+F5SuBd18VN/
ijoZwTc4XgK3vGY3JVVqQwv8bbeRreeXrykiOThkm+CXJXiAREil4jCi9aNnQajyo8KS/mJhpx3t
QJmuObVdJOAYIWr5gWlNsJ5TRhW9I8noRaHAhvQCz4c+W79kt4Hxfg6FERYhZ787kp6GTFhrifF0
cVZF7uPm3ntRNc5RbmxB/gwktOrz+iHo9lk6rbT5NWA4PlVyBrPJ34+ER1hTDqTezN7/ztlhM3QO
Iilv2xV81sHnNyHGeQjU4jKUvjegtnC1/DwYnjlKIeg7n+yKQPigFAl6LKHtXsuTYieu3HgJY/Pk
vn0I5YnM3Bzc92g4MqrUnWmfuC+zHaKaYfxjB0lwo2c0N5/qvfjFdjNyed/Jx+l9MEII8SvPXxjT
BhUzwSW1ng6dk7X/SsEH5bQwVB93Rfya+yiV2ZPtT1A+myvXVDb/cMke3JTZAn/amrg82A9K7b1K
VZVagTxssvpUEzGAU0X6m2iQflxrQtmrykUdLXMvZkXHFzjsY/1TMuS5XCvnBC6U1XlGkL2ACchb
N4GkpXRc1tpEb30bzRA/GHQngRaLGZIJRFpucbpjaWYphCG3qukvQY73cKWLaQuCGk0tGu0s3E+K
N8Nuc4VbscynqC7SIPxeC9aiZQLhw9MHZ44/7FkUy7o4i1ao+/mwKnMCHL1cyl10adiOTGpZT18B
vJEC/4ktqlhDuzchPffxpnaZr578hLZKE56jjBq9kRVJvg1gMeRcWY7pdqcnljATnwyF5Uk4thA4
bJIRDniUMg7/kLXEVM24IJKJCXPhnB/4LdplrzAuKPpu+3YAwLFagXeEfFH7h9V2+fWwwlydLBLZ
p7/yywkXtFkuqkvmBP9NLxLNN4sFDRCE/1qmJnRA5KwWAM7lmtyTvv9eCHhf+Fdnhyqm3dkOAHjW
Y9/SNmtGeLETpp74p8Rn3BkBzY+jnK09T5w0rqr15q3bFBoTfL5fvbAaUdez0F4x016rIX0XPGda
K2tzk3zkReHmZciZeYwag0lkesc2rvlhV8PVkeIpCsmxdcR119J2R4I84hy84NaFCYZJirMMWqcp
CYTc8BlJYOXRKb7tzEuLtfQvbRQhumxfe61iqhH1cwJ2U2W42Y5RlvG5MyuuanR+EbBXVlvfnFGB
1OujVzU+9ncUN3BzcP7I+XetrpsgBnTQWPM9XbF2K5YmDF0Ba0q5Zsm2r0Fje3MR3kf/r+Q2GF85
kxiwwqW1EgrZXvXXDBMbXltQVtBV83EqeNrxGtl79pyxACu2wnLfLL06tmKTh1Omouv/6Abvd3+3
jE61k3rdwbqQBG7gzMmwgyfe2mW0uPBQB+37nWsypStCKFevmC6zBAFQTk4LWAJKw1OYPmcMt36A
Vf6+e+gfwrJve0ua8hsYstMLee8yyBRtdExiZfo2WVlbtMtYCXsXdH3wFKHSUtm3R+HVzNxUloEi
VPZRlHNeuKeC+TNZt0OGDzdFoZOIs/jJB3wJq2Jl/sIr5O2+KOlZXmm8ysVBGkhpaezS/kmYc4GT
w1tD+ysMGzowVHUTRG9pMDOdnp4Yi46xQKuCLTO0I1zUgUg2wcvV8ee3G8RsfPmYHJNYplQAl+KJ
UYckl93UPn7HMMVY1r1GsB3Txvnjj8r/sROXr+6u3KAGYMGld/YR9hBx3SdNFeC7tWwoe4uJxnQP
I/mWuN0ycqhsBxijl6T/o6bIA7p7cm0AIO11biH9UU0WYNbTOTT0lSUFbNoF5dBwcmQeSknMvIJm
OdGzBmN2/HfJXdsEVr+odewXO3cImRsuvWeoTlPFH3kaBfAA0qBPwMTJLMvkuKrwtTG7MMjraNAg
WnUAMyGj0y5XfAHbzLAfSppE3cxJBwNfYoFQscWSS9OoJYoD2JSlIIpqhl+RYgphkm0riVP9PtNc
pXLcOqvirJyNUvZFxO2sVTf2RJJCbzLMVbDMIBlQ2tD42AVsK2j2Ugl8jsH4vKXumfN7Wg8hnTL8
7xW1kP0ONXKgE7AcV8B4URvfvk8syD2hn6hEdq90FwTinJ8PKhunvtqfCvavu+nID6teWjg43/+7
aLrq4kY+g0AxvBUbJ5QIZED0jCavn5Raa8MmySH88vfTlS5gIP+wD9rn/p9sxEU2cwsfPNxQiT4O
kRliOooXhVjgFIgBBJh1ouEusA44z5ohxAlD8t0MnDRTlYprEBHOIkGuTd/I0zrCx78qR0u1UUkv
kVYywlbIQ1yVIaF0PeD5KOJ4UFdtZ5uMhC/cxZqU/MVDVYoVkikhbmgJff32iJ6JYDYtd0W/qfmA
+D5JlXF/Ito93PsuDnNd85w4OaT+6POA7kA9A1/r9jTI/VW+LA9sp27XPGcqNjW/NgZZL5jqiKGL
5Q+oQIU2unXzqRgLXqgL7H4Psf/sJO6akinWGggiRr4Y3N27SWi9CxrzrTbc3DvVXNx/9RLZLPXr
jp2eLQkc2F03Dq7SDaV/wTdLTjnb4RaZ3QZa5ITBS+SDw8WP77tfXMAJz5MEiiIBalKEuTSCe/+c
Iu35NL3q4cATwSgNjJftpVDO7H6Jkffpp+/+MwfVp+DoiOi5ziKG6+ZMkp9uN27YN6TcYGYydELp
2cltVvZ04m3CUH97j4tJ75A3q6c9Ts1RE0iE24ZEWWMDQzCEFJWroeOwGxrxQdLzK7bDuX8UPuBz
GSysRlhv2C1rMsV2krujntpwBC8ABO24zcn/+XhpgOQWJr6xnQURPPsvyeIxOqwUwF93yuuNpJOa
UNvwQ/27sT1TWD+QVgVW4uFY/1dSEmz661CIJ/VSlwtRSDB35GJbxdd6boM7yMx/lszLB81ZZXmj
KhOzkzK+H4K5kQ5LMjmhBKBk0EuPoGv00Fs2kanGn1dA+jhMSRK2Qpvn8YlqmBIA+gk80svpznBE
S7kB1HVJfi5jLH896HLg8iGFYyF/iy5v+3xs4+DmuQu4i+NkzrTiNR2U0Z8r+E+2C4x1+U2dedNO
zyOxctFHRVxTnVpoa6md9F6MkIg5oxkDcdM/VzxkffioV+QShyYHtd2QZh8r3hCDvgBAJ7O9pE9w
pvxodcTBlHObBpS9MnIQIZuJS0CY/ml+1KYJOPm0lOZPIwzGC0ChEEYfm+g5AZW0AT3QUjiMNYKF
WeWima2naMOh7VPEYdnnc3ojou2KsGGMNYAT/HrpdE8XR35fqHNAW5Alal4ZZp8qFXRyAxqpwC5k
ltKL+p5xqXFrC1Lq1yL3UcJX0/b+SpnCw9hlr+JjIdAtNWCIIYbA+ESEeayPfm58Mc1ze8TwVmJK
Fg8huKFV3BVuoQQ4mBHfGJ9JVI47o/koD3OFRBS0k8ZmhStahGaB76swoK2eIUbVWffwSKffPALb
pNIpe9N8FNm79hY/ipFne+eSypdiVWqGrOVA0bI5m2symzUsx5go1iNUN3K1fft+hlWBeDaszjiP
PRHR6C8Fw3tohK2D6GVbNafQBWFLVq92ud+L5HUCurR/vYTmfk7ng3ICiRDw22AVZBNolThuq6NY
4aKtWOH26ZTIvlPC5m2DYNcZjgnLO0/R2TzCJJTqysx4tkrcltEn4FKhFQ83PVnp2ZybN6dGjcPt
4OVjmCZTWiTOWsGgdApfLoJ32vWpCtF4NmBdTb8EoIoSEVdcKSs9JdpM5HBhaiYf1d8AC8YirCy0
BcsJWftSFxODiVQT4zOxaKgJY4YKiLs2ru3rRP6JYWdhxpZVt6RxfPK611g1FkIUP+b1e5LYSDTn
V7hRsWKsW4H7Qf6JSUzhmMYbl8wABgt6mIMIdHxo9VBMV0gWNZ9u6dxnzoo4XgFxQQo/CLuAb6Yu
uFEXncRTuWFii2GOXQswT+sh2riQRrkp8RHeZLWn7kY6IsgrbSDzlUraRBY6IRAIrWcH4KAOLM5x
MJXP1TWGQmY19fv976z3IjnOexhlA+faSxmCEunasWALW8EEcVC0p1qvN7DG7s38p+f/DRi3bFlW
FAGwFsgpslcFJGBH7wyBMQzBQyk9mVUSIgw5quB7M6YoUUCy770jf3Ji5zM+M6pjJ6gZuUvABGHn
yYya1WF5mr7rfVH46DCIvpH7ZQm8/+V8Rc/GmjVSIDSZkpCmpigUJc1HDlmAzeZ0R0HjDeNxgWeW
lQqmpVCyHXlPWVIsrw0ap5fOpBfn5pVYiptGOYF+xNjus26DFzuT6NeulA/VPdwfaGq8w6BYukul
OQyJzLtkGHfbLhAlY3ZDFr27JaaCHBqVsnhHrRlWSvb5rWI7hRpV+Wwbjm64qJY8oS2RSMFDo4N3
yJqv042ZborqPYlhYfpv5OgkrYEODQXjdBoQnfFjCTMt6X1kcBjUxfzm6ReEkQ50HLVe0ndnD/nv
nZKLwFZLtXZvXG1L0oXcoXW68qFY/+ikDQPbMw/1wrssAu9Vshwnk2n/2lszWFgUYHcuhXw1F4j9
Kc8fQHXiNbTkSXlcjTrhR8m6cDVLJDYATq3cOP3fcQK7m1wH+jtBoKdeEBX39Gkr71IXvbtqIuyd
TgwMeLHZtH5Z3A8iPYpiUv9OuWSfY8FNPQPHWwh78Ah8u5DUJI3BnAmTNUPzIFCJV1Mrxzv+J5S8
1F2xYWpQQWYgjo771HeDd9rSYEm1HQq/48PsqdVIwyOA63RM+6lfZf2BeSVRH1fyXJQXAbb8n3O6
JezPa2DWis7CHm15t06rjnEF1J3NJtUheAmv5NTh9QUtmnggDrsGMsdTMQEwINYUMgZQwMscCq9T
dO+S79ZDvXgRNeOrX60fkeEZF/A5KrVFE18X7TEgOy7NDMwV3lMHPQQb8Fog6f0qB0IOaXhhwT4R
Hz7QoL37dBJRJwsCdA2wg2/hLFbrnOL00wI4+n3NYCwSzIe7YQG2pWQi2jOdN0ZHm2oPoPQcElRO
eyPuLQJvtD7iRNZWqI9y3l4+lQKiJPLxyAJ+LpWlg15db4KX+5Z8iRGxfm5tR6ixKIUdv9i9LmWD
fo4vK8wBErWZAZxGDFEi9FvgBhxTcOL8UJVGY4GTatVWX0Lxe06a5IPsjB41ZawnHfD5rubuKhXy
yYNQTyKxOCrnFhaq5bapSyquMKOSR41KOOhT/p8/QjuWvjdNMOiRtG4FUI+YHX8FncWL/CXTdSEt
YtrQip6bgW2BYnWdYiJteYAqoa1VOgV+NFal6aB2rkJN4ZEFyBUOhg4ttWiLE+jIZXZDVZt3I8bG
OM176cxCIydjOGA6q3L+wkTwJbObtoW2HoZVoxUMkaMk6ymJYQWVnL1x9jZ3OBk6MnHwtRnV8CT0
Q7Qv6or8x+wEPEE9mhlm/O/2b11Ix8heQawLeVIDwJc0+pGHkyZfJ5IBDcwt7OUjtrPyWsMXw/0R
gztzq5koe3Lmn4/foRqLeL1TITApskbukB62/aiPDuguwerAsX/fggn3PfPPTskVjFH8xk67etNm
THvLQiPcka3szFqSSkjmchYqzB7KZd5K0yqDDeejSjFNdaGJ1ZprCiDVOwcys3KJb16D6zpOl9s9
rJJ0+wfOk6iHlk8f9j9ObYjDL5/y7GvH6f3kaR5vQWv4OENyEG/rHOMYNrU3acLs6EkkTjSPSKax
lemefknFKej/UIKwWJH1CcYA8jQ8qhrimCI8kZp9LyVJL3GVSc4O7rEFYKfSB8vJUE/612TEuAtO
hAkWzeH6NDkmWUT3uTMCkPmenGvpIbpo2618LJI4emMzVpuHwGaHrd81yUhbWOwJYQn/iySYLWzI
taoEDieLJZBDipTYdiKjphfsgLbeDEvCjFRrcGZKAVjavPAwH0LqWkPAiMrN2dgZC5SXSRFpZfXJ
Puy7w8BBP+M+fO7spvGqp6EQ/4QIe7HZKirPx0aFee0BaxqqpjaYwbwx0am3solOl2jn0B3eo2ZR
TETKgTrIo0uFY2c0H+BVy5H5Qg2Lzm/sxVoPv9TNjDmqjO2wi1yo86xG8FfMSoWtK6pwR7BJxCGw
/86JDxFEp4ZIyJdVwNZFdUNIeWzvoghMou+DYlh2fet9YuQuuPC79+5BBLA6mdTxq/8JHQqGYSkU
j3ZNsUfjy5imUky/mxW6XTbyPNPhLDL2cgvquInHHJtAm9KuV3Dsd8yM9l5YKi++dV6EcqAkT0rf
cB9eNaB9ob8838CNWHKf8mZwHzIIMWO+qnWkL0h2elpSo8T42urOQukYfX+7e+Cg64/VayHHfUBJ
nTvVp57S7DRBzQ4LV8Va2lAPK1Vk24xnqhGfjdN0gX6gYWS2rChnPBQd9kvJW/KoqpMwL+18Eak5
yIpwy3EVI95Xs3daiLZoCnJcVzXLCxOVXc10vv+iacnLsV+n96BGrI4qQjEqOJ1WEKo9SHZnjvUR
Fp5jmVN9kbljTEt9EGjSKkFv/xZtOdYj9kDwldQFOMoeHXk2JD39gBmTjS2lvECLbf5zQ1phDoXV
uKnh1l2EkM5OA5ZdXjXGUs8jOZIwKw+Gspx4l6FO5R/VE0FMSiCmp5ERZu54ntz7WrDHjhFsluEb
jimzluVtmU7K1tfpIt1iihsfYcuSP098N7mHzSldE2yUsOGl1JKUenYO75XFyrNsVyxEcE/21FP9
2pVcuK6UZlVxj9/fqXRfK5h5zEdwLEYhck3HrnPBy/EY/IoybbFVfVwtgJxE5PHsLgBWi+PeCwDJ
7TUweHCVgbXcDr9whzUNLbYDRbD5TdnKGTGWPVUWFqv6BpdOSd2y0uzF7k3+wEHmQN7l7EX1O+q5
J12lxNntma9Niz8wXuWUfDzu2O8sWryTXBftcSUnYZzB/LNsfeMaEIf5ZVaHBVjtRGlKnXzi7/YN
8yutYxqDLlpy4OjKtYzO6RinwCrYHphUt3GpxPU4atRfuW2+NO+Z2a+EtVUDZVEOOPE4UfNUUqD1
BbALHQOgfB6tmUVcJVfN3orChjEaBCEo3WXtqoUhPdZRTvQIuW5KPT7znP2+Gnfk+HKr/9bMUgqw
GTBL4eGOrGHvJ8IXXnOIWuuX8H9HiVc3FKqW/4Rbm/4pUof93NT1ZmgInR7jbyR3Id/swFjlOTu9
Tpf7fJ4iq69MGynqg7e4woovd7orFSXKxcff4kEEUsYt4QY8EhHChI+2qPLSMO1YlP//ckTryOBk
n4UKj83EfBoBfD5cAqKx9buKV6y7hlLnrTGN6lczyI4cIuDsP60vxXqVm5EFwTmBr1I/H16weY48
NJzuuFXPUb42Od5t8Tw9sQvVvpaC5ggTxYYy5WBic0nRpG8yTiEeLimvu5wp7eAFbg8YRmZbr6x8
Oiw8Tm1MaEc/Ud7DtLA+BLRg4T+PU9PXbORA+6rG0DUH+XXlmZgDJiAIpNdvew/YXMgS/f8+2ZTD
JRTfPRX8jorwe/3u7UdkgVjlknaZDZTeHeiSUl5cgQWy2bHO+Fyxw4Ef7H9wQ7v1IqjBQQTrvqTc
lqMigtd5eZkLfBS3bAQRh4/Dc25hzdlC0dGLBtzkCbh/c3ZpOoI72eUuvP9O0i/1Qnwov7UtQ/iB
oX9ooloQo70Et3o8UmClLOdRLx3G5hZM445Q5Oa7PVQO/ggAsH6rwos/QCXPJpNstXg0GJTCPxfk
MnKqp9S31+PTruknxXoteuaq2V+ICei2BVj9mDZfqxS5rFSUBQT20/IzIt7gdWsbWbjykyKXP+pH
CNNC7E4SB95Vp/AV5/3Jqm45+aUwQtnbsDvAwyoTHv0Ex6wbL2IPN/Wtfwh0uBg002peYwzMHIIK
Hg0PLv6AVFo+pGsBG5t/DjnH2ZecPfV17NiIFkjTwftxfnlaEjVpAKJq9ElNwll0I0kVKerT9j0g
jM98+ekn9qsA2wFxpCuh0M28fvoRZfVcq9MdRNnAvtREeZLuoNHfB8tQgxtNCySZLhp30HurNUg2
sS9plxXxctjP3o9AamQWjf8yl75wYIGAw5QadZ6wPVFbQpL1kTiHvas+C4U6WQ8V6fK+3rno7EnI
WWGbQdyBK21AT0AnHj/hNqskehgwXIpSbKSS0SbcPFBCOjXvpKQcjWpXPEys22X6f0G+KQBcP36o
EOn5mpKNiOh2ynGZYNU0zUEpGJtDx1+tkxokagchEde8VvRqzG9PwkHJz7NJXUZSKeQPJDZVC8vN
saR+MdjxYbk2bEuzF63SzkoUE2MvMRLOiVBNazYWCGB1J5Fy/r0qb3kzvRd1k58rD/53J/RTYBp4
N/BA0vnn/o/xRYApvfcCUzzAZFPJ/l+uL3ZJOOChFwm+/YZbr59zd+i/qHBM3utRB5sWm1OUjS4N
1f8VOCBC6cOvDNCMgDdCCS0Cvqnubtm9ZcbSl7OMl/L0EI44RS3oHukc2ctpriFDACDpl2N07lHZ
WFMyAfsRZ0ipCr7UPOTggGFUQY0W2dzCUiJfFL6BP8yxELSVPFrXz6JmG98+uR+FMID9puskS9R9
112/0Mu3fq2JkLn1tD2O+bHRB6iaNi6ACWITvyOa1WY1pB2suWQ1sEC5474OgogjpEn0C0lzv6x+
xmH8xlMV+ca4GlGyodMcBMzJqZ1TKHDLrcE/WhyB52mC3pVMBbsLMIqFUlTSgwhAeWhLzx5JJSnG
9HYIjje5LbaPxsvH2snK1Mkokf8zAZLENl+7iw9khy9K3oJK6fX47bXgwe2D0D1B3e6DcHDBWhGZ
f3g5yFJpRRG/rXsLm+xA4rlzwaGhrSVywPya04VJ0CJ1fMZbGQaSEavi8eJ7SIXS+eKZHLBhNNk4
YO7+HKw29bVgsQnlTXVQAgYL99v9VtBXoatCXcvIfYFiwWw7UTO1TeWu39MHf4kXb6Uo5VrAlQW2
24IjsCpqsbTvJAh33V+0fWhP6USUxqgcfjd2wEQ19jLTFod1AcL3MPNF4LYCwrIXXLyIjZPiQjdE
x9C+1no6MLoymDqLxFbwQtUFDg8XJqfvlcZ9zt3tW9/eQ3E3pz/qkDKaTgZNepsUY+gYhzifk6FO
/eLIpq1tsmGa+sbiLlIodblG9CXpHxdF34+gdbVSHXnuM8nb4xrsdsgsA1hiCDXivgizK6xYzNFg
MvjzT7Fa2HR3J9PsOT70jItkyv2K6MiCFM2Kdq6HwEkQ6MA+2k6QqLWLC1Jj3WcX/npEbOrsO0QM
KUwkP3o2MrgNM492Jyh4somj9RP4scQyMQgBwmdanJdJT44/NlL4RTVwuyd6PwqNrQzRDlcXydOB
D+B7t44llGTxFpd1uMzvNpHsH922DWw9pWpSDLiIOndzo1/74NvHjxT4gRujJLVtlegIjgVNittv
ypjl1r3ATKrcDwESs7ZjirRauUfG1OklU6BK7k6sVMjEKm1vx2+ttZ3P5eIwEq9ytQ+m4mo2+w0v
sIO9M283Wav+QQ6MqLd46w11/tcvRpLdvsLQ63GuXVvacvjXn+guYY3T8RQyDuN8IPBbmdfBjPj5
FhJiZ5FHY19B/w3tmK2P/CvJ1JS3AGhv/oTv3mESmMJBkxlmBzhqzr6n1gqRfXspALRbwFD3kJpT
8++fzDhm9aYEuzIqvc0a6ulh36F4c+vfYrbyjTIUTaTtpW2owXVlkzKiy8Dr0lz9KoY0t1QtTJkY
6NqUKRcFI1kYFMzEMP4xv+KHqavE0TVaUvZpOenjxNAHxErvkqNCjZCtttfnEHKuWh2o3exQ9SNg
P6S2i4v307GnNBcmmLqLN9qA8NqIXYHEIu2C0pmhou5yGtn2NXnxtTsNTJLaD9v94nBU5/9RwUx/
XR4H6+BFcYFg764jQNTxDuHJMFUmZZuL+SnfPfBZsXhEnaOt0JOu4ylA6GAWS7H8GxDH/WA5injW
NGkqUEsea+abk5SeTFRaaMspQDxPHHULv7hqec9Fw5jJmXs9cDwhLqP/OK69CEThyeM0+dx2fQps
1g7Ao4LoTvV/bqfTRDdAXAEdQknN6qDLc/Suax6qqMpzmu9am6yJjTW71dI5nGJTQcLskNlkAC9a
ws8XtomQwvJT/TPszb4NymSl9R2qf4DaTGYK2IHL7fIZ2ATip/9JVuZkIylVNMobrC1R8kexJ+V8
bHJirKAG3CpWetHLIzC/pvl0EyKelWNoB/PDp1WrAmiXuR04SNRBw6lFaYFxi3eRI35qafUPi2Jc
qwIF8n0W1LAcjdPe24N8FiIC3BqXlG0K7b51RmpxSB6+rvi8wP+vrhOcb47c4zwP0WfR9wXNQTmJ
Qbew98p4B7Nnsf6fXptAfbjxL6GdSzNFqve7Bcl0+hZvPf36AnJE0VHOziHgGV74Qo9lqHZbVxBB
slOfmsQwPiXdzC0GDPHXk3rxRapvodP8bcuMsGG5TnwB+DQKrkaaG6HtRV5k8jdJ4C+q3D7YC9V9
PIyQxPBeFB1wbni+rVnpc1WAwjxW/dgHeB14upaoe3gf1BVTcGlK020rLXxaoyZpkuShWqrj76sz
M4JGATWq5+07ECe9dIEMhCKlFD4YwXpJo5PUIJouN//1bIepnvWA3PERRYqUnzA6dV5ktCoyA13j
ntdexokaLuzWLyBYulUKWxBK3mJplEiYVK+RRkmGDf/rL1HG19A2q4JYu4Q9JKrENhsczENbXFRg
m0XBPpYk+QMPlb/lZoqnna10UwsWVQ5wXDrHNlM8P+wlxavTP5CVB7E5IHvv7G3VpqzHVmo8gg9S
wsMxsVsBZjckhYTkPrDRlriWBbHQK+tA7P4JN5rom3E8s12BKkfmGE+/zQbDBXKM2wN2DQ39FoDT
8h1QjK/R/tQyTk6+66Qce18AP7YLM0lNCd+SjBZwhfJkXpQsiQ54WT6XYgdUpgLvSUKxjdDwGmCu
L6tnJUTGA7P4uLDqeK+waZyArSPIkDNudF72eO/inMhUWiKQ5CnH18BBlGMSYbYzwuBqjDQ4twB0
fbmSq4zCm2g0XIZDW0YUpJczpBeDnXKcG0+E9cEDjqSgpJVhHXRmUL488jXfzrYbdtqzF9bhJFXo
/5s8jRA3q0NgU3Ge+b+kkbzMSh9GQNAwEvTINCeB7wP640qX7W7TFhApQvUVrMhZj3OEOcJ2bD9T
soPOn2MmaTjfImkh6++H4xwoP7zLcIb+gXySCHYMEPlBzFbDxZBibZIqL6Mifmp/YgOAdf6iDgwV
XDOm/7ceRtUZr9faHBMxDjKsEV9b+lHVBgg7YvA2e7ml6uwZFC5Kd65qc0QIQr9GLJuUx6ximbFh
pqL2R5QqiBTcCERKVZfB69mIPH6K64EpkzEO2QhvkMTMcbsdj9sEjxMeyz55TCu/WdHAuEt/iGph
b3iKKFPqprRHGH/ra228STlevgjUVMdz+Iv1l+Grx8NpOo0SD4Okm8a7q2NmlEsZ5AfCyvvVFW5v
XcJRc85/lOQGOLDFefgsdWQb6lRAoWCbe6HZYOAYYge1ZUMYdorUEhSOkW49wZ5Tm52K4pdlpMcq
/LwDoXEgP6XjpkgXv/wnZrA+QU3KyiKiB0V5Q/6Mla9GlD6YVJTNPGVQl3Q+1yFYsysy1CEzxB74
uJEfPLPQqYPb3yqvb0YV+h5VH+MSjzffg30EkZ/1m4dTDcOrgT3UDtumQIVvYDwA4UUnxkh+UejB
uCZfSPIdFazlhpYNWaH9mckpMituK7c3gd0OEGdQLv7RDhH722Vljzv7egn4VhNyR5WClGdxKLBM
lCAVGFx3VF2P5cIEPHpvyoWu8LGPH2CJHa47tl3k/YS3m/Eyi1gJhYTjhNCSPcuHi/IMPZpGk3Xd
Y++9asRI4/4QLIbLWuF0YqtOUDXITav9UDdrscTULvlchN3q5Bxd/hZ58RfTtCwkJj8l/oQcKNju
kiCN09yoUbq/TpcNvlCVnYtJDz8MTbgO10FsE2APGUatUsezvd7ludn6aYQbkFy00Udoe6R8TNaB
1yDUv4IlUA/BsEMKDXZwLIRt1n2T2wjUteGJdcdwsdlZDPBAFYwGWM0jma2aR6fTKKyDK/md2863
k8NuWoxYWQujMQLsRSZrikpTXQR3aCxPRc6a6Ey63PShgKIsCtW3BBF6FCiHSDN+l0l8HJBkDQ9P
T5dIq5bdfgX4Anbcw/WuwcHWFAd8xvKPyglVwuzVfcYnkRjRb/ST60UttTzc/7m8MnjBNLdNe4kj
R8cL6iZ8oYFfHzq0+s8pUH2c8OinmQONZyJkLrcESa4ZXmuOY2c//xwaT3RNVOSqg8ChO/7NXKqb
zZMCPaAd/3Y7QdLug5zhdiqqfrNxJ3IULlRKr6PuPUcDBTaFvTzZ3s1vlPpb/S1neJbXegD5FPwF
+J+n2xjSNjLYv5T0J+VWhGIG86+b/UnVp08BF700CMqHSUa08MEWdnqMC4/gy1d9yXsfr1pVEbyc
xkdP1Jjpoo9TRGcNY7lECgbAm2YZ2NMKiY+0WMNlO+nOzcgmlJgQKb57JQ28695koPR1Yfr13V1N
K5GIKMOvZmS1oowQ0HdASoLUPIoGBNm1HGT5QwIjaTwAf/OuSDtLNciVjwvZpJAYJ1SwtvYefUHK
ZhAQeeEApLtGL+iB5JAipsR6o76BwWsh8U9gcO5JNuWICI3u9eyvgESTtPVYDqu6n8raBldXP9vX
/Zp2BoqHw2GOfZZ0KQZEfxwT5Kcbn6DmQm93P6bG/imOgDg8H9wjdHx8JGpbIKft+x5f1xHQ6XDr
3uvmw2atTqAobOcZ6h+hw8e8xtibFBgFHeKNimprPRJnNKZhYkQiCF1qox9Ml2ogrFPftuKnmY7H
zC0ZBBxg6yaoRhROBdzZ9/aXZFkZfaTdQGiJ3EypkEoX7egEyhJSniGRtCBu1djz0TPSpveppPNv
Fj5TYCYbpGhnpGTLT93ZjjY5x9fHH71Ez9FbHQqs80UlOcu7Z9/N4quC3cF6cMMOH+5pjHqx5yCu
qoT7nKdKf7XEvInbjNeJaFaE/KjTu9Bbz7wa53SMBygmnQTA3R1AsniIfrwHtArR4fXd2w5avsOy
8o4BgvQOA5tigg2DVoShPvWe90dN3LH0JvSUm+7W88C1s3f39+VLCAgyrpUKCwqUXBGiVQmwtByi
b8F8zekiK14/cUddzlyxRSgS7Wr3usTX1MYl2tH/wRhGq4OmfeB4+SoQ2dwhGB+m/XBVFZof84zR
Wk7xUWlhicCOCB592lka1WcPjIX2L1rU1tqxNU1Tx4YnZF+487aYENVIf4MdrFB9HDTz+CbjuLzH
rtSSzA8Am1cXOVivBIsdg1RL8Vwm+Q4BFoaGkUbnr1eDy6p9mUzi7tBcVwWSJADBkz5ayxRg3mKs
b6POzyvKGmrommFQ58EppVi0FMiJiHnYKIuLsfyGjMrGEE1uYbAzY+4sLD8qRO3neEM3iLxIpU2P
c7LsDo+9K1QCwc80aHZhivBvH1NbobmeLL1vaTgJkAkFZ2T+YJRV9LkOTYlV6VIOGohwzHH3BhHG
ZzNMqCHr4JZpEVmBkCcD8XH1bDVnXdr+6QbHRMjRjM5JcrOb6HTrcBwue8PteE67+AhkxljAspDJ
wvm/b1KmlwBO0dC0SzRew9dM2LXw1XxNtiJkw6KOvHpV/DG2SFfavGjqfNuxrg5aaBnvPfwYv5o7
YQhcyoScNiPgssyFr4nYUXUDr4DGP9lk1b6rQj+sHGnoog7+MhkCrmgocNbgxwj4/whD1hcKaMKD
WXO2j+TBlFsG7DOg13rufnPdUsJO+f8icmlCq93pMvz90It5z2HurrODxgKWVOsNyKvzVpgBzNLL
hoyXr17RTN+VF9AuZlaZrB14gRqSrD5jKhL4OzBuc7kBvWngIOuG+nziG4SMoX2IrNLu6Wbb8lZu
AfxqALy/bUoV4WPRxcinLUyDZ11B6em71uWG78AOeSMmoBX7Tn5Rg063A8Lol39Ag16Skho6bN9D
0pzg+Kd6tfCH92gWtQ+WMhkZLLPPaNS/aWwmb5rWY1zSdNHSpTawDpXWvOcDkt0pKr/PGN/HVGGu
+h+QPjdPvis77X6ahgMhtRpKe7hpxIZfb/kftkzE05x8hthISzaBZ9mH2SB8uPTNikq7E4u1zqkz
LZBN1cilxRaSuO+dNjKLkxZEC5x/2VAw1rxQ7lcNnhJhkz+wwEyzRn9AvUjaKI8Q84JJPihpra64
ZC6tWwmKVjrnBfyIT8Eqt3IUHNnr7oVnLvxv13Bt68hHk6/EYwB4EN9ZReGkvaW+Hgc7rlH9xzT7
1NcwpKFI9o1522UIaEpfG0/+BJuBmJKwYHZvR1X6zS14nq3KWp3LvQrRUxowy747mIx4esVtCm9T
pD8es7Gg2Viu/NtEsKbDKANhMNg8sNOKLynIi9arqwSM+fvJFimJn1cWRQyXz7aDo1cjGqhmKQgz
zz+dmVv5ubUZueTCStqogTigMOOP7b0gdxm2HRXPmNRbv9YAHK7ajIH9DFfsWgKS2TtFovdPne7D
KVzq3aRi21FEAcGb99rxUSLC6iSSIP6wES2WMnjuzdLqdR1TacFbxl5NAGNQcVAGOu8sZdjP9hzU
U3Bjnlr+W1rjQ7Fv7s8qjRfmgk+q4sNu04rj70F4QzD2rHSoUI3DKqOCjc4G5B19LBy64gLx0B5Z
IIcRa7JyPkvNHjS4K1oHV/Cju7qdaXo9TZiESnacaCFN7daJe2PisRqW+FNWSMTc79xN0q2/mmHA
1bhpZzI2669DTsFQNyhbRbDMhIPqiFzKEA4VR2ka+EEhLcDM2J2kdaXAxCnRVG8oMC2Epu5HC429
EMpy+5MPZd7h6N7ZdPWT0X5qdZCTJ/mVKzmTSXRN5RX1x0xBCjTIN1inngfvf2zALDQLpJkrUDpD
zVyp3hXKtUfSoik4Qo33+cH0x9KIpUVAhpbA0TWU8YNPGaINW7J4JEOEqiXTC8SkMuLgmiRRqgwl
lCxsc7hiMWWeaXMjq8wdViWb4k0qsVnmSLc2ZmT/fmjnDBtJt01s16QEzKpzkny3eUcqnuhbveLp
18upUmN47AO3dNUT9mzrKiAMXUYqRI5w4JrngKdYFTe9b4UHhYdhp469xwPmHx0dz9OcHhZHLu8e
f8cCX7r/pBYBpF8lRQZsl4+CC22Qt9J6SsA+EteygjUDQZVJeN3aF3L4+68+dH1rjmD4rHFP1j/V
DxRg52RmOkNHJDOvC492C0Ms9eBAJdtvoIeHdNo+UhWquDz008GploKVxWvI+cDCft/wsnFqRklm
3L1AIAN4R8iJkl7w+XoyLpn0NpmeFVwUmcyIjYRd1P51ZvzCeZVjDeDxm6flRUWhiCGxGGDHOKiD
yc00yQ1OvNVcpN4s2VMxjgQyvGb2VkkbQm8WGw5D+YkVyVtwCTgMO24quFoft17Eiu2iubcEOUPw
owmB1avcIFLq+tqKcHlExBqwRopeAEohS2XBiDCObZ1BYDMEJAR0WFVRjKI6HwGCH4CMBaXKIjYu
CXxaTTs8/HgIqbVVeO6XRYBs+5bEVvMoQgA6cESTX0ZjPxF75rB3HqAQ29dhN64pMV2k7XljWPOL
TCSfWTXie4E91pKcy2Z4j/bljoKU66IREWDd+bYO0oNOB9fRXrqXrPr/2ZwgaNwrbiMbNKvir8TF
XxK+QbIRee26MThrIjUPZAk6LJ2+Y1o5e72AI3RNrzcz4jU59SejfxC/4l22FZoLW73MU+0CcBEh
Os3hLbh2x6SvjiibmfkGTPWY/m68MzORe1KsXIepzO2UZSFlcn6X3THFeNg9UVa5Ey5veJxGWUvl
VOL1p5FKprkahBCC6XDmuzwHDKv7smZfPy6rbjfQBMkKROxFVWRgiM8rMTYpjVVZ7Gzf0KedzAf0
rwdcQHogHISPIlI2tYkiO0BHFu2NyK6xAP7LmV41GQWWmHX0UlTtpMj1S3VTezH7uQpYYgQelzo5
M9xm4Bb6nCsXBq2JoIZjVsAMfICsgZy4ZuFDPs2bBhFETf9GjMhoX5yjrYYxXzq6TZWyRskBjVY4
jBjQzwhXRjkU7HEKl5wPN79eCAeqgInE2kPf3OvsztjW52TNlS7ehKd0kD6I6hO62XFwhqNmkVcx
Q/c6+G5QqUh8CKwy+OXQRMqfHcoFGqzMm0HvPEa5cTN0MhjEgpgVE2rD6lIYSqukQReAcEzLZMTx
qHdljWwNUvLqFgFC+xA3RTKXBC5CL81Ys/MU+bK/iyQn7jkzoKtCeQy40keP+wkRFtgTw2tbr6K9
XGKRnkX/aIekUTQ5/CpDzi1wUnrkpddDgAQspGKREAd72uSiZAljFuW+s9RfgbcSYsBbn/upLW2K
qsdmPfkX7uvo/9/BzqIfSoAInegelGgd1PDnuom23fZEl7k1enpXOoHVjRlsNW935BZvvrbgnMgr
a8mP4KpfPXXA1Jtbu8Y0Rx8xzLH8wkndqiatJWoue6VqOgW+mICrgXJOu66E+7yAafmNqJgkkoiw
60MYGUzrQa69JrwTYFGkDepc8aKJmBkz8WcAcjxS5O7YJpKWPlbc77GtMIZOt5b4+/KyDg5sED64
0gJJrv5LCRlHbYha1TZoQ9Lh1j0V//UHPexV38ncQjhgOa6Rt0qK2s9S6Jzah5ZOc8icP8extLmr
FDEGQeQSs/dwmxUtBHFpPTIxWBX6ak5ew8wlRv99vJeMVqg924qJMU0eE2EcmROV9nJ+ZAt+pegc
UPRD0es6jYlvir+5VshCH7lNsIn3Rf6A/2Q1h6DWdCroTzcJOd6wS3k4uIsIlAfr5PES89oF3Z6I
MIvSl27S/G1SRPKaiXR2T+gxsSBrFu9Ef1P5LOOslaM6Vs0qsjNRFt3CHx+dz+Lysm4/RznDws13
DjyBVueFI+ksWzGicLARXyvXq1MAeDmZKMr9nIDCtVSkhhaHxYG/x8kJsTEREGiuTeQ3TrLg3fZ/
xEgcWwgSk/xYUotKxcMR/hClU7aaygxcGLJefHp9Ign8Tsn9DR3CrWG/Kwc623FlueWFHTlkCkfm
6byJGxnU2QdLVQU2DENGWU4QURwlpo2ReRmU9ypkMl+4xBKeK5iGX+0Rj1je3Qb8HkjMMa+1zgFp
gduANeCuMTg8TV31XD4lygVMECjNCM6c/U8kKuRRz6vCVaYHmlBc+3hvNZ67YeHwR9Or3HIPwpbk
eSiQuE/h5Rp7Jdlk/a/fOSgWBG/z0hxYBipZpByIuadwOq935eVsKDtxbGtTmXE+RtAOoNE3YapM
npt0Tvl5869ZP4oL+CYCVb9WOSAq4XplLE2F51jTTZbaf5baGnPCO0u3SmWqkAPYxQbctYgnRIV6
17rXBsQPHwxLQMpMeHSKS6DlZrFlX6cQ4MPSmV4hVZMV6EyH5hskgXpVxQWf8FfFvFLsOPC5qck7
tz2brl8mpmsKxKtBzdpo3anW3P1iJrRvn96O1RwybFCSlcmIyKm00DSxrqZjnDA98VNpEDJz/yq4
aX+FXSxbtuipDsJheR4N1vgZMf4VLYqHAsbZyOxN1u2nnFPTKfjFkjUZ1FwVb9/00nszRQ5PTcHU
CCN5zndPVjqe9UFeqZgSt4fYI0/OqKQhOZLBwIfo/Fht28eMWqREkHFRKHpvuS5/s1Is4tmhv308
p0ZcP7Govlb6YOlv35+WaA1VLAv3AlzKU0NgbSH6X03C4PAS5YWXPutrdD1Wau1C5PeA6YzRvovD
MXnv3XF26+AcsUzCIdu8+p9gRAtVliP2+LvU/Vkte6RuLvNj0gKb3ucxxWqbGfHqOIVuLVVDiOKX
Le6XOAsDVrjJR+5GN9TYRzEyvvllmJNystHsCaLcMTSdtqRj5uBNNoYykwaEqh830f/2Kv8PqvJs
W9978n4tCZv7W7do3d1MdwyBdtEvwPFRwjTAXfVNm60rtscDMs67GdE8KXDZfl+g1dch2TmhaGXX
p9i6lNWcL2xIc3CeJ0pO6EmaU2ct7q8EdoNrA8KUUsse/gGG9N3hXVz1tDSzuUnSUlUqMupuqigg
ERpE6Zy65tonc6PN7eVC5h6FDlvZ3KzgZIHJsC1A/1Wm8El7cPGmUnwwmBmKncwTod4MEyw5wVkh
w9l2V65wBz4/JjfXJLtUpZnkivhl7DyR4yXEu+sgtGeoW46TddlHXC8Wt8FGo72Z+bWDSKtfYT60
ODn1+mIbDxgbU+eT5oTNbDTVAKb9ZK/fHw/Til/nAMMcEPGD31P+u63JdS7U7hP9qB9jX0Jpa/F0
84jLI57245gzKyramIR+FiOO7RULePg50iiJETJYD7Vp1lAewzXqFYRF3LbXXQvFdbTo0urguuZe
DRqlxek7PJYk0B+uGztjSpYOAV7ITTd1HGJ+CxB2Vh6q6ciwmPNX+Z6wDjDQpajfqmRA79jnP5jr
xj6+zFls3+ZRCDPl15akol03rpiQpzc7jTyn7liLD7ZDQRNjYZjiECW1lXekUX3CwOYxQCvLQKMV
N2ojE7C0YM6D8VFdViewbfezM+BVFbEAdNIzzbOhEJxHzEN0mx6WHoV1njH5LbBYYbJPtL/+pX3P
S6re/4DBDGA2OkyeuCeEERXXDg4wSEQc4ciPXQy1cy8cHiLTq2N6jlTD163yYu+7qgGinN+0vFRu
2RRgyKK3SViwisq3Qe0AAENS0jQmlPfBlAj6cvd098WRrYUlEqI6fxC5zPUk9Th1WnGawhVTdwfs
R9DcECPTp0SIeeJdMTKWyHbtwzIHRhoR0gWpmR2th3xGxCMvrmNYfyyrt9p+kuxyALxHBeuWdfxb
K6/5fJmDIATwPPX9ifT0NVBlMpwDHssC1/Cfv19i0LwRdhGEivC3phB2FpYnzgbAr42OmBm/JGMG
3Act0GzeZ+K9xEEmZhU7gzpVfqhEWSyf3g/uSiCIok51sL/Nhce/eg6ibXJxUFxKqXDDZYlzeXtX
HOKAJKtuUMgwQDvqD9kizYlUwQgahZ7xnOqA+07Og30uEKWxX8+brjueCIzM8KO1GJ/H+l8oA96k
8o6w7fqWnlgQzn9TXg6gwsroGQHg4/TjxzLN72SXVz4eYLIV8OBmoq0tMlTm3z/PJW+jIMFyU/HM
5KWjUR75lgvwQsFToVQez0mdLjc5+9v+qaf4K21lTY+v/48radR3vpNnRXyIt0AB3TgFXwWf13uT
j2nN8T6wl0/ve3RchFA5uhbj0RBNaFagskEVRDA9lpHJMBDJuCb3nHxBaOUFXnf/3ljp6ZnBcbA6
CtFeZvHmsZg2Q/LaqHrO3GzfczM2fe5U/5GnRcAsTpCNJLVramOT8EdVPoWoLq1WeaGK5eHPnueF
RWrqCr2j/9jDLg8CXAQEDV58Tosk8caieJJHm2GUsRbJ42NmT2qL/H7zDIM4OrcxSs8OOnbqa2/b
wgiAoo30x/eea9QOD7OAo4JId9qXc8BttLPXYu4vWdUA5KfRCSjMvvHTGuFfLtIzfvT7w+43WAot
iQSSkdG9SK0CpeOv4vTaic6XBulppAcF/T4NcFMBDwAUEHXnRwPjpxUEHykL8or53z3aTkUGPc9c
N+dePy4VI9VbN/ScMbCHUsbHldsm11ioj5CgHOA9EhgeLopbDKU/tlJuW4mk1QPEYX8gZPzK+VYn
W5hZ3+yInAO1cmOcyE17sH0GPYfAr/WYO1zvdm9Mo1zjp1D6Zq4YwXo4F6FL8aYnnC5C3LoU8gh7
M74VsgeXc63w1gLNkgCAanwohNX/e+jsQHEgG5iBLNsGoEOI5165Yo3utKrqAok+9qRpfzpGW0w2
imctxHQWqnQeZJFbYbf4LG7F0D2ZLrzoBFpCz1SQeJJCCDCZ1/1S9MiPPjiSlV+DQO0xj1QzeppV
aq3HvHIGv77iViIen475cy2JY6hj2Gztd2iDV+vxwG2SYBhIrCQal4rPDDrSaQUZLfaXx/ZLaqYs
OV7+oHy7w6IzVvorkdrZBiYL124ELtpcpWuWr1Gw3qtfy+5w7wSoUq67kGlzT9vUu71vkrHwEhCx
pKJ7WrIVusf0lAKDnxnt0qGkwwMD5tY+cnFXD9LK7nfrHSYJN+mCajWxc/+y8VM/TYvsaOH8OYGm
IyddFcLgmfohQR4JZwAzkZ2xdd1tcP180j+2Rf2Ma+N1y0iirOT/mJDmsQuEcJTnKo1EswvvW0QW
SjSQWCNWEe9q2sQTDJLwLEY/8VqdeYdgm8gOkyafAAP8s5y+CIL3uUQOdUX0sNAfRpZ+lQrJrdA0
YqONYqAstPToTaFSJavW07CqGBVbDGZDFKT8JoseGOdvHljoYg+MQacP4P/jIthUiAImRjoP4yYM
VICI25Jx5nZ0R1OPFApwCAftwxJyb7kxOtMCnnZV20BYDP611s4mX45jT+QcovvHRRH+98t5nE05
GV8AZd8zApQOoEs4H79NO4JFMe7o8nl0tisoFjLCP36XSuJnWskV95fEjCBvEcShK3OMmbFz+Ybv
LZTU3YUozGR27flzjWsKRLNsnYrfGBVgmHK2vj3t1oUB1uWDJ3ZYlEFYNegt52o4+tTrVtHF2ij/
12+Z9NMs899279RhKFD86ieWjHQVeSFVyJO1Y/06z7wbUe5VUqnWfg+5PUP+7HhQN3slKBpEtHZm
I7RJ+PsLDcNscZPFKsjKdUgcpR5oNuDQc3Mqf91CGELoY/d4CaO27ZLc6Jo+755GOUrJCTxOcajN
tp71m0HEpdKjumCRvs6xnYZuoJNipI98C/A4JVcEhU20QIv2GDIaOZfJdpOSF8BNOp5P/QaRE5M0
uzGm8kgX0Tj3L6QjMrWWF5fztfFZZ7FZtQJmQNosgiGhVduujV3OoJzJGleHhFLTkPjZQGHpkYYK
lhva+BMND6Vw1kyYn5rTvOyCHC30bGwfr5DcbMo5ri42gy4+/pBsr0QjwKfnYfIxRKzJNFusUqXN
hUBqHlYj2burP1AOXQHlc2wyhLY4Mt35N9pZoGrf+Dq/An5VgIJCHLqDyHG3fdyl8HbL+ILhe5E+
C/2LGj0ihKFLpqR9vHznw3q0D5bfvjrLWiamRFQLILRf6rN2E1HyurAAagROgSyNOnJ5qmEEWPpL
e4cTTNpIMRA4pKef8+Oa7EVM2Wy0umqTmb1CjqTfT2QZgvJmn7gca0N75YbZZ3b+iZyQK3OflZn6
nFxER7LUa6PdhrKkqTM2u3XHJeFHO0DgK0bQtnhsaJlvhxDj7PUXhM8/QCE85QLt6Cdwfcf0+T0h
bf5tgqnNZpzDkmU/ts1CcXitjeG0VKS4CzwDeeLgz3uzAUM1Ucq/LKLwrOXITkfyQKYdYsrGDOoi
03FPjExlm37mvzv8rHEqjpiJuy3qiAFkyUTQZtgzHJIf+5jNlnhKMMrGKh4XHDqwNlMrPXybhplE
R9vpRrRJDTSLoPhftaxbvTxClvC1sagoxm4LQushCtUzGN3KwCwKdxjFogWn2DpktcWENX2m93vX
1maU+UsCZNinpresxFCW0svVmRt9/q8+O4wiUQAr2itdMgBqV8BmFfSRTbB8+dgw1LKgyi37YCb9
m1iJEiiLAwODUkrkqbPGGIdABCDgUh7LkEZyzupSFzgZcXnh/C8okCRt0iH9TuJRI+lON35tpSEw
7JMNl6fqcqTKVwxiy4HR/ag2LBk/JVw4zisNF9AcCyUBA+nMYqUtr1n2SH3GUcd5OOjEg9MVxCEj
c5JLo/w/bHOxwbWjKf/cOqb2s9pjHFk2yXZrgID0GKQH8tObYF5b8cYEYyIhGGqlVuhY6DdlNrhI
luj31P/i3hSaIt6rlqTyXUe1TEr987LCxLVX380hh7aP/MQYcxgV4bF8sN6BXT+eqn1AG4jhUD1+
M9MED8/Q2ZJa2YxJeI1NRaahGYwwUdS5rvws9H5ACkExd3V0M1nH71JZTeHR+fPqMWKTOxf1Rq5H
GUQwK8dfy3uE8jfgdOyyIQb8joaQsFmqvp6+zPsbClm6e/v4oVQhZOj8HzEoZSAVZY49RYXtVayi
Y5HNU4/KJwBZqtMG7SBHNaZm6HMZoYjOQe4JPGUTYBi/HYZBSLuw9b7yfejFms1FBRK3AMvslM6Y
mUYmOnr6G71Oe4pXU7/VieAjyoL3iJnJ97LyusW54m753qziq38NgXJdoKMKnXvyvQ83/d8lm9kD
Z6qQ7fjB3keNBWGg2Xtpw57/y2Zyov/HEL61lTYnb87cJnuMUEIxo3rn/GHsBqUKOFQQzftxq5Xq
JmhlQIwNGFwyIgtl0VmqK4q41XLaQGMYNZSPP5fwTDA2DPcW0E3L/a4WqSac2P9VhjLljKYOgkDi
GnP4cXU5mOdNHEnf94jKGlF0VF+JOBR2SFmAgAtizbI8v7cAKhFEPZCbFxXd9e0gXzbRIgYR0mSA
O1nSMxcO16Zi7pTp8zWjjeKnxJ0ZuhfQFJZXf2wOojVCBzEoMUFCO4779t/iGsJZWganxnOWBoHJ
BTfEK2aTuqrv4yC0pKPaQrG9ubjQT4RtKaAn0W0yx7kgNFNRZb10jKYvcBWsL6jkcUSEq7GxpK4Y
JlKTB/EEli0Ul2awYYoOn6Ayz8qQoJO3zusE8Sq4DrTI1CO19cEf3XHYtxU7Lek9Z2hFT0RYCa2y
N6Rxz8Ub47u5qucUJSkkRzHKpXhkcOW6ZARL4RDCOfMOiu0ukyov6UahMMGY9hB59T2LMcQEfwL4
7qOUMxOFqat7YKRr2FZ9kQvLs4W8TAm5WoV4Tq1KvENA6VEu8w69KUyn5LwKnDDNsBfQz2qWzRhW
aUAK3X/iRHcWRWTUKxgxvwi+L60j9PlQsSzCQcGhY505xSKtQ5nKouXb2dNgCouuMTvquaLChNxU
u1g2b+sQZ8BzjRErE9dJ66ADK9Vpb6pngLpjDgOhqr0/QxB0f2km0NieUUetfzjQEqegwIhnRU+z
WIOsVulqgccMtB0b7XbN+RPekD974xnRKrYmTgyp3i+VoZAPom0oz/vl1jQgQfCbm00P8BG10V+L
2eL2DkDirwCAh+bx1i7rRBNQdzpLy57JW/RNCotylyQVJxgUSL/MANZSndYQrMjEsj1BAekiPhZx
FtlISwNC79CsEuE65E4d8Npun/8lyNURbORXNeNKeX8ij/euX/6NbCwrGmC6FPil6SqCxemrEEQW
l66RtUNRWt+DIiSD4myT7HjEn0WcWQ3m3CJGd4CdunYLfeCIZCp3Y0hwtoV72Lz5PK1rZP6BRo/y
UmPwyxNb9qAwMJ0MluJgNBdW1dfZMYYYamRO/uV4K8a8944hzq4lXJ6wVtlK9Pta9jIEV9Dgynoa
txEeL+al6P/4PVQ/mrjntXlh93oQylJwlZ+n7P8vmFNF2uVKbsusk5iCgaACPGvvZJjdtLzpdIDJ
5bCDlpx74HBZbTfzrepIrnhaEOIpxRvSjUAkMTSNflAhThAkU7yytxyr7YGjF7iDRdC8xUUya/BL
qKzKro0cpRIxHUplsEkUTysdl1SwMaivoSLvMHgoPA01qn3mMhNRWlpog7TW3wI9OB/fMfQ87WJc
yWAmIuTHV2VoFHxm515zanLQAUBeau5wWJ84hyShyTcj6cQo3B3u8Bewk8VJrH3pm2drwLCHr4KU
KmgvENW1Ob0fDuSC7Kz8gyTIkz9lgoLmRZmLc2p98Mp+JlY9n+UUDGY9HBQVQOVoT7B6A1HDGsLR
+DuQKMPmAEjyGtunYv7hK5Jwc8FrYIVfIOvu3sXig3yKGIyWhio+BuMj2IhSDpfXVvLaJhZX4yyL
/Zj9bxlKChHJIWACSLRjxU7w1rGhkqOzHTCTvvEhiGTLNbUTrTjff6j8sUZEVfh7f6UZlzO6qKIx
BufOeynMwhOeYnxW9WXwHYGxYOcLRfVj/ucrevoQHbmrpZY7JmZrptss1x15SvY69/enffK4cgzs
tCOYHb1FR4WaiIAs9SrvcoZMsRaES8CJhWvLnIGwtKIKsJeNzH6gfGd+udIDY/gBqmsMOIFBUATh
xGEja+EJBALx/twnTregvnvGjFkIqdm6XOVBleZb8gXIEErvrOoKi4Hf2ssN0IQ1rWmUSyC1u2a/
o45WaymP0Msy3Wc4SRA4tdMQ8X/IbqLj2ZuB4x5N0bVaEMstFSyKLJJqJf9f9IW+HgxlT4oBSoGL
HHsKof3ls/MHhPi1yF4FgCGTPfFZexEbCEx5u/pm9hbzWANSNXg92j9uDZJT8H3aRCPctuvcmCy3
MJN9xp1B1u18zUVkUAYbxQEJYY3BXIHMaxJhJf/xpTqdrWgABZiDBhKy5b4l6vCXkwlIgzsM8UVP
oLGJIxujFPtNM51okBxi/ZZEJ7nrvdgT1s9WzBS9y13bM2rmj4NWaHqdIYZLjAN+Eso+IUrWPywx
HtZ0UgE4FMEbz5jPNACveD1gKo8SkqxJUHGn5HdF5hztypZOfaKHiIg2ELpX8cluhcwTSoEbWPyQ
HXu8e5Ah5aWTld1RdS5p/mYhpSkm5F0dws7/6AOmIuEqiTIIUANHblJz9b/NIg5Qy5PufHdaHZmO
5r/BHS+2Kydq4Fip88UfpV8au7+RG6M7W4DN06/mewrl5kmpE8yBjOIGAcU627Qrt/x6I/NQY2Rr
aVgWqphRoRLWkN4hwdZ4SoCemPwV8A9JNTst1wAgUUK8JXpHxgizloGlnaOFC/BzVImOV7e7VgwS
eT9A9c4RPPYgQWkXq2F089WaCJ1iaUXltArhY58l1FAgQdNSFtdihU2amdz4MSfkBkT5XKyTMa+8
mkkbn8xaK0FpgOZWXQoWjy8URM6lX6VK5H/hAsWFVPherRAhGo46LWbZNzsCJ8dT/PW6m4MZuX91
phEWDGs7WfjeVsFIM7ttLCSvbmg9RdDfHtIFWtiALEkjHtiviRYo71c4CAvRdHnJMlLWLbgeZRGe
RbQUJcJU8hajB9l4BWewQH2YQDMfMAdNsPiAMKdhzlKwOTQ0h64Ctz8WgWWZXYJxerO/ovS12ZFM
/sWBN86IWyY/2TH3cVvNAZ8f/G4LK/nuHLcI3o8kH5dckBv+6Kg8+0AqvlFAm2/e6GvHFEhZP9fo
xuKOcSGx7xZBC0Xkl7QtAZS0ZhpHAf2K7sBxWD20mjwEnxjBlY/12xgZytDOh51qi1yPzm+7yLv/
I8X22R9F/+n20cmxUb3eeZVRC8Jwq7OMFC3RhT4kR3c7ZL9IbWG/mgLohYnVAsiS3K90rGHwl5ey
/bWKlJC9sd4AT7LXN3YXw8nNohh7HoPUdFqgO6zl9tv39GsEypFXtTi66J5+PQ5MVREdiE0x7xnC
rAwKoO66imnTZjC8qPdPOCNmjn8GCYLs9aPmPjnAsNBfPmcRmH8o+fmcl467p7ag4miAsqHXDMee
AN9qx9L908IDAkofeYukE43KTD6YNg6NFkHE32JSp4+HKUJX1v95ipD4O/s359KgKlXx79guE6QJ
oBSJKDp5g/85RPC9Cvk/Int1PlVKpJPhEqP53FLSaAYh9L/EMiiVEe24DkteJyqgZo4wCRvmUII8
hxkSI395eEYTi85MfNtzIjQ/Jl0VWOFjAhJomzJEXmxaZQ0tdUBa0JR00X5IQVjs5KEwybHFWMk9
b2U3aSZYQ72YmUBryYGc+cB6kHl5Ph64v0BaSc0+TMCR5EqR5+VvntHDvNbWeDPNBd/ItdzVHjBM
quq+Cu3wjqq6zoESaShclTHctogkQ7CY7JfSqDce/1rpxC9ee3CLwhTFS9ladNJIv8q3gnttf+qA
P/Fc+7zBjMYVbDE1XERdMtA6MLAABx8DUkey9wgPc6zRWNXm5RVoqbt4ImpCvHrk+ltpLhmXXVa0
JiHiZuaegIdx/McHwR8VqUCAzDQMkNHBPJ6tc/Obfes7SirPg5n5Dzw//vYeS8U/aBw5VsGEk69N
grrEVzJU3jjVvw2ZsalSRylS7IzW3XI3tekklkkyPUzHoMzBpqO0WiqY5v1gGCeEdqeSerhsSoJt
vWqaC/B8m/KCOGMuFbbUYbArYidWOGDEWeFSad/FDf8on8a0k4jXqM+koFSChc4OHbLRrK9iC/Zx
XmXlfWH8DkzvntA31CLi076OS9OF4LZQEPV01ta7Dh4TIvkzuL7BRo5hOwMPNT4k8GQUW96DGcUT
KLUkfhZqG/EOADcCWkk2Mn7lx8aMQTWP2WTij+hpBweS0D5VAXk7d1dXYacUoNQLPjcmcsm4ZvB2
beF32ARNHPNsX/7xzId85WNU+wOPEbGRShMh0FPRpEQAaqBxr7+YrVkpz4m52M38ugtlvRlkkWrb
VV9ffjzy9/ywI4WErM/e9SYHU6LRZ5xohngYF2eyrYMECmM4C/GKm9zfnU5xBG+Wsn2tQpNhr/41
pWvFyHQXiZHjPa5RxBUiDRFhUUxAgki74DN0ffrQ+IP6WnVzO8hTZWBA7zGxNoHQtKd/JCggb2qC
nx8csTgG8oNyF0lIAIlTJxbV1zND/05yBo8B8w3vYZreBXqABGMONx47s+NjDNu786r+FdquRsn8
BU2UAn62Gh19gZZD9CKl6u/bn8oY7B3MG1BsvF8XLZZX0zFCtpnKp5E3BjU6GvQSeDh9DQ4uLcl8
zcpNxhjihyrE4UQRfNEMrSYsjxEU68dgGRRifyMgz0ig8I3yCDa/5gUiUo6hssP3hIuKhRAyfVs3
ji2YKVPfn21JZ1fEla/mA9HtMWLuw4SBXezLZB2DRN1NBdAwexTxR9KH6HdS/Ed3j6sH5I84z9QL
3aDEhAKolb3zzEPucfWRn8+L1zS3sNuQ0I089rjOLXsap9JG/8ldEDlHFQoDphSYxKFOUhsqXCg6
naMCG5OUU4Xxph0zwz3SNtqK3rRq6oqpoZMD5Wh7EWpgZyw6E2QEpbu+ViW7uUOl51xDilUigROs
xauBc4qO08mbs0g0v6vce2DVx2rR11oTqQyqciSa5mZXTHmEt856HIJQ2ga6lSq1UTVADRsH+Ng9
fFaBg9cw6drly1J7d3FP3zQiYAcnsXxv6ILEaNyAK9jUod8uMDI7tupQpl7ixheBzBIrk9tCpus7
rOwPdnoETkym0/1ODnyCx4K+EFNQLWIvXKcbDYdg9WERSJltqvwaLMp4HMp3P0Qae9V9wY7a5Ae6
utQb0UyVuwvYcE1qdazFu69qASZkqqbjrBF4pZA7V8JhinYeRJj9u6qSWmOm8K3oplQtqKUfuG+S
QNwppzNklSg8PpiMO92VBCckzDD7yxgSVXNIrdRwRqAXr/fORnR+zEMgQ7JKB6NhK0O9KrurJCXr
djCoIE/gZaxYDV/1hGLseDvKzDw0iDqZDQWGvxv4/t1a5odrDI4D1Esw3v4V8WAF38jesGbS+vMp
BYlP96sX/EYloSl6W9uhYmYsmt8Ilm8x/dLex0Z0442WwXj1baLjYR9pLGODirwOExUleLJwehYF
IrVLj2rUfjAIVm6VMEV7y63qKNiT614Bfvl5eWAkG0cYf2f6Yk/lOm5eSPu5egS1EH8p+tXQoYZ5
i4M4w2g9UoYSY5DAWpyPqo9RZxzAzV5PXQOscsg8S/I1G64sv/qrKafUiAzO6gWodq1EczH7xj4F
cQGl27ghOwSKHkzrnYG5gbo3G49z4i2c82JmRPxhCcrpM6CsuTgg77K91cVIrVfm570CW3AV4BUl
sf/ydIjAbNp1IJepY5Zc+0sYheeZykgYsaOV5bSkLPz+8WRdyUhppgKa8YhkS7MX/eX+OZv2hTkz
ddd9S5vSmKGrhlmNYXr+uSW8joHxZMaEwRA5d3Ut+vHsz2AtdjRRyEutqyawZhKfX0u0A5vb88dR
sb42EikcejCq2Y4haxlQoLLTDa4gtuve4dGghbCXukspxoWUgxkGUL4L2wnCHVJGnj8DFFKnzMVn
nBHmZhVvCbVktzxOaPXUdrRIqrx4iIJeyp1gtflHyYlMTs2ow2WktV0dJQp1MzbO+Af3I1nRqEM0
q8XWv4y/NXIe2sjnLCDn7shb5yw4JbKZ/O/1s58pHTgkyRhi6aMOWrdcLN9oAOt9+ky/OSIB9fBe
/tWexCBNbvxg7tXxFkKQUtk0u7f1TTKxZdqAktr+aLBqwvjlk1uf+5rSjTkBO+2qj+69JLaSNSkA
2MtR8raFo+1EBBlhmgtP93IuL9F3ml3gcZ8XS90Dsavpk5kSJJn2I1ra+N2apS9vk/PEZ40klCA9
IzSY2hjy6wuumfZIrmNII3UUJcdwROvMwl8ta6TnCdOyr23IO2tBfAWK+sNkAl5TAvKVZRCsuH02
vSRmJ1u+iN+O2hbSd79tSwMB99rGOlZauY+45f1wyO6km0w11iSgMItKGB0aTsuRAixa0JX9BjJ8
/fbtZs+ndca8bYckE1yGMSoRYTrMRQ+SdLex5De87YjE2GcD5w1lA6JJNzzThuHjB9yS6zXrm82t
3RDqE+LcFmUr/beycx9Wa+OfWaYAEQxlRbOO3F/+/TcJiV/+m4kibYis+2HsU1LaM7xoN1nsFy0j
nPHNKHJt+ljrFYgTNZNQoMmp/innUnwm3LW90miZtcoEJBo/tCAlRYD5/f1jX2EbiIlviGj5/94G
uavm8pToVZWFrtjCWsr2IGinMq37xVMtfUVDhrEwylHRPUSLKcwhpWA2cY4SgTw384YQ8v997/86
Pr16ydn3akELIRejSXJmxqVBZCmNp+aZTm3dOkpQRPc6HE6ufuAJprjeAEQIJMo8ltv7XXWwq7rd
ARVEy5FxvCb7V+JcdqWdwLlxSySm0sWzSQXdxU9eI7rw0m/jo9RV/2JclZrSXGN1btqxfmI5tNrz
QtQmYPstes42x0MaMXRAm94okQmziRRY4XJ29saRYiKRm+kDd1ZA9t1V5exKl0CCiWLh4b6n1/u6
vDmk+G1Cvi6toHyPKeSlbJHXFhaFSmjHb6iuEILcKnV2lRO0fb37/EhmI4DIKBR20CJFOSa9x4yd
QpkGi6q/rJ+T6BOry/unx/Jqk/bKZNBAlzclMubaxnQQzmprqu0gBJ1ekyB9P9ZqCn1Tmhu8HtTa
Rl83wCFG5iNWCNgRIuOc+fwOBQSy8cX/3Q/OW4rGvueI6fgs3b7KdCR/Atn4Pd4d6tr18wg9gZDV
dz/9qZ/5IanNh+v/ioe7/t2scZGxwrwgecAhLHBqOPawI3oVc/TmpB07aq2mVEb7bM67ksLefgKK
BGyrarRzmk8mPenK6b+2W3GLZV+ttH1HckMn4kXsXiNr4Lip9qxmUzviGum/kaloBag4zXDPmRWi
evUEk3kT1vC1o3kkBLu0qDtCG3c4j8V5xR+Z2IvZ7SRXLTJlz2RRpunMaw752f3kPTfddQ6ZKn6p
CbyKbdnVirGdGKNOeSlvDe+7x7IeZEqKjzPW4FOOd0oXqb4VJk0+vkE0HmEubN9PDIMs5vzGey1/
rAYyWJiYoRSfV9cpfOj5iBzry+M4OQe0lW0ybbjl06JwcI3/BuAtpGdagYzno1jPBcKLfQc+zW0g
9E2ZV+OSsYTyYcG4IpFsGpZs0eAAY/PTb+ydl4XhGwZv3rx0auvq/sp4PFq7QdME2XmeRYpz9mo2
HJrh6x61CfJLpZbw0XIw9oimVAQsIAca5CEje0f/AFbk8/8Szc9gpCs17yiZ8Fp8Gn1Dz1xiJPzZ
PEp/jmY7gH04KqrOtLoIrs7oYkAsN8I85mTA+ByQGVGPIRWJEHmAdgjEM1/hSgiTWXp/tgAyUBkW
FGfUp0HQ82rP8+1FHLvjsRdhm9trlzfHZUIK/Q3SJW84CJGjbIZOTdAfnp1oy4AR+mWzuU57a0aB
HekNgC86FdLMXIGn65NU90VUHUPvKObKaKOxpXPqti0DEpNZ9GkW0G/UEvmIhf/cO0ayseDsV/Eb
CHoTokl39kOsKN7eIT1F3Z+E7OYr19UQgQ9uf+MgHjY5U0J3q1swB1QaMvFE2vRuiz/Pf2Xx9qTj
x5eEa0D0CrdDavOhhWfktHkridVtgghl4byag+0potE5vVbpsw+uFBMP9SnnQIFw+CHDfbkNRAzC
pIEGqFHD7MlPR6WsNpM2ZDJssRUdpv/RFOyoQwxoPeWEffelbipv1ruUFcdz1Qnd27pST8pd29/L
1aYisvYDIk0LSETlSJcJvEdDGFQiZJcVnxitH2Zq5pYGfw37iJvB9/JzURg8S0J1u5IIIlkxZSfK
7486kkBtjI2geGxIP2O21cSSuyf22H8bdxY8pxQ3bYiMu7soMayHj3NvDl9ZxlsxBHkEuCQZ8w0i
udBsrwoCvf9oxUcOxV0kbM1pDtThDiWEpr2R+ejVgUVYIinTMQSLxObTYNcQnp3yrPLuMCX45VLe
CkBif3RvmLHSAmKuGhJIa5+V4Un6E9bxWGfOSNlqcawLv7hfu9kWLgwZwb7G/toK6/6C6bQnZPzg
HHIjAyt8VqAci3RRkCN2KEy9RdXb+2Wp3/BJTSfT7SAuSsOagZxRl1tQsbQuIHDQkJHbeyRb3iUv
RsvJSbR+46LKVyVDlgJS1b9RFNCtx5zGruhMWqt/es0BwU5YAaGcH4Us8veel/nMzXH9XjnN6dTA
ZCXxq/XlrdwZzKY5iSz8D5621PkR2lGTZQ+fn4GOeWmiy5hzfCsVBECD906OeS83/flFBfO2QJtV
vq4UTHPkaieC3sKNu6KgJKvd0+cRcFH7sfHhsB2nNBK750l+7mF8dlFV7jpecQway7Y3ePjJcmVu
oLlntz4sQjhcfFAES1X/DNS8v/zI5qIn/6DssPUHqMeU47tc3Mb1Yg6jCoNAKAI0t491zln1l/LP
N4f7Xv9MEUMqJ6xxWS5+KVaIHOUrKX1Pm2Wc03Fj4XEwcPx1amCK3Y35Z/+hhHaxLyyL4BLCTLgM
nyWJv86JMyNnaZJwhXkZBAsSCkoPAf4GtwmNRz/RjKqRaxceNDEw2/X2AJZwa0EsJBMwvZ6U5IgQ
duEsZDmK4Q95vUmGwe5rRiK3wNaQ7STkEgOw4fsHVYrQstKXxsOs7wJEo6UBWvCpnjtEOcnRLI9c
qSuUqzj4Qto+Qb4mxbKjZsYX3phrDILUD4+dQPih5noaBuUNiZcrygUaIUN2OwN5ZjvPZrbKEXUj
ln73zFIZf9uStt4PxJmgTIp7HFEbOjPva9Svfxt77PyWvOYqcsBO0Y0i22IiIs/jXeTp2OyC4mqG
86WA/ZH1LuzSgVthwnVGlJT5ONPrachyppGRRE+WbOtdLBCX/ffqHaNhnKm4eKDhfru9ExRHWEiW
9a3YCZLInn251cxTYEz6GaZyaFf6CjIcknfTaRbw8ftG/LESKjPowBelWAWynUkAZHUTSYc5RcyB
hu2qzxsS512Vuem0NY4IqcUP1CvOmHNd4Y5BgP5VjSaxwSjNPInFykhqlgOWi+06r1tQClerzx10
riRBFVDDmxl7YCfrkEIeJ5xERLh3b8REhiTAzB2ac0YQwRxe0NztUsep4fyWo/T+i9xnQSJoTVAo
mZFWQlKu/U/df9j8XRekDa/hTsj8MYLYmjm6OzD3aFiXmTjyhCg4i4nWxM3RuQdJoEvcANlghKPD
95rW8QaxXqK29w0vegWEYYwQiQNzwZswKjC7zBs/0fdfl7ddG4fZnX+q6ZyUgixaiR+nFF9V+rnx
9rGQQt90iKzpdAy25j6nJ1qDdOjIs7bh91gGjpplUslS6E07sLIfGtzxk3kwWdX2Ld2y61YAavzh
U9e72an8G89NhUnu0enx0zVSrh6lF0zIpFwbRikL6FDNhhVRXbK4/fx4uyqq4Uu+GF5NuPd6dZB0
gL3vQdDUEYPbE6Ijho6/OQQkCIiuTjS6sbu+gPvMh69wlm+dYzfWdFknppxRIYFm6x6b7KVktMKl
CPy3lBhFi4sjH5tSwwfQxBapQmjNz16ypGHQdgo/wnEYXBS8Ap2pzl1UIk+Ma3bNO85wMve1wkdw
RCGjAc/hcnRpVyf35H9s5FO0YSnJ14P4EunyvBiDSfye+dlmKWVFEZfy8a7RERC09dPjtMhhfeQI
fVTmrzHtEATR5LX4fKnd7MnKRHZz8iHbNfu1lOpiQHWPuB2poi1tRVg48F3AzMqt4W3IjwY1C4Ph
Qi9b5yfzbvjxyQCcS4DL33H/6XXhzbO7VGiE/mmFR+4W5YWb5CnvTtHg7dv2OQDkUxXXbuIN5y0R
E3u0VZY8Z/h4yw270WzrA8Dx6wahY2HA8PUsTFD/BlW3Fiq2kB9YJUYWscQRPFzvBCDyUUyZrk5b
ws1KHdXS1AzI9MsFJbW/yrwXoJAnc4Bb2fGtyC/m5HIYbfNfJCaot36GSx1zL8VnwNZt6buP2CjO
ApWAjbo9kT31g/KiVBF0Pt+b2ibXTXPf1DXDs5ELaypiYMGNXL9A14yPmp8GKtDeU4VZzAc9178t
LwjotbERU7MvyE6y9gqnudfj1DzoOJ0ZuhiaOtwARMEIu1s3z+9ladcWlH7efSYcWx4pHU4oqSeU
1h6hfXLKNd6Vg2tSfmJz9DE14jhSeD7ZLZCcr27XpL0CZ0qG8YFJljAd3BL5CaaXlqhKWmB2V++x
P9iDlKcOc92hzXt9EvqcwbUa1tJr5tZO87i6AiBiH5ydB3w0Uj4Tc0IZEdzUvUiLEywVJYbFcvV6
d/ebXf6n722wkfwd6quf+z596kJ2LH5sqeBwyUY3jq3fNPxyiVsjguUSfXwwY4yTiei1iZ2/xy8j
DjBLj08C8iIvb4ho81eCSaNl4Sbq/T69lHGstvc04swyJwSJAh3dy5x/ofGzPIQL+KcE3cnrsk4+
poQPR0e5nPlKkXl71Bw42r5MrJHPJB2l9FatTguBRmS2P+keNTOhfqzCFPViOq/fSbneWlWbKUzP
2ZXZk6ONqB8pOm89M2AA6KARxjYA4zweeFnEZSKDQRlYBL84hn1ActMs0ggzhAauHQ6+Rkf0pjDq
vUXFJendJ7lRtFa3kIYEcTByuqWafA7TyuPoPmuQve48V+1RKTYR1nK2IHVgqBO9znj6FXbfkRMr
64bqgJT1LxH9Bd6ULlrAkl8FKl45WXYggJmfECX1dk4IpPFg9zUGN3RXT8FkO8nZiIC1r5CLbDy2
kZNcgxCKuFiVaeBz44yPM+EIyUenEY2lHIbuLbKZ1lyHfZlqNpAatuETju4XT3BcFtaMKTdWeA4B
McNtV15vGpM+Ftq4bzbWokW46ZzV5EtO7J0uYHkcPSYl57WhjdwNQt227Oq0ZwC8OOl8TKBC68As
l4IfHwHX/tQjez5uLVzhIVy9IIhwUgXqe6JEGQj/KdJSdObS0EweAK03M0iYahoe7vA/umTaclF+
7RAZtpaApJIN4kfpixNDHTh0lpXDLwPOX8XoaOVYKZDHeXR/2VT7mPFYSeodcMmNBxRdJu2JIoJx
RilaVFV9fjR/lHu1xZEHZamRfw30IdY3IJMSFXBb5/RydAFOxUEAjsmQbuDRBXZ9smBv0UTqJ5Bu
wjQnOuTQxJ0qCU3wTWAMCSj9wGwzxQsGLTzFUfPWtx3Ibw5Acrdb2es6Syw4vV37qguyYZ2lhdQS
Q1NjM8K191NwpfiPlz7VioohkMN5ccgd92W42AYIjewGQ6pNUF/WZPJwE1oe/Ot1OzVokFhRiwui
keRpkiSoXUBn1niiR2JypCRtBVKK6PlRN9W5eicX++KdnZZHbdB5QzLOxQC/ioqtplEUhYf6KTut
iHfQb/XJLiwNPSdMpNi/WnZpC8D+JSWeNBypuHf/+etOB/YKbFUrb6prVlHDGww0U+sDhkMLkDte
XS7FtFU9pxVug6t5cTQNgtdrYtW+QT/FksPz3nHButuUESRnh1YbKCHYdjPxeqWPFmePTziJSMro
Ai5MWRtGD96Klzl9cg3SfK6t1z2EMFEfp1bBviOEASk/aGvL7Imr7KEpJQVkxELvYiFg12AKS6wc
ykALIBxzpvXEdseTNevP8TPvFitkzlmuo2nlQcJk/FFk4tCPLVmxb5+w4jTqUmbM2tNbv2GaegKx
kKdARkQqrwEEbVkZITTNxpgPGIS/tIVTeNHiGCnNeQG9yxY0+7Q3C6QId8FrZPIGiPwSRQCgFsf5
Lk4CkxLiAZ/39pRFezW4MBwqgde+UXKS9oRQ6E+0sFAgCley9gg9KF+6+/NYYv7TrqTZKAQ+az07
7NlRChx698KU60Zsa4TIBl1jQ3qhhZ5drwEuXEhoTRcTa4UF5woIk2ysTPBSUEqGxManG7j9H36x
fGEacLvUizkJywqgQ3i8w5mJFanrqZZL3QSSH6V0gX4FlGtiNOksyMRkrHAk+9B0lfqAgWXggtxZ
22zKJ1NJMnPk21oAv1kH8Rj23pOlcSbX6bCiYut/GC/NxQseX/szth2bRSG5NdOu3r1oLx3mPITG
O2XSLM1tZEut661EQ2g4rV/63JVdioF52pbRXrgEHD+RXwkUFZBU04QtDxyleECl7Pdmwl9NNEaU
Bu5VQA58qBSh6iVDn6r4k4YqDPkTL6FuApWUzaBuo2mcUb9BkxcWgg1jwPR2j5VypG/kBtrNshcc
2ek8h/U9koY2xaFKtO4G2IhHlGqTN66vQVf1qPnzPVxynVe1CMayj8IQq8aqNNpDWU/RWEtf016G
ZWowKec7afOeH0N3DxQyYvxA2mYixyhtn4bkKtmGqZIckzsllPNxGSlC7DQ9pI3Rus5r/4Ha+ZIg
HrCV9N+UDaLVe3L/af7xB8lTx/EFETHmxqOeygyPW4js2TALca/pe53i3t+Ie5WAikEQ2REgboUb
YaVCfP/IrOe39d27MjvnfX+2S+wXJyYqSR5oT7McIu/US+2MQnd9noC80tqs7dRV96ob0X2ARgUs
UFH7KRjgDFi2UDVvIIfSS3jFU5UpA6xt58SxnegWCHoQg7A9xhnT25Y+en9yzbHEu8sl22p9ABHw
Houtv/kLMHWksMz91wP59lOlPhrNaYbUb9BMg2urC4J6R3xje1PQjlNv+CZpkEo7Ueww75h0mYvi
xjq0ie6tVITj1YQXPyf21VFHMa/F4qffa5GnssWrSJ3JEZH4FgdqYBn3eY3oCAfMXu/+hKpeBNgv
vCqGegmJ3+HKS37BoCMlmEeBwF38Pfyg4I+FAVN1Am0+IvxPULIYsmXr/qd4tUHU7XRz3EI+rGQE
hmuspCylIT+VYbv7XFyz0LhXG9uJEUvgJRnh1awMZgDtidf8ON5j/Nxrf+nG/xEBjETR3wZx/U+r
X+W0nm0IHHF+fYDFSHKEjgGWr4ADeFS79fRrKC1tROz8eU0f7PtJNJ64Mbtrnq1Yq3F0J6PxUNbX
A7z6tVfDnkx/g09zvq6cCvJZc+6miKNzVey0YTqA5NlMB4qXG6Z4aPQFEHSha33VpuKyQZ34dsYg
yIjJESgOawZUULZCait+UHO3CUdUUYWzEdLjNi4MuJN1Aa7Qb7jbF+eQx/9F18wdLY+MH6E1D4Yw
Jl2Py/KHKrZWb21BjXfWS61h4KBd4FIBoo4lEl3/tPFGlYz9h9CsaZ7wmfrrqDYDLJWD/Y0249YC
frqqTuKrWN7LSPUvtLFWkWkO9Tj4e8y/p4WHQUv2393sDVYIayiOZJrIUD9m6diZjzvRS9Bdikwn
4mCGNO5aHIpp6gp68CPCLHXXZkda4+qO6VxbjUTtZ6A+SqNfKMuhTLgga6xbTCXDkYwOw1c/yg5O
+BKpMp7EnlNxRz397u7Bs9+bwGwUzLB84qno3d9lk2aiE/zxstNLI5TVz1gq0J1cb0AjbM+7CPkC
qRLYJ1LLJe0C0mPb7j7tdHYmACpoQY+eLqUG8/vzOsZYm20xGRrGyoMVVs6NXczHDmA9U3pCPL12
+jvjIZALiB3ToIrckCihMsCmOoYRk3PFUNrlzkm3v/p0x+XuM4ZlAaTNasVOSIzT/MqiyAszMEiN
1xWqZvKUoxvX3ALtyOLwoH4SgOO79Qlw7ASfo8zO0voDNdozCz5WDgFsDwxIyQuIGD00hyJnrfYQ
P0cLRUXE2powvox6PLoafcfA0ex5UivRWOaMbDOjvk8lSVRodXP/REGGWuShpHuK3ZCiUVbCZkrE
tMgnPGe8Gz9VIpyYM/ym08OARs3bwgIqjBCKO9Ya/W9cnZ2rJy9E7LX52ChE4HD/2YWhKfx0IFeL
DKAuHbpEpSKDEtaHIcR6nloE1BrKkacodPeOie3NSyI3+MQsFRSbeRCBVs26g39+Iig2/0ejSkEY
rv1Xka6+bhRpvXHNDOGh/fP5wxFOQSCeS6P9HAI0DIhP8MB1YfATKACG6bv8FYMgfUmQtt77HXEy
NesGKJNnPDWmNmByEmi3ha+/3duTGr8BiVxyzGKH57BxtxcBkLodCLNDz5AAqlB/p+xVr+qapXPx
gafWEsqqpJSP4XV4H/h4Lg4E8U07LsPKQrB1X/3Vy18Zz9JvHmtu0UveDfjkt27q0/2djj1sTjVY
WdLSV72McpabJ3PhTDupkohrkyRbIa0BqKVBmh1eWB5zNPg7peFs1RjSFRyCQdE3pN3z1YT6uiS5
AAcdnxJtkMJPljTg+j4eiaosVAHrRAEzn0Dp52tldKaa/ZFnjDCwP7aAT+LROhR/L7Hl5ZANJCB0
NC5IRXm6XaVLhzcwafCs0Dm7D0jdcNzorVGxNFk3ra2B0Dkw+Chs6mftHeIQvMlCLHgSf3S0JZ31
S9mWWeF68aL72tL0vA7QM+xLZCXb5g8ra0tnTJnaCh3lk5xS42xjXKOdAwym/rMfp75oyCvYSzN3
KunzY0WL76oG5cOcXGqzzwQQoWMIsCcxbOuhYbPQjIB4OWdew5VfLOazk60MlRTQP8PzQpQLCWmw
EEchu2dvBcfmAJoe1UCRo3RTF4WV1VULNA30oJdc+hvCuwzA6WCTgV96H0atNPAeuP9Ui6/aY2UQ
AUicB+esEOPm2yArZkT8cC/u/Q4OGea7z6jaWTxD30CHNDLNdbb/bj3PWQaqbcM8cvBbHEGg9kyo
U+Ya0QIw7VbDVQtxqlCQ61PfYCnzbM25cuKQTeegx8/NuLhf/tzcq6jHV4yZ5GrpYBiN41KZf/FW
T0i8JBQIFPBEgG3he2gm8Pnln7OtDQDCMjvVgJvgA3vDay4adH2FPxRVAHGQYNXLmgGoOvg5WCoS
rPs3oT65CVlOZJQQpP5rDlpGaK+Vhol5MNUVBbEG/8ZgHXYf3RLLtw19UmOcCbW7f6XZTXFj8QIw
6woV85Oxfb0XcdRUlPUORRegayr3wMkghW+u4FtmBRiGtaUJsYkXH3f08VhoWukdljqJLlcZLKnv
Gchdk+dLAMZ266NTcQp0tafA8drWMIT3n7YijRnaQYR8o+zIbW34h7/zGQiW5vw9K9BeM6htV/SN
wMvS38/UhWcwdgKBVkXJwTzHmKOsifw3sODmsqAYrlweiPgn9PLs0S7ZY9U8ZOMkty9dcCdbCKLh
WoXqmnwOByA8LUvjYK0BrAlQG5UPBRisIu/R4c+E4rbzP6EmAeXZMJcQpVRD8L+VLYYbRkTP6jx7
18ebwiE8kLFtztWVWBk7KZU1R5dtPyPh75FAmgcNlrbeY7zCOmZhkKRX66XS9/lqHwX8WCHQShPR
9oxrfy9kofG45vyK4s1hOJFQFu5LCFivZ2rkAMr+im6MBrli5cWvE2Bc5Ukpp/SreLIM0TaH0PAn
scZLrqTTiTduQzDtceu6Z1jjCtdHzawum42aMNeCRRNTnQUFON2SqcQ0g1wp9fAkYs86yKFuO0UV
/H3dIAK8Xv5JdWZNn+7IYO9G+yrvG/ytZxJjxrej8V50NWEH968JzQUbuM4H2EjwooslRpyS8eIr
qRKco+orhX7x2jxK/l30odERxF+/H71c+SXObTnKo9TNaVcNkfVsNaL5GbQAEi9kSrbEkbTdLGme
cbwtgmPCUwz8axW9aIwh4ZExcvPFFS1nUqv5Ve+dz+UlLCaCepJtiE7f3WweKIDbu6Q2Uggkt4WX
wRw4Z5PT7go7HoNuP48NFlO5ApjpRM4BzWnfScJDZZV9UbKltj8NqAwAb0Owu6wbxYeDoZ8wufoE
APgb6a7WrfIy64vRj3ttUgIkJO8jxYZXjp73e/U4ZAXcdDCQEaeBjtiuTXZrUeZMjTQc2WjTamLf
mdDmGB1H3eiksfLVAoK5TUeRZYDGk68yYuVouTL+ZokN9aulwWU2gmPVQS/WaL0ztSt3OLWP9c4F
5UGjkfRk9qAt9x3f1sICZuwHRIEsWqTqD4zzhCufOIPWLbD2gQx5xdST9dYDUwJO4bH+/W2o6PkI
vsEUEBrKo/RWxo6L4Fx0nJWlXKafTZPu6wMoXweU8i3JsXwXSLBse/oFauDBESwCeQyU0cGDfxjO
2U2rcmOpz58TIzb9JuYDxka2ca8i5vFblZ7ALP59wcl5CqCe0Q0USuvsP3r4L/YU0uYXISLhF7CO
9OdeZKyJVysUd9kXxpXgAYEqcif8DZsd60ZBG9ccDlF6u/T6F+iBrdW6He11bKWGHyAncCYjgk4z
xIro/Lpon5vPZWPtDZ7lOdSrhvGmXYENfxbZsJqdwSB6a5Y9jQSW2W1nxsQnXz1y9fic5w5lHM7S
SmM4i5qe40EDz96C/xwiJMcUs+O0oqOg5g2Kx4DuKkb9lI0pITmhByY5DfkQW0BoEHGLBCPmw1bk
Qrc4s0A4Ft+Grw8i0HrzVJQVfO0ZaETPw/hkU+kAijP8mDiEm2j2HQY2ddAuBbdFlDMkb8FVQYCE
DwUwR4qBJBMuYmeS6QalMFgLfHPrd7teAZTrudGyfG5tSGeatyq+Uw/MEpd2iuyVg/UNp0kspu4i
RooAOUa6SiX+R4jH3Mn2CjftFWX0/vMKrF4DoOT92lDRPDzHYqaMRdzPoXs7zCP68TcpIeZD81Je
k+kUX/KcZcZrz/+WjdSIGeTcCEbLwnGgiYwU7c4FMGbSzVA8Kv6ZSDSSV70SUsAJNZKQY838bPfQ
p6xqeBr4C8Bl6j9+eqQMn84/c00bezYNQXKA9M23aCvadx0olihxt76myTBjPy9JsOn8gE+cTYj8
up0MKkPnStoSpKhHvEtoPZ53hLQ3Ntd1Fbty+kHPQ87J7qpT85hZBHRZKhUb33JDT7D/hG0QLJ4g
Gxk2H48OiHPvm+cfqsIppNwyrSWSnALuK2vf4egBOdOR0AdSO8f2AManxf9shYdhp8zeDLqkJaG+
8F5Qz+R6pMpA5en+yWlEO+ojHKoq+8hd3qfuu0VEWuZbJh+WZuqgZYlauSnK0dHa7KfXRz7u/3SK
evzrqQhgIy6FLRb4cWiQNbKqnUd0wSuJMn09s6GlWCqbMxvtDiPJcCwNFWBNxy9o8FG0Z54EBM3i
tomR19I3PFz0aB4i400Qy0QOc8b/X0A5j1U5LYAx5gv5fRlA6O58M0TBKp6wKEdUBKSc1yGS05B1
DH+JbXTXdyUqZSTy6+1Vgk8JDQ51BIJIn/wv4BeoXuqqjACdf+R/MMI9pUGNteWdiYBAo7e+aXgm
/13uS/eisOPkgsrIv5k5aquGoimNa28ufvZNBjCfj9KP+o7rPfLZ4cLS7h5Z5k+cvLBuWoNzOKo/
OMAOc7m/+EadU7/VXfztE/yCXj8lBI+sK2/MZrLgWgSfGmcTztgWb1bKAd93oj6aNld8WUwPrTKz
wSIeSPWJ9nCnkCyXFYCHO3ft/giqkgEUITbKqIWBr43c56ojQgxjJUswoLT0oKZ9xRPS7mU/1v1t
rtiNuMbsr220TX19X3g2KPBcz/Smxt1KjO8teewcOcXS4dnEOueiDmzwvUvxeWxYUp9hBPI+wODy
ceMUauNJhWxS2UjITTipYN6AZAW1yjqabTGVohOy5csLcmoTRJ5oMaUlnJvayNbjbA7qmzCM3Mzp
G0Uqf2sMYQrtjWoZI6HE5vrjNjn0yGMbnkACGJrnLzEg2ul0K2egcproPFbBA2YceM8i2S95mPFP
9e25fZ2AxOER97hLWH+4vygoIdFfMWPfqywsNIqtG4MSmLeoT4+jLp/RF3f4b8ck+WTSpbUfBFQz
4FGWVMFxQVUEXaSEbOh+TvcYFe3DmLET/tR8sefiFuKx/9wdpdBPrHtP+RcDURQuP6Bjo5UAKdso
tRCaS67ePNejSNPlpk9R1L07dus9MYbwD01pxNjGsbNfcoaNBD9+NtmBda1kaTvzI4UiK6Sm9eeW
4iRVNbX99JPKhkirOYVP3gJR8nQ/Cpe3vB1GuzzdJXaGkU5fitMk3yd7/V/RPT3lS82unEnA4DU8
y44TGnjZRevpc9LY/qL8K5FSJoekSSJbCQAlF3oS1siVsaB30G2XshJhASoK+Tr2oghyWKZWQyrt
/6ryuar+DdV5PAG7yr+cuSgcGajnzpBiIzeL+2ezhcaDhEoGVRKQKQeLDfH/gNthnk7/GXdGLM28
1pNnzOt76LdjlGTs/BCZKTY7/3bRz77YnLZhaBmhmb8zWhZ6p5sVlPGAEHo35QGNuftBxSf9IXxr
VpX+BYErf7i939phCiJeYSdFIRIFw+24Ro8Wt4r8cnyRexiM78uWlbD7VRxWbCheYzrmDFr3bpzA
7dajYNyu5BM7OxhQmLPI9wF1ECjebeJLi1Gkdv0LN4mOW7HMgH4iToylo70EU2H7IlK6jnadyx9q
EspApF1Bl/QTqc7YcXq/4FKAjOroeidi365D/co/abnJaBAJYuyXVf91gAkz/n09W00t8ALtFOpS
Qow1BysR1aoSnUUvQCr/jV1QAQaoPyXs+cm/6BVaMtcnGP7ovcnRd52MdkM8op/CoDhZRf1hHxC3
lAA+CcijNuuXdiHUAzhgCP1FQlp/BkG7L4qmseJI5WXzCnGtrLB7zP0VT1mJN8Frr/fYkNCK0pMg
khWLd5Td5dXI7sX3Id6sD48LCMBqg/G6am2O+5zIKUMsj+9i0GSmFQlSeqz1hDt1wbRAHXidRl7m
GvCnguPvK8WEi6zxPPX8mjiT27/Ri2tIIxhOsyfmnTWPTXGwXyC2+2u2oloEldEIVpze11NZq+91
R54QMUyGIQxAJBnQQqmWY96VFSqouRoREFKGpeRWHnDq+GHtT9AuGOPyejb/29mUrpKbXttTBYTH
Vj6loEiQ94u+xmjsE3QaU9DYxTkO+qTosnoAsaT9ZP9nEprF9cXWPJdDY9qwMIZvdpykfrfiDo9u
usul/Y9v9AA7mn+7Z+PXyezHV2qTszA0Oja7X+gJMxx1WMFmmNGiUwNu8gPVqVLc8aeG+ELt9nqK
cyDC4tQe4WS+gxH/5lXOXDz76t2Ti7h+CDJ1x89N9J7SBS5LoE5Yv57bkG9wMqQyy+I7hKjOk51C
MFFG4yRzOuqCvQa7DZ9XBYNVCtMH2mESTSCVHFdI3kdJOJPofzgoW7UyIajE1wqp7VeHyWwGvj9E
WWIUYTkC0+fnQSjU12cckTY4sDVr5CdUfQdSOu8hVHsxeNbYOw5EUAu3kCPg7nGTKtpRGMDoyAeK
3hJ+fvjPizlWNz1U5oE2u50pp99up9VtgsqUT3Xz4kALy5fq6SeUethYNEdFcM7Z2VLoZkU2zff/
iqCa9EysvBChIWNiolY6J4JZhd5WzFic8XTrPVcUNA26sQXCkuoj1gavbP3RD9DVIQWA/s5YKNCY
oSyzAj+nae0Zj4nfqKrgq7MJYrcgqbdJwyBsr97GtMmSBa9ONE7/ZXIHgHPgBAPZOyZ4wJRdFUZy
j5XNO60VOzAjvj8AM2w6IzPr4uKkNjusi7tmYEq8OEZWjK8g11YzSPY95w3U1xhl+Q7/HKs2EhBL
a/VA+r1E5xb2nRpvGys5p8HFE3eaWCvTw3ujWUpmBdW1rzhkTmtCPCtvNiNscJJzI18sZqhBTt7V
3M/agOF2sLT1b7F5+0li5eGWCiX0Viw1G6jgE2254CGDRXXRljHiUaEz8+QZYs2PnCWG8UvWwvK5
hohZcwLvSDuR/wiLEayjDBl6WCUEUkobbjlXJt1EwNw8xTzPE121EyNHWUYmxuVFjs5scNY8YkDZ
jFUIg1SRUMbEB7P3sc8dBULfsI8nW8dxDOUO41/87JEb/l04OVjjU5B0Szcq1f9nWEqpIcRDfztM
JN+oVwfZpU9lfYWx9TUKr/bLyU35J6H2KRVIJtZsHYNyAFeLFyw1GHaqTLW/x07M/Llo++uYsUWr
hwFKj9ELVZ7Oz5kqC/ccHobTup1+K2nR0fbKbGYqPYLhylVdHiu+5r9DgWzh17n1sNmcd3ssYEdG
IRRy6PPihCPJkEtHP3FuhYMkyhjXo2eVWV7Vss4zxD7tBIwICdMyr4iJk4iozNOuP24Iih6fEYLu
G1u9VNvpJKgiXaR1FOPVcgUErG/0vKgO+inxuG3noScMfNhshvOU1z7ef6Qf92aeC5dIJKtxog0x
K4DwEO6sNN5uV+MUies5p/nhAir/fcTwKE7zS7+YIQi9/Cu2m+s7D8+zuI1xYSZ58FJQHodmHgcq
rvX+4qHcOQbzTviCiBlPiDSWaiaFGXEnDrA6k+t8hHJBQaxV5Sh9cllP9t0mUf6nMP0vxO/9+PqP
tp5ui8tr8pbW1zIdo3Akqa5StqYo37MT0Kjb7zzRaD6dfcvFTTyHPcJ9aapqonDEyw20SDOjlbse
pf9zTMmR2TMTVM631sEX2RNkddUEEgKMkwRXnQWHuwm/lXgj1OwwXue7d4zsJjkwCKQK1Unwvt/D
8V7C6RIiIJiOIu5pvovbEyQLzueZbic2B6UyDvUYJY98Hd3jSTYMmEj9gDV6MAkT6ap3KMA4Dzvf
DzEI+aQ2PSVwsm2SyjxSNslYjekq9QwUA55NXFXWc09q1Y1rW5Pt7D58qPK/PdROBYco3znzAIO7
MAXSPfaFKanUVz/VSmztUj6F1AaaQsYOz6QWi2Vu6emGpg8182oaJqZn6VOE8aufQA79QmU9pLEk
avkiYVnf41eR7VOZO3y6Jtlyv/gF7HVVheefsJXTKdF2lMkRMwIysO94lSRzryVMfBsaxdLQJlbv
KQ4zSECluAKCGfpokszchT8562N/HOBWZrtaY1eovMVeHtzVJNrgf9ViDRrlseap1gaN8+6dKdnb
kL6p80IOh6GdYmW5deQ3fR438S9pCfBz5l5oVqI1ZcS3HhYx/HoUNLjVRt3LQjyAl4h8jirt1ozV
hpxhsLPmHfN1Hn+NkmhlBb5iIS51usCIqgN5+dVCubLi6pT98P9hpnLYhX12TLhEETdumi14Mz99
ex5RNdFWgpx7ZF2lCkMjRlJDEKqutmJwucaadPk5yEVHV609Qlzs6NsGwVScKlUmjb4hpZZNEwKW
DNjrRAFoZWQ/6bVJNNzosrAuaXzJHoNTCsj/NkXfEgH9abLx316a+k08VfdVDYD+0IUjVR33CBaV
FD1vnU7/MxN4JOWqKAsfy6/utNcWoHl4XLhyR+2r6+QPl/QW8Wl3plo2DVwiE8F9/nUVMBAG6rQ4
7q1LxtfTt9b5gZ00EnTA6mGXQ6k2QnNbucxla/HOkXtDRc2wgjW56DPmn13/ARSCo7CbmAImYkG1
PbqqTrLFSS5/x/qzEIEbTI0JE/MswUZxFe7WmPaeRY1pmH3vjGAWGXcKb4pGNLEHe/YPRApvdaAG
6hviLGePuAYg4NQKaJulwNPaSmMGjpFNmJn8Zs3l157ndC7GbY+irosWIWcUe0iPqrw+KYT2PA+k
zAjWiio8/wbx6u2gN23GvUxipbooyyyBt9ukG34maN2XNCGmu77vF+O8+GiGQs2TjiA6ObgGaBCC
JQQ17/ZazuZDFt2YKkyhVd8y4mqsCE4ZxcZ0lEVKQsysjCyWdMkY3axCcgC80YXNgew5wbLqkjJe
ikIw5vu3HLvHA6zfV9zP+EB5usyITOVyC0NE2RK0jgPzIXfDPasquecEDK9WB4O/Bx1dJkWMBRcL
BByb+1TKkpdmGLfOYQtUk1VA+VRrk1Zapp9d69HF2eGg8aumP6pD0ru0Mkw8T8+YrZOuHR7mMyw3
ZqeRbPx/xesSmC37KMeZjY5TUwfVFSS7hzCocY9xER+BHN4AjQv0Aw0Ayn7ehWVHRzzS//+GDQix
FL1r0DpoX8YPOUR9u7NS2adOyfp+IfMPxbtkKMidMxBvJch985VUWjmhSuEEr+wvQXo03/ocadL+
Vk2n7yog4kigHgasxqcIZRGNXlwVb4k9s3LSAbQWmSAQS0v+6doT32Qk1lv3ce0A3u4zaU85T9Ci
kcOzkixCPQfaSlvID28Y+be4VJQMLgTceDHcL5q1gNN/20I54sYcCGNc984KUGrA/xQNFJZzpzoP
U5tSIuxuqVqlQksajNLJyAS0ZH4v4TK3b3amLEQ9OGLS4cFv5NBocI1dEObRlR4qU3E3ZuSC3ins
auyCfaJEyt/JFolfCwM3L6lT1Ko5oJ/3W6RNx2P1H+cvKDZu5ppdNx9fcmGvpUmXRgPUApKexgIW
qjrPA4Ni5EDXiTrlRUdCAlPGoKBK8D7Klvbbo34iLSLVF24/RASSyszkLaFdtPAtXWlPD9INwXrZ
+DBx0aZDjgogtN+CU9VK+ll+u2cHRjkj4XRChRCrhJq/w0TiRMmHJblGnaxVQmyvqiGjb+skCAoI
i75jQtAb2DKEl1j4e1tl6D3G+Cjb5XxZDAg43ifTabqlhuiLKAPHQNmbifN7cdSkzn3ghQNnHStQ
dAMx5J/Tkxlq+bHBipaUPCWxFIv/pCAge4/N3yfxj0IRizuGst25DL+KZQBs7RpRK6BEw4ReJTKg
Hy5HTbEXDe0bKZcRbeRxBUhwxrF+mGqX9hvXiubtrYpP+WLcAtv0LAU8k15FLs1NdsFo1fXY2dJU
w9pil6VrKu9s2/l6FRlZsZr15jCbNvHx00NbilfS+XCxdEOaXOu1O1auDNUGSyoVaAXYWpHNj76a
6XysgnrZEVuwpA3sCa+Z5Sxvn7E4Dd1QNdgSvOtOluNzzcRTCn5s82W83GmJrjLL8frMTOFSamTj
yQ91/Zs1sYOEmQETPFxey4+YnFWKhHBuMc5OybhnSGhJ6lMcT18SK7cSssi5U1Iu3sTrqfDXwKwB
4C+yhO7YnsVgvPPwjY5tjUkLTKOLrqrnVRiq1dw+7tgjYhz9iq/HPQ8gEZPrhrZqqxqoT4p2cvs5
dIQ32gV9smQDmyjAvPpv8EBrpYKCxdcoZBSEoguNBtEG1++zoDapB7gvPsr76bCGca3G51W9R/d0
YYHRyw/vSC3x/GnatyzQYgkUBg2lnGxEFcVL7N0C2ycSIW9clol2qs0eNTBUtr1Pw4d+M5eyswPV
2t9UAo6hlD97o1CAfE//beRPZeFbkp0njj+x+3y7GIqqQ6MqXHGSMrIFUlWJmeBOQqKI9CIcJ9rk
1RGyp9siXguAEkvHOcxIQu8jr0RdxYv3ISle6ab8hz2cOhS7Cvpp94pPhLmooGLYY5J+onaX8dsB
TjEjY5b7+O5/SnVjcWeQion6OhIKcSebYZuZ99RsL3Mwcf47ek2WXix83SmCiiTtw4BNNgcRkM0o
5X1NC7AyL2bM+VagPKcV+CtaTqmIT5AAFduhaX2VsjHshz0ANvRCPnlrRV9GNG84b5fNYUZmxT/D
Mr0TK35j6ojwQR689M2Eer+IdIqTw25NCd/wsNCOrL4Wd7+LObGZPum4RF49DYoz/5H84jQOg3KY
caUaYCFV4jm11r5UjRSppZItUd6ARg0q1Pj3Bsrmr0UcpYlp7rXDCoOuLipPkyg9WPv8ASP2M+1I
iRemvUGM2k5gCM19h4aZTyDhzjaVc0xmrTMAfOmQMG4/0iyZx7SUYBSk144UbwcjUhI0QvKTmKij
xuRN6uJGCyzLloYDFFpOCWgouZQBK+d5rB8aS8ihTxZjcap9Hj1wLF0SekJr0aGDZmOKa/egAUKw
kbDwW3agz3WyR0Yj6IZ8ssfP9HrEk1vdieTWhnIrV8Pmn13QhjzUH7X/3CdiMJmUMBEzHXxgcG2V
wfLD03vV50JXwgcEnRzQfcVxvPnoov1QGshdX+zi4NLLc22CrzSz64ZpQ+q1CQgsWELwXIxtDLev
rRfJYErUlK5tAKNUqe7P9OBeNsqZi99PtBZKrI/uWh4UsvLqseTfPxuW6B+lKb89AjnRDZGnAZcq
+ywnWdK22LsWzf9nB8t1Jvun+n5jV6fDORqhE+lm10OWGyM2i0AHTdkdd4iF4H7K6x9rJNwpEMzj
BR0vANAaxcmmUMpHsAenSEf7AnKL+iiq3dcsXBoQFGFgkTBv+hoRYq9XBFtSqLN2jTSp/DGALJrZ
MsOhIrlhKvwHj4vytwSg7t2Qiw9bNW0AaTg9reOqR3UiGLThk0uECUOsrDitwPViQcPofOAsp7AY
IL+CnW8pqFnbPI6ilu6w/wkInFGlFPjMNuCoNCRjsgUFIHJUduiwtdQBNpW0ZWM71YKYqVY4UrZH
YgwYEY0ecBSqHAx4FxS1gI/qfw2lW1hajtEDLhkwC2tVeAS4JZzCe6YqdrdGCTqrAMo3HWrCqe47
gMhymgEzEi0krkwUEk7YVGjEQ9HtZ/cgjjh5y5mLVE61dD7IlKNjZiopYaWEbICRDpPRH3c7Cctq
3LetwiYYqaDVLQ6mECPeXAg2oQd7c9gBqYnGl2Mquyb+BFVN/jfCurkncZYGV7ZodfRsdjObapky
5JgWWUYd60Zt6Jc29hBDZsDbDChdokMgsAIfkkdmxFjnY0Vj74wH7i2NpkdJdvGExvqg9noNEh44
mBgNMQbwCoVmlXEQ/zWT3XTl3r0KYUVXPlwINIttU69ymii3S/xMyHtN+7ArNzaK4L5gWRAVplfL
Jg/mAt/OPMgZLjkPSsTh+IXY4cVgTF7NIOflkLIkUsbb0gHNgO6LjJR+fCzxDUqvFunFsHLstI8t
XiRCkxsm5NNMeDxyYCr9dGiUpRs71JsW0U1+LmIUaZna9TavpQ2pcl3F/2+zKK9jzND1IWtaxHwz
R031hUTVYtSnBHRWdl2Kq3uYKUVJ2eWqZTmyskHziDPIbPimgKH8mIhA0csBHvIlP0oukry5MTfW
LrBKVQmuBxKwXuepLmlHfiJgHQk4EorT5lbUKSS056ewFAnqTVzcEFOItzXNzYnHxdFlHSkMmOnp
HT1njJZD2OBsjwchi3LY757hX4rNpjDyKU0s+7hReLOHv/jUGt4mMQOfKO1Mg5dyg36RrWlTLvxn
plZ8tfZyIktQHsqI716F2PK+WWR1YRC7k+G20io+CjImNb3L475CE3v0gqkDqfyKWxebWTEkuPA/
AMva9/3a7ReL9WIdZwBOzFXNlcFL6iFsRLD46sowgAXWw9AKghQSEh6jqXm3rmcSYqjbYhtX9vpS
SuCjxGPVPTE8k6Q3wMpDKSDPRPCR+MGMnnGms840V1aH655f7e3wGNt5DLpo4CJCv3GnkNXglq7V
xLviKbDiDI2qhqDr8i5lO6guvGJJ2fksLW3Aiwzyny2tqoYALJgLXkRUAFu+z+rS11dW4RLlDEqV
6yUmcDxWFWoNMV0iBBHTEAiqJF9xNzaBiMkDvzvHyZy8qwf28A4vj0vuOr0e48GkDGHMvusCbBcK
QkuuaA0oPkygwcUAPCBVsm9Vi8jRAq+CFnjBrCD2j8IZXmhwS6VUANcXfzy+jJL0C21uXadSIRnq
/vM921uraHlIWNZkVucG7umXjRHX7HOIHj1G25oHxzdg/KtcV6s2gr/ci+nJSmgb0Mz4tvnja+6j
Pf5y9Q2XRS+HpoJt+ZYBUNhN2SaAttee4Av9YteZWF3QiV8cGrAQ8C/iXfBOuWxIi1PzO2j0OATC
CfdobhM099l6v5/kpSOAHZMnixXFbofA3xXytVmu1bdKm4RcK0cfeHsfTlavZsEpo4zuYD8Dkcvx
cRVO4HIAwCOS8cNwRY3EkZOfzt91YSUTcrjKNtI2mBpD5XCwkLizhYbLSj1i1t1jjkSnOoM8HoZT
zJnqg6uFqmNvHCmsnZa1njvp9dUh/r3Nis+z5hK9zKaWy6cDbH+g9HY0ODjzk0WFMWsUVk/PDjzf
4EIxBmQauW4/esbVnaapPfjdxFasDyKfnaVM9OmsjQyXKEHBFbL6qyqtcCnePFWIoq9zffdBW/52
spqUgRi5hKDUM1rXXI8IHVFuZw78R45AbcRveR0elGBVyyez8NQz6v5MjUSbG6fY1RaUZdgK85eo
gRKfOEhGj0tY8WboPu+ULRN+89zCWAyk/x71YNCJFqVzPQ04KGNrMqL3O6hkl4e+L4W47YqGbsE0
JHMFjh8yqp6FNKq0WcVKM+JNmmYngqPsE4k6swTLMHfm3JJfv9WuGpWiAK/ynzsv1kAau1v2sMry
IQSDoC7ZQriky9T5aXxpfCEuZt9M+mo36l8FBjCFt4trQNHwPcp0yqv64K7EVauQDwGdXZCa3T5b
z7iwW7MI3xS/yK7CEZyVAdshLx1sZY03IsUgzRzwbJqqZZKhCWyNdQPlQ04FOTMdtDeVK2qWcXA8
yJgDQn8Zn9OfsmbMgwUvmT6PbyC4uu4WbJSSqe9Q4HqgiR5508JeJQVInCcrf0IvKDKQ4zSxPC98
4Y1ypS9k4jAC31cfuh6hDw9vijH17AS0arUrszDDilP8PZUmg8hT2b/du0SQTmjeKs7XOu5l10Am
ibCv2N8gfaPdOVDI7WptCFFiws58EpZ1PRq3FZhtbFUct4iMV5N3Sr0SBpYlmqc3LjMkoztcgUgd
vFfcFE6aAdEHhMcseT1yXggaaI+cyIWSP42IqYU2zHuoCq26ZpT7raZEKXd+XU9OuYz3t0i7jGca
4Yuey5pPJYUJvjshfdyZJBwBo9CbArVaP6/ojwAPUBlwg1fuFI0c86E3+y+sBjWRmbKBIcVWH3Q7
J66ww4O8dqCdFIFAgm3Yoh5EqeSC3LQt/cZvqQ1LdOgxxHtZAckHvuyf67pA2H8j/2R+3qBOymnz
b2vAPfoJ60NNRNUJFYj303h97hUdozQUhqS1HqlrHYEbyIupTLAVLes752tsocs2jvNshloAwSIw
VjkETJYjzPxese/yNLsfSiB91rwxAYzr+K3CHnJXAJYQxTXDjkqqxRy12rV5oN19j5yd6mI306m3
sGOMo+mcqDc4/hoJORy/+d3YxUxm4OtcgyKmep1lp4ejMdvunTa3tTwZiaYQ2pL6npHvYJZqGlbf
nEiEMYPIW+38e0/O5pdOt+p5DFOn/NCoUFFAewob1xjDVUCPpogTY6/90J9A5GPBgM38vsn1fB0M
QSKuhsK67BbhuCmAmc7Qn9EuYMIHam63GPjWz5zaTkAnf4L20kVF5aWFkX01VxwLOmqpn4UpF8Im
sQLgaf1c4dAJju+35gTjDqD3vhYilI6eX0oSNaQlbi24K7F3jgMxtyZE5UDizhiI+L1G+Omv9lbw
r29npJyON301FBrf/Oddf/jJfHqsLuU6sA7r5+BS6l/iOrwJqL6tQatXFZuKG9QnTVat+8PnCkY4
+qocByf5YfyimFnmtoEBdfCDOdjliYOMKp9gcf3YQZrUN4gOXxgkiyMzrMfa/HC31ZnwCON7u9O3
fkdnI2HKy4ciboCp2sjuRwytJ4SOA/V/KJaXrwfTG8i29+wZ01FcE9PXEH1Q1edrOpJkeffH2MvR
W12twtVsoD0izp7u/Bw9iZTyJOZw6ot2cLlJRicUENzj6XygBsp0htcBYRaFeQ98nFioy2/qNU1Y
Jfp10hkPOT3F2Re6C+5o2n2ZJW8YaGMBs64YCGNyIZxJRHdq0GVI72+bllGz85CDpdJFOyln5YjJ
cBPSWWeeV/W07mHUCAwEr2FBq8hC9wOGwDsgWFf1Mj5udgmcFWWWxp7GtAJEs+LFMHkIpI0otK+7
GFoOc5kCej7DhZ/kc/PgW4yiw/CmJkEvl/pIm7mGulZpExGyygGAjC1LMIQTn+W26GazNrCbqYxR
GFtQmg8tgikltpaJWd14MMAPQdwNuBFc4nYMOXXjX4/ip2zOIfp0e9X2u4PO7ZPuO3fhqwm/Si8c
lgCadOx8Jil5HxWyEcl4lz1jn7XPhXYuuxbMccHvFBXUG3dflm3S94mea/IuUqq+agvKrWxojOFj
FDhf31eRE6/BJm3QsxqTYfTMMJlOMpmvI51ommgQyU978gX24+4ydjtMv4sbWtiPSCTBM9V3usrH
4gc/+zAYIinmQIvglAlXrqOTYSp3wsp5gjOW1eWYy95ToIq3hHZpQKZ5WTO7u1Qc1vw/0q31LNF3
VCz7nqHW5j7NOygQNyKVz0wW+EtVph/5AgP1fOnYo0jHuY7RhUlfP6JMOV7TL/bWFfwSEzjgcnBW
jkGJDCNc6tiV7ksl13iPxY8RNho18jVYqHx4C2gO5CVgRc4VbJvrsaVpKDsZpxVZU/T9pWUo5qWb
m9GrI1hMaWEa4xOHno9XmnmmiASZU5nVcCk/7RmA4tb8Whu+aCRXzYJyvlk1Ig5qCYfLHlzOphd9
fPE3o1W59V493i0gE2SsmLsF9Fs6UMvxXpV1k0vY2CnYoXgfzhSBimjIqj/g8fRvwzOhgUC9EJvw
ZtFDG7+8kuv+7oQqn21NRe4f+g/tDky0624VXFOtOIvk+6LNYC6+A6F9+N4l4KIMofi4tNwR62At
DCukVoyq2Xr86KQO/uz1k3ij6Ym3bFwXv78vDdZ3i2m6nMH4Y6oiQ/6FPAUNikoR5hCrvu5VgIOJ
zhvmSl5+jWMhCOWf10GsWBE2zQjEAlDnKdpOyk6IGoU2o1tNmqE+mHJ019M4rHhGuN+kTKtt2Wcv
gMtr/BCXAtKQ82+ojCyspMKBb382kjB4sP0vIRLKjcG7Af7a+2RADwkRlh56qd5aRdn4RG7+9bHH
gBDWDhXQKOrqwFM+bXvP4fSa3H+J3CM57/paJC7yOmZd8fd9TKiQ5t/BC8kdLs9+K3yGU47FId+I
8sSz/HQuAGkvHI2/pNlTko5C14fIWmM1BgkIyMP6z7FXGga49OpVKmQSC/fHfbDkzzLuQBYYaiG+
giV21n5yYpfrd5i7FdcgLnp569FQPz7O60symkEW0AXNXZzTDGahSV6omNfpP3u+JJ33bOrph0ao
I2sQF2Qrx27dpyiw0VpkX0mNY9lNwlDnLYO98iodBiR8pHbNh30srrXEGx0dZps1lCQjUW9sNaL2
sUUiOXqvMahEy+MVktgx9LtTf8WZ8sRJ+/CFI78IWH6qYLJXnQq7WiOetEPUCOEJ7tGXTI+zfsb/
CtmPe8L0KyTUTOGzOUEbgWJMSCgVQfqWuT/zGp74j1SO7QE4dLdrKBB3mTD34PvjwZxhvwzBmtQa
ck2Gd0aLBtQw7SwaAPxWvNb3GjQewJqAk2gtO8hXAaK0wk4DPjoOLRcVbmXFxquR1u9oqnepUpJt
4vgYyv23P+uTxhVDZuVgAlvzca/stsELhxlQLRH8Mnj3cTMCcWy7EVQN2DrBI++geh33SeABvn6k
gIePZN5VX1UdEvjFaDGZgJgDZtK04TEucIZceTSVdjqlhzlgFEpN1J1JkXkFRCKhA5OBXZEXkCiE
rrWq17WyrtXGB09/0seU1m3XEh+5sRBH0lkpJiQhwN75uZgvHebC4/lw2n1HbMcyOHb34oAklLo7
MjGa7/bzmAAJlSY05b51g2EJ6/pRBphke55YQKhHwcTkvmzoo61sutyKUnO4b7F1SF21Q9IDrfNE
wocLKjYT7U/NvtXI+Vq+EjL+55ZaiqlgQ5LA6UGLL9gbb24qKTyASoxDFPhut30BGof03YHBXbJt
HBG6VSgche2WYgT/E8W69Z6+FDeGpju0r+KNToApggQwOZLrYXszL1bNJ85r89eQZYTjNUuYRq2P
hE7Tca8JN98dO806kBoOgaFa7sd7LHU9nUJPQJEJxI0DBEAbo48emfgUKkk41WD74JpZP7uPQpzC
ummESQ11Vo5h8RQkkX90j0ADgQr+d/4EtlIX80zVjFGE1sj6mB4PIOy1pBT8eemwi6UPRQ/rYtVs
wA3qXHzsnbbwdD4uadept5FpT5yjRpz9LgXi+N14JrGnqaczg0oFg7DRTaAY6mihhHXWmn1kFyIS
jMZ0jBMlV2ACizl43ULXqE4Sms0cUDeJjqcvwSRA2B8Plm/YbbySQ4zXiNWtEZvBamuOCM5A+c2a
vW131kgaiNIhTaOS/NHnIg9xC9/pz4Fndfr5F8Wo4KL2fRgnKcRFfEiP8CmNpuX2R3TC5TpW1hER
R+82FzFgt3ASBT9+C17nts4QXnZJ81+0w51ryqiQhJwTmjDOF+9QgeZtvwtPSBTk85s+IIhsy7Pz
rNs7177mGGQ7NfVR40Qvu1lSX6wDh/R63VRWth/PH+UuowwnoBlbnoy1sIHuhHNW1bQvxjVA0OFH
mxg+ErldgsjWl2xriDehpH6/LunRilfjyXbzfrH2CR2vOoQhHI5DhA7dydBAwWnfM5XUcs3bgEyE
foBGdrRuIC0Uw+LKzDWDpVfG3obMqr3djOYAMNG/5zaSGMoMwEbeS1YmIjop5JBeeMWtHExUtTga
MElCuaLBV0OTJWDWfyMEkT+ZKaKgYpT+b7fgF2fN/Zta0HGvTx/ccY3t76f5TEVqVBjrMsVOKjkF
SG7EgosU7K6LyR9g0JDti+oQcWnlP+dlANuJ1ac9vaiwdauICFbnclNc7BqxJDHGuaIe3mpdrGnv
utZYoPUtOmHhgZCjJ6axSzUL+fx84KJjAE7bDNxBzjtno34hQ+sOxZdXQA67OXc9VgPwaMxpesUy
jP8LMylDgRyxOVR/S+Wgv3EMMiF5snHYcKe/VB/7Sx8OmVaaRSZfcQv5yc4+ufqJ131TibQ+NOVq
NAanoTCeo+G71wcGR5GRWSCIVpqv78nyf23uprS9Mqvmm/6oKDu5XFruOSpe33hwaCZAsgKlnoaL
2t7979yG8sIDT75WjOw96FI39CC1G1gnLepRIPvW7riZHO427D10ye24Bvjkv1HiPjQLAB2UY4lr
Mr02aVtmtmIqUNjXz2eTa6S8Z9VO9melj6+x0FokW+VX5oc05nBZvwY5BjXcVou+wz03r2BR3j1w
FO+J6Dm69uHZkIHAhTz80I3KTeH+3rQvGpyjSt2cRQto9OzliVS9FjN/gVr1K5zme+1bcARYCmUf
5fOKJJOXNKZXkutf1StyZc7jjsIPzhRHC9XRFDi+nAgTqJMBTk36f2ezPxE+Mo9sp8sAGMpWlrqL
xuo/iF3v9qXZkEo1SuY2G0M7TSYjSSwnkVG7Ue/PNWjPLk8qpGq+co0lksZ7dUzm6wyeUDaFJavo
I5LyxTg7Qq3Fk+BIu+MU3SLPGlyrXD/rOey7S2tl6xYE0OgCepy+xBOfeRO6NtNvnOfzgjMYmIby
lUKVZLrKJ4KgLLUJobBB+5pKHDcPBuDl43/Z1AcAiSBbiD/LXA3Y55WNF9nv1FBe+L3t66GpKefT
b9MuBBWhA4kHCuWULrNbC6MKY6yoX7okD9RIA/lQQt07pFQZzd7W9sPDpcGnd30bBWMXcZJd7In3
Bn6jwCn5Wy43USg2KO3DGBAIxhd6K11Yk0S7dt5EFmcuZAubYUo7oUXYJtJtqRNaUZLQVb7Tn3oo
BLu/KKKgXa65sfbeyvBBGZqRUdXTtVeIkCgv+oHqSfN6lbYlSlo9OOpoaG299AVHNXN9Gg+KNpgI
CpY7ZSINVwJPOPRS93eTy+Ov4cU2EoRIekvvB3k+AAolsdYOeILkP9p0XtrhfdTL+viJTH8NL5c3
NQKScy+L+oGikCxmc8PMQyNo4GM48Kpv/2hjp+bUlJQS/shIQ71ICU2Vk1FGeLehVK+5ULhR7W/R
xBB0X0nUeWJLxn13XRjChNKQWrXGvkPKIX66dSicjad3P+FR4wbSQ+8FbmKdqhJDbDf0dB5UplrN
Q3aMafNcHlyiSZ19sS5KFo4V4j+cTIYBqVrFX2/iOsELcVBFmjgU6f9yM4jm/VwFIo81fZEX2P5v
BPrgtaglduOun1pkZxhHNZHHSnECOBMOSmzs/Vo0YHf6yok/GPd2Xbbfr0pHdE9UmGuvvqgR1dTq
ZzGn2GPRyQMK7VNL46n2PNAot5LXFVHlTaC28YwfBppeyKSwU5R4gApmF1uDR63NJFryG6ZBbwem
NyjXVJULQ0baR5nF253YSywozZqSv9APj9VmX2a/N5CEYGzyB6tLnaaUI1jvt8dHNV92CnZP7H5l
vIiXqcHVc/U28+YtJUjPCHX9zbjcsQ+sJKq3v6RUH9WLkK4Xe2QHmDM/5/1TN5D0jZBlACypLXfg
xU4AF0lg1nXR02LyjefEIJwU/dyHUJas7sx2LQG2lYV8bJoxOZTebZudk2pLZMI0pUv5HCREy2qT
sHcSJ/GchrSTeItmYEKeYDJ5oQ2hnhDlPFZ+3d5rSZs5nyQjJn68kMXk6/0ESLxJTCQD926b66N/
g2KoRazKYj98msKb5n87tlWIBYX1enZGuxfNDf4kMDTRpXVuYDCuglOrt7ginK8l/RhtIagzOuM/
wK8X3oqWTfc5T4JxWkBGGf4G1DcjnqouihY6uc6NAnOB5ucUTuT5+dt3gmgHxSIIe4v+8tzwqHUk
Xsk5bRp+gZLCwN66wjnptav7hG+fG1yVW32LHGjYV2V6doHe7V579OUePxpt+NxoM3aiLeBE4aSc
ZKsC9Hn3JAJUQ3eSpgS0IFen10XMVFMl8C0aq0u+tok2llsctD0YKg/cz8OQOWnBzpVsdABKFjHy
Q++vDCdWZbPNN6D742A36VrjxJ3G0bhL+FEoG5h7sPyVa8hfUTv3c1fgju4H9UPQjteI5l3trPaB
sqaPEa9jUc0rSGxIJa2bsJyN46uhteVRIqlr8EbWYr292PFOWAIS4OXX8Ek2QJpwNJ3qqUPsPsej
rfozGcccQAFHd+rOJq8yMkMP1od5G2GGSRELyZbdlKdFVD6mjvoC5ZJVsyehTfrAiBH9xK+wVRPo
ffDNNiruHhjTCxknbY//z/8ygX9NjhttJ06ssb9H4ah8wvDOfxsc4GWbzNFLXROEYyKVcOzBaSLC
E/eZFmTFDNrbAegrbD5rigiZZtdpYK/7VBrxzNwBWMv8UqlwdeBUOdBeqrL/Rt8zECEGkIPvLtXx
FTP53W6IHRKVkYCMQ2FtyMZwKaOKjpiKMGc084QetPIZ+4jSN9iPR4eASiG6J9AQAa3Iowl7hgns
sR5qp9dK1KVBoqVxmFyM0AxH0gKaJYSteBHYvmkyq87znoFr3T/mewfgihBCwic7V2JeiTsiB4ld
oWOgyC7bplUzjEJgZ0AotF3pi2s+FAD/jDjAWNdcFeXL7Ylh9us8zX4J9eIdRU2KVj9J0oO18DoH
jFzqUfvqGoAIT4ozufeqlayKEp50r+ECnPtQQB0PEnlJE7kM77QDaFW+ZOh3kT/s0mxhN7UdLZxE
Jq0CE9txUbOiAolGVK+ErK1lQILgTNmcjpLwydcUHqEZ8MwAb3Za+F3JurOuO1G81PVIcP6O7QJU
RR6fNfLmBlMnTYiKWOU92u1jA9ohpM3zq6bvSXYgPbfOlBTBQvff8pDNlkIwsgZKe3Jvwnc6u88q
YwB5SPuIgoB+n7/6ixDpRZ3fJp3A43hlqJCPHuXOOZ6Nd097ToGqWhVoJAna0mIyFRnJW5ctJiaD
aDyTsRvdO3qqKkoUlZxLPSG9OtobALz9lMuZwvL+PWjPOx2lK+EbcVB+RnI5lPfPsQqQt5wsHKsJ
d/TK/xwLJMfZ90U4Sh0tu6Wjt1ExmMqHexRYCTlwsMRf+3ivqGpJfABPjLWXKJVub0IGXye7s2LZ
DCqKlsAYD/Ju7kpzuZOIDo+8MjwYxC1j/qg3kgSc0jIzJBMRbjdPsMofKlg+t+RYtVdPb6SEgTtf
bET27vouq8IOIUXQGO+7pSkzPELcjIT//J5diYj25E0+JrgBw3hKM0ksKi9CUdrzdSPMcfZ9rIEU
y37q7xYb6SaGpmzdEgVM+G3+Wx2kk5x26LL/xwX2X3BQ5ZHNHZUGuY7NhMuAyvzgHFJEhyRTQ3e2
msIdxqjtazusmyAjEHqeOn24NymC+/2eOncVNLZgu7PQhOUD8czkBZnw3oUg16fDQbQ6R51/tCRH
pXo3SfXN4X1SABAnlfW1xQfksc1ZeV4C8Z6ZY852DoFI4QWFQDZP/anmHJqmX7v/Bp8Gix4A75Xr
85iyBgva3xeQ5TaNjH7DXKuhRB+QVgnu4HLP1ogaET+Y1Cd9SgJ2Ls6zkm2ZIFaxJC6Cx5uqxV+H
DlX8yGiaFveFkyomJ/cikvmKLLuTowF2ameWAUAVuhiZs4OQayZKFop48eEYrYup6FSWhWN81sbi
u4/NrTukDooBTVYgBhso/w3O82QTQO+o+ofPO2hHxWEkqqTLUqSuYKw4TDjPBLHkfMTGy/x207gS
PH48NQ0gbq6BbJgv1NXq+ZfKPsbGMWdLx8io3AEcD5QpOfgqo9byNttqB3zUwO8yzBZyU4IGz3zL
g6Wh3nKuIvOU26Hl96ToO44CJqp/xR9Cemiei3+YgXZUGW++IOlOeYiLGe90HWoQ5UjkoHK5Eond
qEkvMoYaJ1aueCY48SLVtaudaOxz4oICmvyH2MjgLoRGEor4azkJgdOswFwDtpkxLRDOqpjwHUys
Qf81PbMRLY+4mr2O6oRvHbFNfZMAtgXQ/4I8TU8GuiiaGrQrAYXhUi/bQaitZo3F7BP5HqgCVkEE
ye4RxGESdAPR/X/Xmn9wuYvn7RAtWyfukk0x9LWBX6/CraSmyCT8JdrHMfp5CpOWuGG7lnxyun4C
XJShF7KWsL6keY35QlAyLCT3JLz8ha9iskAjfHzxfSHuBH2mi03aGJoOq672ma4xF5qGDq7yxtzz
XaOmhyJ2l2/lyMfPNdEGo1VDzV9eO7qUe6jkjrV/SmbcmGYAOnsXp/aR9UgHwihk2wMR7zdrxLqK
wDmEddachLp2B4r0Qjk7IjbhWh41GbBROxO+Hk2kb16YG4thZKqRcH2cyIHVkjsnm2osirFXbXzl
9zpNdERrLCV1ANw6KLon3bLRCHIzXXVHlF5HOi00DQJzlZl6YOjkeG7Z5LZy2kxvsYrL6bwe0W+L
gghFxF87PlHX9coqVNOhkVmVNgMK6qhUgd0Z07Mbz2D+PtMnv/zdfv6OSBxr8ziBRjdppKWJ7u+U
kZEkHaf8j5iW0Ku0cLIGrfb2pUL4fm0IM6N7Colqfbgohv47UED9in8B9eT1/Y+qHQjH6dilSuYY
Dazp4D0oOF8fOs0YwiFvP7veYUvEonGNAQj6M7p4vuXJGittv/7N9+um9uBFj3Fr8+Ty7B7o7C6O
X/+szFg1nfQDyouyLU6bGekI0KT6EoFQp3LvG8135Otcj53gJrkp6gHQ+qrnKVGpF1BqAWbJN/Rp
39eqNzuERlqVwkwqNIUgRdiJfYyiZlhLHJxo07Wjkx/wdsY9jxoiptTxrUTct5RJ8P8Yee8mczZJ
Bhw7wrqkN1DSekKUCf82FwpADNnuIOWmTaYgWcm1uAj7UIBchEvywsQQ9lZRvCfHeuopjkZxjOQy
TZdweM/WJI8cvIrKXbFh6cToZNKmRUXYEZCmjeen/+YaB8sQHEc9l3fa74HX0fCkOSfgpPvfpmSJ
GSbUszAY6pzlBi4hLmPrsQgxuAb+dL6RY3XRCw90wHEHzR7L0Dbx7IRpXiOpp02QXnth+GbOOd/g
0svXUzFlam/pOkynT9kbu0dF6LDc9AGjxMtE3Y/WCpOZzZwa7svy0LdKlBXmb1SFSNdEbCMvbvxj
fljP/5veltTVz3IEZCWkG0A+q8V9w29vVPPjGXNgNlUQzSseVvhMKkTYCRkztUSFOe2DVEnw429T
3lyn4/AIJB0sgn+nsUsKJ3v9rjSxqeiUv3q5LIz6Y4Iebpq/sx713uwKufWF7GRpCDAVzNQo8x+M
V6aNWVH0ujNh+3bWN/zJGuRWfv8Gq/Vs6TC3+A0DS9dZkXSSMagQajLhI4xQENBwThExGVuxi3bq
48wctEs42fM+pfzCm2VL92gYMb50Rs0iaVJ8iYo7WyqVLSRpHkNsR2DK3Zlk8x+qEejw/FirlpVP
/xQ9pv9x++osHB+BvFGvjQ+eihVb9MbUw8So6rjcYyPwgSVgRoej/GuweYYb7JuI9+x/ITahqejV
q7FDgpZW5ZPzie+ZdTvhaFhzw3q6UpqYsLFh+/IHve0tA4/uZNsJTvdeLIE3GVCwAtDTY1cKLOdA
IyyxJBlHFmOLbrtxWC6cf4CHHeo8pHKvczZwgz3VxeyYiqiRc3qVD88Y+8W55ie9CBb8gHxzBo96
eQSzfOpqZMGKxz9sbmY8VnRAw46cODNc/R42aHrGf2An0x+BrfcAjpSItGEa/nTK59EeFeisZ3pH
SrT2FLGw9oXNIP9PFXwS3TVe988+vc9uzPZBx+9NwsFQzZwYYUj5+54AQL999YQIKZHVddJubWXB
7X5x2zBZbDtOEDnpNQz5ZyLBF6lnwZ6aYr9Q0ENdtz1N0XDUmLHZaUOFHS4t04Y8tKuQmGf9B1rb
/bN4H7zxO5Y6MM7JN+c6GVdMstR18LCIPz91L8H3z1XplJbcH+pia7p6JBzjz9oB+fGAAeKqmgXJ
1AQsfpm2U1+lfAaXLZ++oRjRe5quM10ZR477E02GBj6yHZvrjKIBJrBoOYFi6+KjJqXxB+CZznEk
iXzQK0XOD0x/cnzSIsWOiIbeNdWBxGunLRzV4lDIUrMiZ6QRH11I/GFkyaoyCtTU6DOjFfXS8+td
aqqMgRCwowK/BVpBc01TpZlMXf/kIb83zCtXtwE+wioH3ZXw4FOx5umBWJMeYjIgy2fKLIyI48aU
OV0E67p4kzugK/z1pPoIAgwbfabg5J24OoIHkF38eP6OXMixBSOcqzZMv/SR8pXcjPRPVHSpmhP5
0qZzQwyLfzoOzJC/r2fCHqzbXCCPUHaRFOTqvaI/QSrbFjVHKxAIFHLK9mW5ZrbYqDwicz05MIZr
1aEWu8eThFiFtjVWD94c5GkadWXKEMSxnkxJnl9MdKRE0310tkM5qSakrEjV6cilY6Mt9RJoqlXN
cX57PjiZES99cXt4lMcOesZ4D13FaLbuyJEnaiUXSVgUYk4lZRwid7P3Z1eSwGXBWuUL6K87Oy3M
Mo3sjjhCKXhGUdIgsrpF1IC39+aY5qvL4lfH+fDEbN0g2YZPhi2RJuhcCcFJ55W1kdViWZR9vars
xRiQ797FDv8Fmckk4AtzJDqi5JCUrlsEmMbOyBO7sMtArvXrPKUajy9V3jV4M+OLGghPwVgBjxNd
my1iTDe7u1A7Aq+rPZAVhWlsMz6e3fCV44i5FDkS7F/yEGtQQeZeJWyMRYEG/6XAwJbMD4H895YX
AKcDq0yS+2ZpzmX9E4gRkGuc/xNLduOilkjteB8qTq1DpwYnXcGKjbBA+NLC5xtkxWmneV09XObt
pYYUSQtvjaIDt+kSagDajHyLVT44PaRK3n4e5LwKCfSBxM6WxsHR50vLNAKd5B/Wu3KPHw5Zur3S
cQ2IsEpvo1WCNAAkidxA+UUd2l3p0Eo6k0icSljgeCf2dgHLrUStvPajUDZQI55oRnpu8ZWhBUU0
k3Jb/Mb9cVu+cIoRMaUyF4atHHpjinVTZsEe3EtXdQg80J4mVaQHWuodlkFndDyTfGkCLSxDv6AJ
J71voL1hFzbe5k9H1a27wVlS/zy4HY1/IPXGvXCuwvWsudxuArDvb3lcmEcha57y2bDdqOMS/7J3
j76PggV9ti+GnlWwgXBFHe7yaMfgYQcNDqdRfudMfuM7IDzjOa/DVt+8wLN+Qyd3bTgEK92XZ6kq
VN3N8K0QE+L1NoasLbh2EmMJ1zpAhyYtYB7PJX6fyIrwm0uE9e/K7KSyVfFDhvgSACQ0qPk/EOJK
yKZdKdHmFrah28edbCxBUC3n7cF5tvKlMLqxBlvMSGr9rJMlPwRmqisgUr1kl+aDeBvX3LyWn1q8
293srtxpLZ25T3FcyUvTsgCuk3C+S/zEJ8/b6zRYQ23LXzxh0qn8I/OfdemN5YN6LuquRxENC15q
9EDWJgBLI+NMllemBmZEb0R8O0TberW/HVMgAz3PNn0kVNcl54uNfWnvIiuoPWXpoNB1GeQqVjgQ
LDLkOOq1jr7UpBWJkjAwDWRU8nhakvxb/6rb9hlZtlDydvV/HDTBPX2SO626WolVysrF7dcjT20S
vZLKj4UevQ7qL735noTyPKmbzBFqSi7hQlqEltqa266S6+spKRXeF/56BfqCHX6xtErsOZOKYw5t
Vnqs5E4VPYuih0SPIBWoisCecRyGYV9cU8BvSPJgRgf9XOuFiocsCW/4rzcVYvsC71QTBXs7x0Ix
69GyYmoHxUMAeaJaZ+It6JQo5Fmm2oWE8kE76FpQyqxZJ5Wp/bfi+9D8oJRUEYeoUSkJ/LpkOSI9
y4MZ6xsVlg4lJfw6HVE0JEuQMjXbrnQNUzo19Qg8SoPU8B9aDeRXroCqnJqjPahPdI4hW2LiwpJK
uSry9IUm3wPILl0RYzeot+iZwA29/8tLhm1Z/CdiJw9p5czqR1XRoH/RzdU55C4VUh2qCiXZmw5k
Limg8OWyCMW+tZPH97XBP+XCSGFRilFB/3oQMG/Bn0w3/9sOTiqNztBMEB+smm4M+6m2fjveiuWn
dePCw5pUl1WYo6hMRBtHSfGCkjty6lp+eQjqZf3K0gm3D1MDTL7MXHg05K0h3lrIMPmHgBByjuye
TX6+C2ozqyPT9I/mU2LdVlw1kJh3jHZ04jUwSIS1qDayiIk/rz0118IsHyMgd33g8qB6ErZjrrwL
PXiHfDykeYHSqHrdFgCXwmjRB/JWJVcpmiRI652xO9YzOWI4tddCVFHGaeA7byuahVjILiISs8jk
Jt6GObj2rtAo6sNpS6JbpNdj7vSO13NM5pREwPgiUgJMxxK/9PPOScftMdQdFHdPWQlZ0+SEzqqJ
08oBeoUbjHeUnoeGg8V3EEpNLGTUvfrbSRCbv8cKcCR1be04sgT824sPwwnNMY7d7yb53EPLCO2F
zUPbBj30Iyifl3SifrH4Fx6a3D6SJ2WL0y2gP7ZIivC9QyCntxuJjk3vurR0iM6OfczoBVMJb7vh
1XWnpO2Wm5eUO8ht47UZqb8VtUj0oolxOjuNthTIZ8mE/EIVfupl1JXXOEZskpH1/ffFZsEhT20+
9298JVPKHEXAGYdIgdPHtJf5aFrtFP4LmYL5fBhR/J6prUa40Xcccq7gaeynAjz7Be95dq4k+c5I
cO7Hu8tfOOMa+1vYU56+b/8qAZwjdooM+eI0OljegcP+c4NWT1+B0u2pnO1i3PmPhaEVJ3xLpkEZ
7tpE0nTCw5ixMu9qFPNGnypk597QhVN1/EnrlNcC5GneHgm9d7Qg2rFR6LbgR0R8rBIj1gHDXqM2
kBtxl9LZVn7QRWRdrNZ1xYjUa4ur6PlAsTaj2WHBcEv+sCq3Ckiv8rQPAs+DC0kiArvW8yqsDN46
VnUJpGpWRm52TsXTt1uJ+0XO5QE+m2XU8FLKlNVi/5Q+O8esl0STYLEh2u+J5LQ6NmStPGfIO+TG
/1ZaSGukCWNAZLu7GCyzDoQePjcI5OFD4GUOuz1vov/Uh1G5j8UfOg2r1QWo4dmr7pBThqKfSYZ7
c4bKJrNGHlrHQGEP0IOMbUwWj/ptaXW43h8MOFsGYDVhrUyrzJM3mqg8AGo87NK7DZcdmWHmnzWw
6dxLl9fX3wVhPOEAfjwmQLkcTXE1w+Vs+RZA1NQyxRl07SfHZUfLOfdO9JkMgxBRCONXhL4rBccP
R9KHMhm06542g4GJqe0/etESJUKQDhxHfmtnCyMqZEwG8/0zMhDZxwsl8Rh5Nv+DDAaJrDvkBn2b
vTRcx/smcnwDCkFtm0/MuPnceazWOOoxoECzq4dBqIZX9NJhblCL3RNcJM2UF7Jco5IMwzEjqt7l
PtSJ1l/ZqiQuUM9Yy55pkksi75LO5FsPZJ0RAyEQMrt7VEzSzymVtR10pJ5gpk9OdcjpEt8LtVd5
GCjLqF4Eddh9UeG+Q5j1k9td6fUxMpxKg3/Uxm+4QGAW1WhOl/gIaoc6SzudQtjSdi7THImtA6d9
rBEFyOKBJNh5Q1z8ccUWUbvgPQHNQB0YCDDTTxfgrjV4izmwqBNH+Q6QVHAKV+qDcXbiFrY2EVOG
KfQ0ywxvJ43Ccg77TV0A2u78SKfJOijfzJ1u2AAoyh45o9TQs0dCT6jrgAhV7iL9CDN/W4UEN28w
Q8+LFDDNzsd6neHq09JXR/Itbpef2/EpsU4ew0bd2RlN4CENVDoftB2X4eJBOYtXmWk3uEDmSapv
0x/P8ZknE3k3GWuYPUIZ5bJOsskf6CWaYP2/8IUoZlJW/XOpc++0h44AoO93dQispWDBTXippmxv
3nPSDl6PJA6II7sGGcsyskyl9gL3blpRJABQh3/TCIUuRMu0g8v/AnPZXsmN3I5pIoUI/SAYcWcN
kpOvhxK1YbKcH4dUdcnNBP+3+ijY2kqbI5MW8c04EzSBy0RjtpIXfmlYyUldbvoycKlimVkYpKI5
2vjtWgja84MLLjC6t3Pt3t9tiZhxWvzHrh/XmmuhI1u3gdfvcz7e8+2OYZqiM+0P0doEb2s05y0o
vXnpVya7r9bVuszKnmqMFRqfTVlT47k1/ririrZjA0dfvSZCwOT/OU3Ygh9YEmH5yM1xCuKhZTkD
bfr7AdFNshG5ZswpjytblbD0bGJ/dyq6K8CR43n5P5opA9yB0TYZoPbWU9AGwqnUh90V6se/TTdc
eB+cb7a7SzXHjEaKBeKauAXnnVQhI03ExOY4NEm2rKdrrPkEhloZrB4SZJ1kFaExJn3hbuICQDsp
rTo5e+tciiCz893AQTw9PuPWwuNRLjLC073rfqndd+514Gfqk5xNnB+3EbnkkVZlnybTZ4ksVWY2
Q2w6Xc+Vmq4BRGkaFSE7CgcvsR6gIfcNBDWEJJ6RRXRw/jqN1ZOZS29Josw5irJwWF81AxQcf++n
HBIS0y2XTTmXj6hcLr9tuQrB9Z1TssPw7NhFj4+2agV3faFY10wf2SbVFSK3bxAjmczR3RjhUDY4
yXtxwvbO8osG8C1fucLBMS+UnVh9mT27NxhV7T68+kgu1bvPabA4aW21b4/IsP17TEHT0KH6GqWE
JW5PfFxH7ExOnKj8BJPhnqi5E+goCnFzgqQrV00nk7DDXK7V7re1yo+SbjIfQFSUmnV+tu8rBGPu
VdXUjb+bIoc/AfKxuEJCi+d4jNfTk5wNGq+rbhaEe6jAyPx6qb84UtmJChSvNE/wUtVaJbN5Sf0X
kI7o4ABpxa7l8+aTEvBomfq1y5nBF/pIw6Oo7gbNmUjNMx3kYQexwjs5QzewRBsActpWde7nwoQY
4xn3cIiXB0/CmBrO9cDw5jxj8M8SxcYEFjVdLptm1BMdzms5DBlDJl4V3UZZYRUp7w2Fq8M7Ddzx
w+fTFs/cT47GjpsXCT5UriNIxgLfNjE+yjV6rHNMLsTtcQv5beZAB+n/fha9zG7UPVaAM7IZyVcT
ZEhFehrgGwpes4bk8UlGBzEQfYOS98S8fqFIyjWAWCNoJ1v8gB5bKyiERtmR30R9pGZaeso8pTXx
Fdb5LM/e+9xFvQY6mmFi7z/OVbzSlQCuAM91Tys00ztCebaJvPdttFFLNGUaYNj8HiyLbAN1xRPC
LT7y7bSSVwbsJ3ywbIqwgZ6gjOBGUair6FPscZKjWYdnT5uGgYbxwBDy9g3vUNc1SSuwIyAy7/NT
GoQDCndB3ruZ9SyH1HLD97NFckA1S0oW0r/TwgdaT2C6rU4NMtthpEoCIWyIkrgT7Qvh0kkPEtww
4EqxAV2pnuJHqwJnhf/VlioEU/IM9SMCu1L4pXOwZgfl37FOAN1bWEUTCtjaAcqQACjUuvRChIba
W1dXBykoe+fiEBthtczIWfPYO/PYyZTp8RLJdz2o9cSROVkiSX9O70fzPi73usZWFCR7JuIk4oO1
YOYjaqM6DQSY42hTrFujICeZSjHC0qgB9TRsNH+uuwJXMGFxSxT3HOqFtdGXiyecHr9pQX5o0uTz
mzBVgSKklsmjmPakwew+/BFk/xLO0wvgINDHdA+Z+Kaajy9vnpIWGQNXbhKCFVaWNS1zLR+QtSBk
nWEKk76EarWTuEiSeFhJaA3jZpsaynEL5xHiqNm2o784ct4zuWzqjDunOH1+xUo2DIIDXXl5PJsm
sqSOSrzlikKGyohnkf2eSkufnV2mtwLM3miHUbDYiyjtjOttXOw/+ZN7SR8HB53lLhjWmKAF5UIY
wWGhYMoNZhaVNbrmLAnnnucytuhNB4OqnUzvGfOemT3GB+ub1LIjojAI8ylzT4SUkyiW4xdpSstt
cprJQWCdH9cOthYxjNht03p/6Ia9esStZfybRJbvWVObX97Qf884U7nhs++nyF7sJ95h04nZEGsH
CRrobkfyHHSOVIKSgmWInuRE36awHGw0p+hr3TNN42fJg9L+cynPzmeiE336CR4FBR2oDX9h/OAU
tpxULrn43ocLXYiweFArGlmfrm6FRXrTVF11pj7A1B5OSb8lRZdqTfPHriSmMevrIlSmuvgZrDS2
FpqYlRq/Gk/uTWrnNICgTNHyUWWthJCloSEbDTz+MEFeLb1KbzPJBDTWGjSTorZkIU4oLLZuY3C6
GeIVQWJOR6A2iOBnWmjEoBrbAnmMBFJ87LOMO3p9JhvFWkYTWGikQXqmtVfve2J64aaKY+wJdQic
4o8sRguAICa2xfMUIqTWxboB3cabyY/g6AjBvnptDJ/0RY6X5etmy9BrVstagRRGF6p7VGJBc1si
bTdvaJq8T4FfN7adUiZH3G7cg44WC8ZzDpscSmZlZsdk4oBZw5fAMAMIfsheg7bt20dAKPuQlYU2
/QwAI6GHqcR0Vu3Kv/WSb6CZ1G/VxdnYBPUNthVg+nQu4ubgGuCguWEUgRUOzDJyA43zN5+VWICf
3dDtCRcEmM8C0+ViY+R2ela8IsuX2ZENZz1jKfxYeZlCmOe1BRytox3sUbm3BS7NmuqdZdPPkC0V
0zB2BPJaF5dcKKV0wryPDue2h7JkZQqBT899hRu6rGQI9EoELG+BSwni7qEYzrljN/Q/SE+lMZnd
VelJIEBnBI6xE7O2JlgmHbSoU1Y89LkZSuU7EjVz9iFBVyrFksJLszHBAeWbTBnSybn7gBC6m80+
depuryXUwM094RI0vyX7idKbFMaLmGJ6YPxsphKdoAWfpdmKD5IMxUWEjQm5DwFBs5FvT/MCueMc
f+syg8sot6WHrtrY2aufgaHLUnPLbkNFpcf4DeMCC0XymLJfmpSV+hh5mZ9koizopGZzot7o0nkI
RsTivyXb3khWFYXAdktINMmjsjHCLkztQlKysAEQD4cNZr5RaTTrBJ2g9MNIYHlSuTNyNxgO+C2k
DN9cWSnNlaTQPplS/L6QL/icIURv6/AASJK3jJHJboIpXIjqUo5uHBX+J0Sxwn2HUUgtG1+tJqsA
BE6rscO1vT4sZzI4jU6qklEXMuA+mD9Vj2JuhfBvgMHG2n+ZzL551h8V8Fujhth6m8xi3vnlTrP+
8PGdkLEsaJruhk6lOLwuNhDgErFQMSs5tgb8RtYpxUR0gSujyrRnlhXU0lMKKy9RAIcWxEFKMS0v
zQNbTpSq3BHmj6MCsAtjyolbSM+2jSY54AXF7IxDnuTtHzfaEU0kY2ReUVxn0h8dvDzoy1NetrPJ
/OSRsVGqJIAk00EG+2AVyhqNwwKmatGEQgDpLVGj4mPcVM0wvDI9o2Xaa8spSAUw7vFSkuazpkj8
Q3moQxVUH2AtrvumnYtXgVzVBzh6fzS2uMFmaEAfCjpSma3EXisHl3qfCe3qwx5UuIEbz6arpdBm
wzpZGKfJyXJuMnb9y0BWIIgaaIGXwPll1Wr4Oyr2IhIhm/89aSTFNwyCiaG66C5vLEq+UXTw1zrn
8NyM05fLgCWZ2OuPyNm/ftVl9Uj69l2a1ppZ1/y+zz42OpYi0fxhe6BDDyjBiZJLaXzmqaPCUvgO
dNpOltLg6TIDs8nbRztz7qNKQhkUCzfa+bfEZTPdwPiuKPFStM+xewJBqgrzbCysCBZhAPAdpeyU
5hgwNPuvo8S09O88qzQjsG4u+EjbzcmSD9q00kjgE0ap7KulVV4Je5FLRrguIcXNWlaXk416iRCm
rThpR+GZsY9wXMGGyV2DeP0yn0X4Rr1zInewwdSbKtLezqSGKTGAKSBEFnr33ck6h4H1+lo/XMA7
/210dNUutwWDg/+54Vp9xFK9FcnMflUw1vfwjKfbesR385NUzYtpt9v1TWZgZMgA7v04i+QcRQ7K
feLPzWBRUGQgyaaswLxQ22jVQI2oKnRIKxOjbWvFk49Hd5+2OzdY+t5WW9dCL6fBf0vp5ojW2LKa
1g7heJyfpogB6JSsXxGcOSX2epeYWp0h/Gv0hXAALLrOQ9GI2AecPiuWtzH9b6wLybTIl1EImxYz
nym6XZnNrZjWqNc2O03d45pwxILTFelORX2ywL60RcbKpb00Zyh4+nXPUfBftdYzeDxEbwUDaP3T
HF3tVskC5EA98qQazp50j0y9xq8a4ESn4GBGpn4syfKwEsEcLBfbUfrBhlDVY1E+/ttdaJSZqPMq
yBBTjE0X7iKbm9QUneLyw7/Yd+YFTb7DSpZAHdOtYDQUEufTrlFrYhwoSCv6rod5S0eQESv/PzoE
TZ9aNX9eZKySPlXfaS+1gyTkwHRH5LO+yas3ZiqBpzHXKdFDNiIg+Tivzc/1XVbRSSPDa7ugxXjP
Aj7RAFJz7/CRtb2FTgJap3zd3f2C6QCaiFKE2eRD9GNgx4w+yrvt39Mj1VE3aW74ObKMaeeK0jam
FF9J+qpr26O2FXEhIuMF2yP67xs62KARv1Mk1R02aaCF2z0Gkid7aNICefiPgJdP0PDy/hzTEz5C
0wJLCJ+tMovbELkHjirdZDqALbJe+OV6jEkL+e8ishV6MchffBc2Eyktc4qPeOAzCd4kuUzbGPNH
g5GDDV3e57dKES39jZ6hnCFhtPMzGczDxOBP5Y6Z1ZOnQjPzrWSdC+q3YkZyVX+zrnxrluMdBmfP
lr/O2N1MtFmNMBZlPJaVrlIOiLFiJ87o8XpW12pVAwZjibH/x+u447LjxEQB1FRTWWWKBa5pB4AA
op9JwpZk+6XeXqc0DyHSw1RP9l+BJjNuZYXZGYHthjpvVXOOFuGpajePiJjgONDzeoBiG+8w1IMu
XoeEPnktRfqoXd/nCFB8rLE6rH015JKtA5uIvIsZ0uzCXEdM7Fe4/zafyrbQ7VSFw1xFNDiZOeUE
+aVeIEjRUa4/DgVQGZM0/YWkAbP20K0cvs5UkowCkAtR3lS8KCj74SYN3PQhgVY1HexMrTobzJJH
kpCHZV2rOIl3w9oL4MeFZ+9Mp5zyX3P+mBLftT8xqx99vGiaaaxh2lkYXuM6rQ0pFqckJFeAer5p
7675Gd09+8x+n/aeGNftSdfbaF/n8u07gK/9s0Fk3yLDcU61wEEL877IqV7ts22RTacSbm7oT5yt
tZwQ9e2J3giBRhhAQOG07JtrueT5mCg6aBb/fqBnbLGBePu33xyMxMlTNpUj183AoB+0tYyYiaiL
EOguuACfVuT8qEYnOGUc2tveh3A6hSeygTPhdV2gw3fTOSBMKYFmI9JqI5WSzGhVrhzzpnr1L+eA
0F1oc25RUtO8luywzM0qc4H4lPJAs3uPZkiKyv37+H+v4SLFSYUnVsyGBTOCnJD4weVycDE0lYT3
oiiEBJwZdPHR2ZVdU6UqjiEV/l0O+iosdykVqcpzKsjwJ027iBN8Os/Yq93dwgco6x2GGVaXZR8r
+Q6ZSOOelpTxx2oMg+i8jXsoaqer5Fs0nY0COPb8smFd5X+GzSZ0wuPJuloazX97v8pg+tPX4L8a
YyaA3a9U1wcXehpMH60h/S1Axr4/wRv65VoAmulLLrjkIcHAeWG2TfNDksHU2hh/ydzL4P2xNlzd
WTP3RvuTo+JJ3gXRSXhjW9u/utTPib0XvwqQ/jstWcplKcEopCoG7y0drHmlbC8OpPFW51BzPHx4
Cp19m52Wz13hKJn/QwuTqs1OEBvAlPiAv2yinrN4xlz1D7UEmh9fTndxR1aQhiuc0mHEFZs/Mcsg
CqRMmzo/RqiDtDWpZVIu/lTCThe/eHkouoLw2nzLVV2c7Z1Cp3ctrt10FCWniZfsGC/WrM2zTEwG
WiNbsEkpZXuo2+nCr1VpXHZ/Kz/rcasktwN2jJO7ecsE4QGWRWzxwxU2QVTb6Epuov5Wl5T7xYws
NW7gICc7Bsb7V0UFfsBuX1a+sgv1p7wUOBtuB7IqzAk56xPNjPBbnG2HFeIUzbVd7K9eiT7su52H
JcRycXvB6lVM33V6qF0oPB6oYgczD11zWTpzTsJywor3hNPqpE+asWG1tWulVNzuxf3Vsz5tFYXV
xb2dhai4VFNWAVIqFWNpQk/SrjH9qk+O1JiZiEvYQnDrCb9DQPM9u6YXV+X9y8TnA5uXknEGPPm/
wHA0IsLAqunvp7aQ56ue1Ztq+5xN3XhIRKy0DZgUcrDz/rrTkqft3FGn2qzRaCNOhSZHTUag6sd6
EGRYJ15VvNMaVCH1PhszodBr16S8sYpZTQ1z0nmPBlvaKsy4zwb8YjMvGC9bcdsjbJiIaUNA5LKi
ALWqhQlL2WFNBiFREO5PHFa7ZoLsmFycYuHX/7rafaQWLk9PsPVzqCctoKlv5zGxfm2YXK04VJZj
jhalk0swdZ0LJU1r44ZpBPehepgw748mh0A15jxObVIJv2PoDcWfYWLIqGPzLWmWT5AUZ9Qi4HsZ
IFbqlnxjt1l27CcGq72JoC+G7PZ5xbW55cgfQqc7qQo4oDXjmL2jwqYhHZzLjIbFkZ2+ucyZtuG6
e3PaZm1n8k9/H2s+cSYV6JuPSfEWkuuUoswNSw78KS7q75W0IuX1fgILlq7z1lXM8LszqALeni3y
MxszOGQca8gwdSn4LVbhHSL22MWAhbUy1dcxGL/XLVMjVu9+fmILdcTfNv3sydhKrvzYnRXIiFke
nxuKPNutCzWzd42UXPx/Y7cS3NAO85lHjgWKSsBkum8tDx7D62r3DZJJIGvOzX2pVxVZ6mM0JOb+
Z0cZjQq51U0dnITfv7D524nkZa7vXKZ8Jxpv6+wncsnXeXI3s4oj2oW21FXPTWmCUb39CUGmctFE
QopnFnQMpEUtAdMJIyKKG7ByLuRugSAWej/J/y1AxIomf+bnKGn9WKMBLr7ExThGt+MRd712t0v0
lvOyEaal9PI8YXG5me9KGGDipK0ZB7gnnqYlQH+dfsaT59bN4X44QWSe53cfdGKZ49f+vNvYSgqU
OxHnvKAzpIhjB1Nk/q+UE08oFLRxuvk393cjNmIpYrWDYUQz475MqDdDeqF85gpP7ZfX3JBkBeJC
n2mNFlqZaktIoDUgSeRxcPfMPZWETt00FLiOMzHItAuI7UYCVhpjXKUq2og3+/7J+cobPuVs4pZ0
ygU1SHQJqCyrNcAi4eQRd7BaPwivRe/Ym5ioqbtYJYf4lRL/07NL9N8MupiWr8WPwMdsAKb9+Ngb
Zk5tbAZ5a9R1gMIYF/7uE5kgUiG3mc+7Qf814W1AwaMVRVXgFpo7fVJcV4gxGG8JfvRcuE5cWHsk
RcehE/BZAJCKWmI43sINOWIoQbxpn9zZ+wmSguMmq1GKwJXVZlyyubP5gipc15tAzKowwPBgEcs3
/jX0XEjeThzHT0h/VNRcnnxQnWTd8VRoT95di6fX5628OzmcU85me3229sxlGRVED16SuTG1ywoO
dR9YY4yfZEpzxGxZwXUJwPZUlgLODXEJOKMud/QnatOfBBU6KWimmuCwkfacwVhLxQppKecZhT/t
y01VtcHyW/ZnHMmmkGVAUU3SOdqD1lPpWYvHm8A53v2QY+lzUjJBj8Idq5D8AjnAp1zkrulFgwdx
M7i8Qn1NwdbWYazE7CuhZyjxWTyanBNd6qJkFJ3k9NoFWuo2EaEDeT3Ji7O9Zx98kKVjgWRJY96v
FYueUj4UvWO293epbTcuQ8+03UaHxI3wbCfKYc60YeHbTRmMwnHE6NSPrPv4tTxfJfzq4UryuVvj
Wh52IMvmrNRrb3FVYEBFojXhjQGQ1v8/7CuajQQ4NLurAIsVA+msNqI+cE2iwOpbcV7xIQrbPAGy
HUxXUMr4BE0e1b+gBy1tuHP/34TYMVbuzfxKoe6oBiX/nZLhfN+Y9+VOTfC21A2UXBcaBfevT/f8
0cmK+xLa2ti7QIAtSy8ebqQV7Uh7t6QDTYam0VgoJcWelK+a7kdoZ1frTkbgVb7rA1jW9SqLonur
y/9hCzgZf5abFAIDrsn6cEMTdKIm3Rv2lemHim3/IrJMhEKrl9vU2FipnW7X7hr3aCcLvff/j8WU
AavRb4rsX52xrVW8C0QlyMGk23NBbD0raFHHgA9rHNQoEyso1ivq7cMz/1Zj4neJvETPAFeOSGU8
hYoipaJH3fmFqh4KIKOZXt86ZGOlhh/OxGl4HJUUcewe/0CY8aPrOlOTeQc6cvBQVQ+TnSdXCF4+
mvO4J6cQNx/b0IUBQ/gntUIKXjsvFZWDOLynOxYPAxv3MeRFOAI9Z7FXA2PweiCvsf5tr/ZMzDhq
kXSaSKLQw5Q8qUZS7LHILfDbQwAcafeqdxiFJy6xacY/60R3AOTgBT2ubk3fjOk3DFJy3YuHIaq1
bqiEatJT+DIKa2MZFJhD0wsNpwYRjrLpyahPrYTNKjz/noi8Ts11hPtF9J2elMoejGrRXu4Zlgyh
WfSybaKh+T6wyICbDpUO0ZyKJd7JqbLp1qC2mI1AhtjZs+sIToRS0loN2A8pUbCFB7GYxQ3vdSzo
rxKlzvdTV8N4rLQ/0Viq90wTD1VckV67dbiyqvLd5f39zQZkYmvoD4eYEWY6Px5/4Tb7YcZ6pLPS
PB74e8gufjXQVLw2zTaJcUm7uhBW1BlGk4V9Kw0O3OO2qze1lklay2YoPI6iG2sHmqrLEB3X+uOl
O6YsV04/6tdmyYsTEbsWYSyafXw/XzL31fwnp5GcGg00y0qV3Z5wfhCcN7f/U4xY2asyTgReB8iG
z3NZjDaj0TMPri6kifZ8CwTqhV7qeHp19G8C7XbJajOdvxBGUAg3ce1lzfKhfOxFfYzqYRi3U0dl
xXomqbox0aC4U5iHkIyNNq7+XttqkSSrP0SDIMnAy5PBk3+PTEf0u/5nWn1kay+DtyhMReAeRZUB
VfhAFcHG4HpyJsDgwjmj8IRlM2igoH0iPiO0Mmz6uipXr7eukt/0YUYTVBQW3nE6lBt7T/XSFGIB
FkVtRRPfBq3gGOzKHuQbCqgHpCepLq61ppyIkH8L5dwPAuvJFfjIpdwNK0WOF/nrcVyle40AqKL9
xUiCq0aOp8aogHYQxExKfeSualT3gw+P5neHaXZVva3+grzgp14Uftzi/21ouZZ4Ztb4ym+sxyuh
gDbpW1BuOeB8QEfgGSFfr4NFxQqhLx3NiwqjMIEJZdKEg8bWXZmix4v0zYFNkn09xpkBpSKWRTuJ
jW3OcRdUzwqQL12pTxwJxza7hR1icXlUBiHTFd1Do2d9rPEPAuL60fWd/fRT+DpynZ9QRKEHCtjE
uKp957n+svCX1bKgZzcSKzrxdALYfbRd2NRGLktmlpB1D8V19fw4QNybd94h4LkbuKY5N0d70J/M
Zw2P61JIylkpBI11O/XlrK2p0pw6TjlljHe/63Bk2qdmEuSaoGBZD5VJ/WQuR2DldJX1R4xzIP8U
i44KAXdhsuT7GLL9Cbn2JHivYz36nvW/X6qsgZe90bn8qjXeYX+0GcJ34O5wiw/UiNV3crFt5mLh
NBNmBIelX04dAmNe1AeCx+A/9NYG5qaApEK5f8qIArGSpxV+9sYS16oodBGAULNPxNjpFqbnd0nT
+Dt+AiognrgSfuZ0WP84LaS5hpf9HJ9mirLyLj1a08CaEDpUHOCAgqyaDV/yfjBuBZjt+0UPlEmR
TLa1gG6xgWuaJ7NFtCdFywHKI2FUDNc8QiHmkgOiYoHvhpoEDaDuYjo3NBSa6fn7MYt1Rr7kHuaj
D0253tKk7gyBJ3feSDKpNz/95iJRi4yn7ERi5EwaqHAS8jkYRKm3CkfvyNZsbgMDfafFA2jZluHl
gvh5ffigFP90KQstx6WBp3PztO12/MTEk1CnofUDHEah8O5B9bK5y5x8BJyOFlG23Kpf71aP0n/f
ip4Gc8Bnc250NllvBx2Vo7c5cXkdyI0FABNtRhVNssphZe+11aGgj2Y1f+BTbLGVYfOyAju4Yq7Y
KAlyR7tfGOBSe7/HXq3ujzsPB6mj0vSjLxh80fXuOn5YoJ5oY0RrczLJWcwTjINXO3cqOr5estu7
PHP3yKkBjwSGbiIfGk3nS95+7FItqHmYNsdZNBXI5/5IT1Ot9tpL8ilLqgAj0SjRq/W9ovBJwni/
UYoBHoFwLEHqbfZiEtvCX1wWQdgnC90/jVQIAGmGACwq+LcStilSdqyaiGLC5Nhzax8dGqXHuCdw
5+DYGorqnqhL33bqtX4/AYXsiEx8lfW2FEr6YJrLz7zNsiMYe2PHfLJZdr1qVJ0TMdhlzWe+82ml
Bd8BAdlVs4gtyoJi5p4ksRCsNBIj4HW4sese/FWI539JnHcnfQxPdbDly/QW4UMimZnRLh3fc0WZ
U45KOJ121XvQnBJTHH1oe/eUb08M77hUnWi1x7FcHV2WBCsac4gvsBFR7Y3ErriR4zQfp0IPOJzh
8R9vvezgUXtDamYsrs6MtdjFp6qvq6YHO6A8aqg9DCz/z+MDpLHmjpWfGvJxNvC6U4a+D3jw47VZ
nVQAlfG+4Bnneg5LqTEbz6onvv/JIj/abXeo3FigeExrojn4dAeABPM4Z4NkhC55lSIzPKSN0Hss
oeXsNMCOmeYz2iAB5bDuK1AYCmjSKuAMYGsrpdIptHFb8sXDV2ucbW1WAmIjWWigaESqqmO9TWUr
yxJivQmRTULxrQo20bPw/lZB/QtBRmRiL9U3VObhasui9AlTuGwGwoy0iV/i3HRO0Mt7qym5ylWL
bzIuRsKMmsguJgQZWPTtd9TvhN4kiCq5q/+QzEjUGsNO60PdSLR5wnOzpVhxSlwZAdqIQQhamH6/
1ekyMuOqSHEDBdTG5XokGv/dx8s9LocT7sFFsJfPljx0fpdNx7heQ+Jtz6ErA0k+6cehtZnkxImL
cAf0t1lm+sHMaeSU5hMYsY9zXVVJIj8qa4j3IWtA9q7M44dZYoQkAmM/FND8U3Qx2ns+P+/zqhVr
7K6mi9tzoDqcvRajQPgtEHEQW2d5mECTk1TdTuDLTb6z75nKRZP+I+BrTB8jqBsz2G7QmB4w9wNe
GftooWjebryue73xoZqAK4Qrql/4hI7dZJXohtLljKNGgeYjMtbMuajCfPay2C+jixi97HLkfgZ4
OblVgtpcM8CYZNw47/fEe+rhaQiSiD3uEWnk9XF5/Y9aCL/oirn+YGXWQdtW9FGvf8trrJFS0EhZ
RVogOlGwCzxoh8HDaKGHbXp0wU/2wHec5AGG0tKF21gOMUu2kt11Tx+avuIvhyo6zim735Z1PG5e
FYGGOwlvdIprjKy3PD4L/P2UCBViqSONWe8eyglfVIArVRp62q8yju7elTCxdKKVjImFPGN+CAq7
RVfdcklv4sBWY0y0Qt9nMq64Tl5+A3yJ1wu8WUnzgw4aC9eULWlpTGX0IN26Px8rFkoYSBTanKBn
yDfI5fKbdiRcEeg3OpQpPufIusgSSgW3HpdF9FltfV1nLmGKzi5qtwPuLtIlQskUt1coIS/XQaie
6/84c4iWCgkLqKiHkeZqxpA7d6L3S3IZx9tmh+bjGWovy+AB8EVcAVYRhhDVaIwk/MoDq+nft4d7
bJBA/pzqrppGWWYuvvsTgu7sCqD7QaY3G+fMklKEIyeoT5SoQxqIA5X6Z8anrPgphb+zM/daFKVB
GpaUCXJHWOum9urwtIIwGUFMOhcRrTzListOvLKYrTnvlQu+HE15Squ7HyJ5ejFLcm+ymm/H8FYC
O993P6rkgZyNtvYO4acm1Mq0qNyrCIuj+prZuw3X5b4xrluK8BKZKyj7+JW6UpwYPR2VBY+U667P
qd7cETBR0rS3OuBiqjDU1Xfpe8MKM6M0hyKa+d1IiccODlT7313LviiLKmHiiWOUBTHbcuVXV5Lt
/YNUiiI1oL0rPAiSgr9pVz2bNR52JR3GQP09/9H7Ee3i8Zvq1s9I5bfgYd5UqezpluNN5qsM1ftB
T3zzE3XWSFsxkxak26+2W2sinRyeh90xJnQZalfhL2hkmqyqbaGZ1dVTGA1J/N8JuI3ISX1qKr5Y
yC1/YsOsNjfNleUIEw/6y0vGm2p+ld/KjKzDqFHU+efQ3pRzHUgkfgskJlCcMQrFi3KLLSgwKiDD
tcvaZLphxhHq3yKW8gkP88xEBNHfnycRWt0Yrq9m902daHsM38JxyzJntHauaWTQNku7gK+grmsg
XHKn8FQUaBNp9J94Sq2EyAoGB++Us/XMp2qX4KOFJ+SRTH2cQ8N9o+G9cie1GloXhsmm6RY0tBJr
hPiZ5gKVEv9/hpG9mV7Wx5bg5p4UyYT9AEKXHtFd6rpcADluFw94evalC1U6PMIts0GRiaugxxGW
m3QzTm8iX8G1S8FptNTCd1EbERPeufES44lPolzHHwL5pLQAtHa12sWzb44q+//NhXrrucZguEUY
URuPoYKk6NfxGDz8pKFabXHFpMI9QbmWLXR6QTCU9tQLuBL6X1pomp09LOYKb19jcTAwKXKciKHX
g4ktLCggwEyz4neHet49AWel+T8r2V63BJIiuDARIG+/ovCEfhjndEOOqZFXZT1W/pdEkj5DdlcR
KUcFUTlYM87ifTh0uDdNShNMKGACy+8POAgE9e9Gjicm8GvywyeCdOMfQUltuRbUpgRPeWYW6vd2
jp1WI6ASwwrRFnoE5jemkPvX3v3olClTAzUwoC5cRsmzsj1ugxIWAkTKWnHA90tqQgWdA06DKPw2
SMEyVebqfexy8GdOj5sr800ZsSjx5acoQtQnA7pjcPB35TndBq+rhatfP+7D8R/4Ctuysm4SZwAD
IPuOWcfERCmZaIHDBQ5NZWQl5hNyg7kr/v1L5hnjCs4Eb2xhLY7eqZ1de/gDOkkHM2QiHnGPm82n
OLpFm3Ikdx3U3wdKhLF8+AxEj1AcE4p65OkmcRtOzTVJNnxf79+05MktP5Ezy5I0YuK6594xhSDp
jeKtyMEXulYK/78St6yyRgOsAfqlTfNWfLxq/uPYv92qxmhU1vicvlty/7TmoIRN/2tb/sFyCx/G
6GTjR0TTusdvnR05zZsycLBHacdLHC7WJZNqAKnzT4KOvyiNtgESPU5jEb3niPeSLtdBFSsOvals
uaUn7bMqO7sYTjasMw/1+/SAwZA0aCbQAlSTAPxOd4ez2wySZBguwen0iy8GZbcfKTsxMS/gKcUi
cw/cGTKL7hs25sp6oEovyui8cGTFxtVucPrNKesD5WIa8laavAZXy4ikxmn5H4ZQur+CjQ0ggav/
e8SiSBrIC5Js55i7W87NQWAbQYHZrKhAtRzZL4VIY4xaWNQHxhOfOHba6mIvvpX97vh715YszNuW
oi0zDo8Yt43pR9ViM97vWgYK6lTwYgUM8Tjsiuf6GVCGcnUFdWNpXCgvQrxFmiqlCyPdIcHMDP1M
nNblwex2WxoI5XEEwSJQN+/Ctsw/Xci0WBgbABo/qOQr/S9O6BkakWUQ4dKmDICNrqXw6WMUB+Sd
oMNox5Ch75vqDfkCMcswcgS6FQ4LTW/kSZgqLBM9xpVEefb0potpKgWnapO2Mdw3Akt2TFq6Cn0c
yhuIFIZ9vJK0FXi4m/9/JIRr6+PqeAVovEoAaHBD8Yvme5r5DVjaEKKviFL82bAwq+fMOY76Wo2j
0fMwfTYGIDAOgVJMewZ7QX98oh6VUcRzfL9R3p5QV5LBn1bjR+0ZDRKuIF/dfYnXk+bEKVUYu8Vw
O/vuW1xUVp8JA6MuxyP/GuCmFGVnH9D54DzMedFMwf3qHstCu8WFPsXXUCsf+OMwECEFc0hyfFQ6
N36z5hw3B71sVanhND2VXCwZgh5pUlkKhb33ZzZYvFnOMGMarokRyM3pK8xsgbEJ0B18Q3ru+c9c
F+vJA9T7Cqr93py6P2ZxXuo7d/KE2xt+zZv6ixBJck0YnEnlTdHd9dPC3UmdV0GJ3CWNUFrpw5pd
uw1sYE+Xu5/Tx1fe89zIg+rH08kG2YjW9tvEJebUEy4ZlL/7KFZe8KrEmAV4wwh7FTWjDjZPUwpY
bHd71AD+1jPaZcQHO3LmM6wDkt4NDB//rasklJO8No8vVUp3kQ8Jha7oZuweS8QkJhsErFl8L2dV
ysHWle/Y9ZIZqlrYlGMqeMbt+6Z/x6FG8Hv96b3RGD2bQTimX+rhHo37IltaAkL4gGc+JEDkQwPO
Nwndou1HUKUv+uFU/uTFkkBOkY7BdvhZeOO0HO1n6hNk9Qf8MiBqVx+GbdAJpem+TtvFGB7pAdrN
xZ8LzuUSCUtROfnK6gMIb0ogM/sxxQoy9qcLwEZKAC5zCZyz+RqjogsAvZMMqenXC8+WWejN4vBg
KimGCOe4/0tVtB8AMgFWAC46w/fMYRCyZQ712/tsvour9Hbb6CDm7/mZ/6W6srsM9sFLrlYacfoA
w5o9ZnrwtS4Ou3BWf7V38BPS2dFGV+PmN6K1en+9oQCg2jPKE4WHg4OURad8JxmC4nJSL0PtHImh
MnVFEhZprk0ht9vaYD4jzcIUA/yEYiLeeYj4O80CVyqTsLnxx9dw/Rz0Ki5VyYge2PuOjMhYfZvK
BlQf+oFLfr4M7W+2i/GMNMHCPYar/1QWNtURabkmnzDhXQlQCZp54sdk+aYSlXFEIiduBXSgcYTs
ksELjc1KBE1/Ln1iRxyJ6njsRKAFPmBxkSCNFJYbFmJNOnDAI2XwcPOtwKLVskXgSLivH+09E2o9
vBICMVhTHzTRM5h+O756YMI9fF28fju9ZgmaQaVg0dXx6l+hFcYxgCdSdhf1yzlmmIGHuF8Jg6QX
ltSCds1iVasZoCSNp1AUkP1L/L0v72mpyMhzMkwq4aAJjPe91MTdjOs9xZr0zGVGZZuL9v2/s9ei
B+4WjAs6WcKyxm6YKA+j7Hmk6+/yThY92ESgtiIzZOJjGW6e+8puhzPe8Al3OsYtErZ4sKar0swh
7ZG+96ObwjeFNtFgjR4nXVnA1KXOyy+tq2iok39EQQnK9fRqjrIktkMjwyi2XMcOTzpGEkI0p3zy
HQYHd0NgObJitGsjJbCcrqU6QC6r6tgeKM3hDgzfV4LvsR9Jbr2t3b1UovpTu+pK4inSq6qCkl8j
CdrfUBgLH91H7sVZFqrR6tmh3vIH3ReR7oUH3zq37Kf90Ir3Osg+b2NKJyMVow6GFcX6+W11qG7w
4KDW+3texOUuu9XjKRQC6+qWbxgcQyN5BD58magW7phiDvTxDhw6DA6tbl0PA2JAj+H+NA0esz9w
RTTqbTE83IZaD/e03Mu/3534B4IpmX/rrCv4d4ZqoNfujyf9rupO4e1/t7hHAJOGeoRfxse3tpH7
WeOr/WaFatipHmT/X4l1nUOpmOj6C5+0FBy0w+ufy2DgSuMbUUOidCnMOyRE9koc43BAK10GVWnh
+WngxC52YDbGcaPg8VhCxb9DBd3OfW9+MbNQfJ/TFCq5iI+Hys3e6PLWe2MOJnyW4CMwgzVvNbv2
GomB93FiyKFX/ffNI9smr4EQbYY7s2B6O1BuYduXKRKbJ5mjwFMvwYtdoO0ZgQ2a7mgoqNp1bhUz
V/nja1LTb6I3n096iv0fTpwSeAdxBDZXtUsEnCPX0Al2CAlCmZp6AlJ1b01rZ2d4BCssO+KYKPQa
jgS5OOrjDSUOkRPw2hksya1PbyZEI1TH8hT6wDuXfFGjomhW/RE878Am5f6GzasFv5QLXQPszV8x
EE6xhO+pKoDOI/JKyA/cQaRRyD88XX5vY4JmlSjrFeqgCu2H4AFyfGSj+9nsSnwIjnjXmptePbK1
R3HHVTRmIApNXb3zmtx8oGiCyXtGX8dAvzHgYKJdXkNsD/0QdrFldwP/7S33Loai4/tFSBN8xAk3
nfhDVw/1ZD8ZyVT+YfdCJtAaaUQMr0e5xlVTkHZz3WelCbc+IK9UmIypNwAnDTvW9vZUeqQ8aLXv
fJdxDL20w79IX3DTKs++2UAfl+qNGu5/j1kx2qDtcoAYPjcah+cwKHOqxaed9QajyPqBX8ONn3+2
jp8a+Kbki75AP5iyrs42z1w+VJsYZk7+m0BObhRQoXsQYzw3cCvR2rKe120RfN7zuqUDNJBaKPlD
VYd4CDAjujQ8SM6KLPbKuNczdXdoGRB+lNr7/4dvr4hrPfb2YWT4ue0fL8pNYgYEhRE8eSrzzJeU
tExja7a0L8feYoKa1yTrFtSHXaUhp1ohKMfp3vGgCzjLLFCx7Ixj209/SUUc9dlG67S/QaIwGOWy
e8iGWlR8+4szR+gp957oZRxDxjqrkIuqimjfeo/jSTgXrWEs+0StuE5WZDALX/6bPlttfymKL8Ky
FMD3hI44s9TiJxcvO9IDRdTGwZNsz8AJVBrijS71fWOiBwcolX1l/U9yIMe8if4VY9SGDBd9FUAv
rLCfJfQbQ+RhtCpwQdAKeqNEkW/DNEIFVK1H2Zzvkq7dyn8K0liq5wraTm87YAk9oJQcdcHicKmM
gkTJfotCvVG6aYpNnFWrh3IH9aweBxOFzbpbM8dgW+7h0UK3PF0sLRTSleyMUCOyNPX5+MWWBgAo
p/BSczfWJV5zsqeC3dtwMN86ggtpppJFan1iME0jKsMYlqjHfG4d6+0IN3/kKFYRL50U6HTJUq0w
YMshCfgHLBiIvOiozcq8YfKyUih/ACKvIhShu0MvcGb3QXSt6vRBWJPZ9WmTeY3URe30JdzxHDwx
hX26wAdSCVlMXiT6eA7TAWZuFqZ6IcFW5SNioXhTkr9qMJ1el69OJxyYa8VXlpb+Twxvni9GyVFr
Imrq8/B8jSF72+AaqFu2Vun21NbnvpnGu+IaSUb9A+PpvEY0arony9AuSN4a11wC3XncMP/kiKHZ
VSruEZRmVb7pfrnr5WW8EjaMY1DgLdmFeFwuCqRXgaafobEGCU7sS01iZku1OrSwncxW7FlKPXLi
ZpheDoo3lvGdKfZOT8o5tWQGQLb+FXMr8z64ChTu4daSxU4+CvP+jK53Gx/sRryVPthAWvPrJARj
ZizOoLeFU7QW/8CV6y9ZOg1cBGH5IDj1GIgs7dRwYJRddgBZ3H5BQ/SD15X8Vo7+9RhYHGhCU6Yb
tMMhYexcByh+dmf6ksmxoiyvzYii92OkAQ5OzJsCK+gcQ7G8h+T9RdX77wo5BIRWaoSaRj4AJhxT
k7pofdLPiHnPd+LskxixFuNu5MJtphDcALeKvxi00q66feTIxvX3V/1bf4ZfmIHw3P9oOWnphZTm
fYa5JOANfXC6Msi4leQLLalUx+p9R2RFl5ZsDw8BSE8ynvbleZEWAAJLZlm/SG8dRWbzBtoOuiV5
794pj/w/DcLkk+I9rMHEygcMgZuWWXrIbUhB6/AvyB+FhwnuBWOrdbwmGNbwFEJchqL71VnTW0r5
NXnaUOyH0ZTY/WA7zLk4T6mt0kiXHmhePY7V5udWVR6hr0E073xcex8rCDsZ5f2Kuk180vXwfwQZ
GMlCEVTjZBo0B/2Sf0bZx6szmPJKJHckQRTjoTk6b3vY++bPawirduN0F8Qmzyjmu1G+ciVzhZBb
RmbC2Ki4kwGe5/XDIfgtAz1HInrKrh9HPo4pOl9yWoIO/nyQYSHEnG85h6sBpYy3ndUbzv9NAXyz
iT/mg+hiZ6hPFff1h8iNX4uFXMjYZGBkYCSRX200k1pv9pZ1SzKeuWHSIUIt6+YG0blImeQBPg5m
NDdGXRFHHL4fdN9+pqQdKydzP/xlNLj3NflOQ7ZKEB556F0fXi/jmL1H5Aeh2mjrce+EMxrqjqIy
MVbJRQdP03Ph0xa6rvD2uLM/wTh+pWNredLD5JssQLNmFQPEoHpHFhqVXJTvmgsdCKuq9fVLjY7V
3mnyrmTQdgjDZ+ledy9QASQmdewMYSDU+zC8v8TnXF0sE57zRtvX1Kxa5Nd98QXnguEvTaDGIoPK
akOebwdMOdIa8O9T+yKBoGSmFpvDT8wuK65QvnIy7TeVRsrne9LEKUef2asPX1iRnhjX7qsdb+qz
lJpoKcOz+ZhE8vOZ7pnto/PCsdmOenMpzAb4xWPYD81i2mfxFPZE9rZKNGYf7LOCgRITIjV2ONTU
ETut5R/Y/DTprOOn4AJconfI4sVWlTJCOyZcqASDI0leMSAnu+0jVGSPgNZ0r1ZWdY5kSPpM+ZHv
pSYSjWKy3rW1bAwOcn/JT4ImyFi8SCu7RlVHgul26VYAq95C0kYQP2eBNd2xY4LM0K+SmrQEUe72
FZsMioJiiBCFwUnNjb5yNxKs9VYClCdVLFOfUKI3DyXnn9IHxS8BCRdyK/fZ+b4YKDBa9EWEsz8h
IzbsD+vJ+09EFDRrCNtw37H28/Y5tLQWaWU3rbgHEUSyVSVYwtGqJVzuDiZweGFmtAnM7JOeImRd
ktat8OxvOi33NLLB6iw01hq1oyp6yhJj6V+xHm6L5EaHDJobruKX5XLao5UZLG8fm3ZylrUN/ixU
Sav224zajZMkemztdPIZcPu0RxaURcAjwEs8q1FDzDqLS56H8vT1sp/X/ZktL0j96B3BH1aNpE4J
ErbcPk4xDIQY/Y2D/VBvuT65hVbvgETr6QqLuaFmOZCNZfcXS0R/9QLTzzicO+g6D1BeF61b3ipC
f5LObwPlbWTPd2g/uvaa7Iq5/InM3dEApuBYNm3iB4RQfleOW+HC93uE/2WDUpW2Xo8ICMTFdW1+
M9cA+ngPu/tbAYSEIuoHee56fvOYKQ9FSvInFwOSwRIDgPc7wZX0/pkqmOyV+VsxovDIjCVPWyp1
Pu3piy0J9KKlFpV0An/sotzdKLsGmqm+MSKKT9KLqkJuyr/okXF3+YU1Usb6JIi8rMzDIsXhXd7e
Xgc9bCWeRt7CE+kc60kk29MTIt1qLozFzRcgvJxkUjdoeWzgNz9SuB1wil5JHa2789+tkZmF/zZI
/aAbpaTrsyi4J+jZvkZrBAinBex5M9L3eJL01RsuACh/FjLNyrnuUjKhRaD1U32H/A0nPONcxesp
zBL/VbynUUUJ4qfzCqVp5uV0SFMrwHaC7p8mSdLjTbhvXl8LAIQfyfXeJLgqpfpMNa+puqwF1GCq
d+qbEkSsg+ZzOo7Hrh09yvfSRBuhbl1yoTtRaIJeFB+tUf6ogHvDUmANwhNFTurT46gGmZ7nASwL
tHdAX3/3bboN95tVAjyHEr8a5WeJ97efRCSGyQFjGrnNHGiGml0mWbEn7i0HUw9vtSB7CMSG5kqc
C71t0NGX5Rve7nfnyTuisM1lxQ09WZ6Mds5R9FwbOmfNhUllMQMgt4cWcnW4mcg4p+LN4QEQGpW/
zkwefkcuyAy4vMIPh10K7DODL34ROVRK+ylwws5UG1FwWCjYfbRAUkFXBzb9tT9LeoxvAxVm6iA9
pX+5QE3jHCpoAinMihxXmVRjTTBTynImL5fkAaVKEAcalrIhJ7naQEmq4CkDv1TwpzWi2KKNRXFP
zNojr1V0w8jdTUc+hEpyyln0SIS61YofbUIWo0bB4U313D2yGETWMyshCFcWEODhG1OzbkKQMyxl
kWawofth9DIgLiY/G7dE4m2Lq8V07eGBNif/vFCmN9dXbYT+a4n/tVaIVVG9lIMGQz/JyqeSsHHZ
7jrjuZifhNEY1KCxqSL8QV9hE912XNEWREaiRDtS7NQ0jw/M647DM6roCQUYNRNDQX/1nzN5aQaz
ueZ5wKAOiwCc5QE+qopMcs01AQ8zqhke1/evjEaruBUtK2atP6XxxNT9G8EFdpBoZtvZaNIzIKvq
+0H2CFgCHj1bQO1LRIA/45wrH8sUMn3xEGFUPAZV16Ot78WXh8ALDxjbujWSP83uCSbI0MLBgb+2
kb6CoHk2x6sUKAHJnq87XcjxtoanjBYdZCNuDrh/ftI53ooYed0fC5fGFmIXhNYGNGrzR0CCRhhz
SLixXr1VXCaZC1x5DOEixF/8U/BoWimVX0UEknuStNmAszSd2sjeiMC7gmktBCCaEEPwsCxVZ7g7
CQc8s5PzqA9TTSLxcCuH03b1EB1nsofOg8dCG1MheK4v/B8XXrXDzT9FJ7GhM7Q8+xAmF0MVrrYt
lX5XSWoKzkB/NnWc/YJ/JvlC28NagFdyKBPzmWHfpOlPgaug6djPIkdyzqhSy8XcoVNFgU/Ds/kG
oFMz2r/+FMRo2J7vjX2Qak81TExdGDZOcvwVRb5tA6IrETCm6EX9H6tPAoQgSThCGFWnGy7ETC/3
6n0+PQAFDRguvsGzCJoyagDiDB4esRfIayHN1YGoGjkLQCbkMEnDo9jYuYCBgGxsOxQj0/QP7Sqc
AZwJ0oDDE6dQlXfc88RSmZDV1FDAAd25180Igiwjjogwf+LaWkmHNkkWTxbkLmmBfV4d7WbOPn5+
e+STLpMXEk4VcqgBLU6xIzR2UTQIYx3kJ+CZlN6pwlhZnMO5kYX6AnqIvnBz++xp2TpDxo+dFefW
HpsHne3rTthC5X4ZMNAZ9IX6qbQatL0WVdrmqfYf0ohJGS56CA0rtNKDbhRASMGImmjxPUHydwcC
mXhJ7kEzUIUu3yI1nqd+V56Yl/Aim7S6gXMY0cogBclq1SQOGlYeXdKlZ3MfIy8ALsG444FNV+yR
G3XQQnm2H8L3pi0wPsQIqUjD1YufKml5VmzdwMVz4LSDdca47n+E+KDFXhmeTezHFY2UIWbpbMk5
YqqMEP5Oj5lbAgbjQTNHQFH07bWLLM+zotIKBf4HWDpxtUMjNG+25yHLLSQ1ozOp+G2eykOjhlO5
1+oS1oN2m2ecMDEHwrVE+ptd2M4WdxI6q+1LHF/8X6PWei7OwOH6T3aXQHM/HUspbMwpDAaABuyx
hfQ3Lb8wGrV3b6xro4Ys33igyLFucCbn9sJJ0QqvqxhpbHx396MgamLnteJdvCfbJZ3XPcVlYYNh
iWMZUj1OdyoYybzVaukSXk4HxXn6Cx86ZgoeYtBEXntO0HNFuYyUFICSrRl9SREC5L2Ee7BRRZ/C
qOdBpeZNo6Yu629ZJz2LM5P/TT85YG75s67KKGaVcorXBCTgl/oyHt0fkc3V05tHVzqgMdStZnXe
aky6gWnXf9fvmcbo2LbbSCY164l9ZkJixQIsk/GBGrXB93gF10qrH3DAwW9IvyKVJ/VpPLI5/NOn
kmQFDE+tniXqdp8hxeKvSYDxn7owDAoEMyrn+EZ06qGt+RNcNYSe4lAoBOoAu9WxN+5+z6t9Du56
xUGgxdeQw9YMvgJBBo5o4IyqbtMaBBwiG+0S58KsnCMSJa9cwOhFO2mb2WWcfi+kyAIEDqNwS0r6
qYyz2SWrTW88C/TRWxCeDT/Ov5ZuGGEcXs2B2Ejn7ynmq69NaM5AlAg3Oq8Fes3PBxowJsOI6B2C
e6RxNkhP3ViSRpd39ot8E4m/97OCT63XXwDzUBqTJG12m4nYHkBBa+1dBpOX7k7zHUYNvV72SOHx
1d3rYFCV03g6mP5j3pQFIRMpzs9IFMU6ueKIIlSGPX0crwgU9z2M42AQCDFRCohtlwOn87wUAo/+
mGP57SvDMmS4DvE6LL/3SMx8Hs4wCZdgKKbv0+fowdIWNS8AZ4QpGxhgU2AWhW54peg2ZSF6GX2Q
6jjOM2Z1ODUBdd7HKI3t/jzRiVWRfYvY/kB3xY/HhaAPOgwSReJEai4oq850F/GuUJOhS7KXgzKz
7GYOqO2VyKpG81DuH6YBwvLJn5xPv+OEUSXwXJA/GWycQUMMTmyt7/ZPPv+2QEVF1dZszPD6XpIJ
d5U4VP5ZjtUza16P8Qi9W65CUvCR61ISorg3eInANt0e1aMqvH8I+iRSuDqDOKSVa0v3rlJpB+ZV
2AjWoiamgqHxGMsKG+TAjpsasMu8UUlHw+SqoKEb8yx2fnfD4Br9wePFifpDjO9fvneFNBGBPcC4
KHKgFHGxqDnkTKt5LWIEWzIuGdZ/e6CpHt03ab2I6Og0a4n3DxcLxJSgqFp8wdi8BcTJnuqjJ5mm
+AoHG5MWni6/XaPHD/dty5zuZVeoJr+cac4n3GSK6PRbA0UFSBkTq4F2hf5erJ1oVj9RuLkEtFib
JDMSGeyDIV7h0orrgRfIQmfjaPD7iisSH8S0JCEtd/k2nz5Ybyxwm7BJHrPlXVl7Ub1StYHyrgJo
6NBMAwkd66wxCytLKiV29yhv4Nf1QENDgb+W2iu8zKCESmAB93hUwsZXJEzPry4OSJIVpPUvOHCa
SruDbbOiv5Qtch0I5WSucbhjwbLeue9c5V9y7dxOtI6I6XuyHlBdghsf9CUE9mhCncOS1nztVZlZ
WVoRX19091Er1W3oOHSF0xEycxnaYSDHS7gAFMXrzmnYixGwm7l0yE8Ft/UNgH2I3L5aOrmqoh8S
dlRxQ+K2ADNukQqqWmunZRYDIKRKMtyDnGirSegRuV1hlyvFXzqpKuwSlA/R2Z4uNAVjzmizXga2
53NUktlyb+a5jwh2pCV6RsshiYciiXEwziyvvfbaWWGUD3eXHN7QkdVFsauvBNKHkdBS4ZFk6Z/g
XtnnFmiecdBi82VAhQLulSCQiovesnh8jh8aFAPIC7m8Gt9yvgH6G1C+bCZ0eQ+I4sM2W/YkM6NP
e3ji1pgFFwpJXhVU/cA1yRAzaqTc1ft9LhbBM46/R3jJFY2UvfpYgJo79A7T5RHzzcGDMJhwGVJk
jZTNq1wqvr1v8G4VWYCb2b8uhSMOqdNYTZtnGRb/JiIonnGQp9dSjYa5yhA8aGg3eRpMB1k6otfh
ZdglzVMO1dU2kg10Xr26QuWyi/zDATaYqGwk4cXucjKb+XCKbOTxYEyVhpMV9fgnUSWFGKCcfGd0
iyPps/bBjJg8u5SH272Z/JvttDu/SHM/n11mKAOf1uFreeAGgs3u9zZYsDbyetjCRz47i6e9EmRH
01iqaV4EjzT6/2NTN/wnqF2hicvKQTUnlG8iCUthKu9mYXjQ0XmhTR1H1vWFdetGDRBejUj+GfUG
msp00lAZTMYlj/oitn7O+HRlY2LgFyxmN2h2a3s1e89zgRjWxGkGZo9RHM+nPGyBVN9fWVOrf4A1
x4hOA8+suwHV1bbQv3MkGgvyPk/55batblK2s5B3oOTt6i17GpVush8Vh+54Ts3e1Vi2C8Qc5rOa
UBerw4+K1gYkY34JuV/JKCdUuFijdUy2ab3EsAOJ58bEKOhGPO3rU0lpfg9m9vwCun8+6YYJQykm
bHPF9dKrKnjHLk0U3H/h4tFAthAeM0h72U32cVz1eZhG5Y64RW6aNQ0KWKyKol01KB0oM+Nvy1hq
7/EAI6FZojJ8+0tsU0xXSh9kh9KC0cdAcSHqFYtZV0Wo6OHwOm/cFkaMd4PrdxiboBCfFl7cNo5u
DtmXm/a6Ts1dXJFEP+RQsVH5j0C89Cg9H4+AnHV+6c5FVafPF4Y1a+uhIohPWRviSwaZ5DYU6IVL
2lMmi5rfLtJid1O+whCmjcnMq2N74fgZSOTGo4ub3krLmt1SeE9Z0VpG8LjO9pfILpDrcsdJeRgs
fs6p6ossNPZguRst16tuVQa360GxlVK1T7JqACg0m8i+7mxtlpOunlzhFjb0D6xLNbkJcvvJCKz7
VVpDbJAr7RsahRhapGp2zAqKSe9cpSzFR/P12ShbMAaeMOEYZr7VjmY2iC7u2/86leR56Sk3/OQS
kZbnk0iva7k+DY3erOmvyhxRY9xz9MpDy5tU32ULds46o0vHimzonart6OHd8iPSf8QiAF/Y2wh9
kIS+W9jInne5GB/vkN6FHQEetoh/EBDd6Pxxr553fSHGJwTpvacQJk6BnOurnsBtmKGc5a14+s0U
ypc6ggQYxZhRO6ZiDacZk+eUs0YpzzAkht0YxaLJelqKbfgmql8MRT1oY2633uHviL8jqyutMisE
6rcthrcwEXVDXb3QN2trXT53WG2q4lbfdM7h9xJn/CiRJFRLWIVr3k9KJclgS+jsx/nVc8RSyIsE
79ZIkeVfzcOkMMZu8ylkyKx/e5sPleMjMWTAJ53dLDNk7bZpqSzATzr7z7LUioWSZ4i0WVugwshA
xQXW2iYdUDMDWW1EmmXUuJ16nK+lBCLtsu3ywqkfpL1nlLhUdcx7zoyyOaQRDWqZDLpiMml6yf6x
7bqHFFMAWYEpUFm/7R6VoKboozYQcLn33nOQt2hYDAGZ5JnoZzzUbKwohiOzMhFTZsOuVwpKHT7z
KRF8v4WPAH8e2yDQK/rbIU0/CO+6VAk+Sm+YUNzE0/rnQl0ls37d0QeIvI4naJUJtAZupVzhXAWy
iejrp1pRe7yXgk2j+p5pY/1dkDg57iPDHk/5b7rujYVp0KSQyETlNsRx8rn1WzhBfPls3tjlgv8d
CUng3X7J7ff3CgrghJHP+vGH65QXXtmOH+twrhzfHkJzH255QPxNoTJF2CKIkESx/OVjTIubSXqa
lB/AeC0nZpbsvu1FAiwQhrKXq97GG427RYpbi32Y0bIc1EWFg9okHHrjeitEI6MFaBu2Tg4Wy6yE
x4GgX6sUsue7k7sdiCAeg8B7SlfsYqS6oP6QWwVrcqgamM30f7bPoTaetR/Bs11oG6+1bi4vQcsv
SAlVS2NaXOfafdHcp075MmooOFVt6D92W9U/B0uFpXCD3XnvDjXYiLIwrUacYjVaoZusUHT+6VDl
KdG4fweHZ/MIWkqYIm7wMXo1WFak53wJsgbUT6oZSPMfj0SwhAF1TmIziUPtqN+wY1vniW+f12zs
yU69rFUxFTPZS28wGLBdRw4w14p5vMKx8kp5/IX9eRbSHX6ug0d1kb5CqLa+FigY1V6KpyphMmKz
hJc8yE77SEWKAO+/9MnFR/hZlT2RSu2Jx6orGr1IK4N7EWtfuftSsFc7FrKMfUMBCZ+jEXXm/Mwp
1UeGREISjf6ZOcnd8da+Dcyrxh7JqOMecWYEv89kgoOM2lcP44OVaylfEFR/N+YTwdsSqYF7bdrZ
fOEEPMI8i27dXaCHnqb6Z5GFYGlVvyKSEKj35VcCMeTBTdLxrXRAp+PwoDjnnzjdAHMBDD87SfD/
LzHwvsQRcvxq9LIO114m+syG9bV8LC2cgTjb1CdMq/oX8YxYt2YQ9mGZ2MQQmZtyA9vXVWu9c4aT
AGeYcN5cY6ogPU/D60JXHbByQ9e0rzfX84lYfuS9xroJj8gcfu+w3rYiU7kx8Mw8+gRoNGoMkHMK
7Ot/yBlkPzBGoKc379HO+J8bY8MGvv0Ertg+c+3YE4RVA0ThsuzxErndlPC0CKTdiB/l0OBr8gxY
G1NMgpsDJElSz3qHfS+NrOv0BxJ4J58rJvzYc7oreMzr4iWM2AfFa4iE89xfuFHOBc8Lm5GgvEwt
0gR5xC27/+nn7uw5EtU2g3L+cOXX8T6sFWFXPS3ico6T7leHZZK3jBhhrVqzUqZXmqKtRN/G4ng1
L0jG4dvsNegoNYxXk+zoEtjPhe1oJee8tR+CmVkNoJklV/UKeC9RvmKuNNsTuAMVEWkRkPNfXyoY
aWHjwv4ARS+ix9JFT3QdM+jixDJO8mgg1XJOhhkmQc/4rfqQ9LUaebhnlHDklqAMB2pw9aseAnDD
Nb3NAw7N9OT9ATwaGxV2OXtayHR/bOgiFeY2L0Gr8r1jN9QAeLj98cEn/DFIcV6vFhyJeULvBlR/
EESsQeHybqAS+9Y9fvfvX0N3PcqXkMwWmRnqzxux6aRu4uF379q4l/5TiekE43JciEJ3wMXLFmrW
TAjuPnioU1hTJMJKiLzjIn4dfP/wKTsm+2g7V99fbp5yb29wedkV9E296UCGhFrKU9Vdpq/6OuGN
6T41VXiJOdtwdcpovlmkarFg0hhtf51GnmBFIJcMWNQ3e+keOcdsixO7lOHf+5ijaCC/ptvM8PXp
uMrcSQT02ytV1ZO4W00yvcR5dIrvl0lRbt/4QSt8ezX+uzZlI2JVFW3PYxTK4aNAlAsHsNaPcD6d
6dbmThD8kLSzkSmXEEuvZvKxQuDUVv9bcRz/uVtMXnlXCxhYKLNZrF4MVmQosgmKXAuPUoaxwnKG
oy6JZ1fpsywTT4M76gO647KyDUnb2Jqtq/5r/bEgSx1db3YQ++R5whfVH5wXLryVvEAfGJSBMfPH
26eCfFw/pZrF0w4uL37UL/OUgnMYLGsKZdwH/bC5FOyHQDzWD2/vseJDc4DcVdQCo1zSC6DkkLqZ
9MwUe6wNUSFLdUJA5GQMgdOsO2HRA6dKUKqWECBtYoFpvvps5d0MQUvZehsrr805zctIZ1alnz4w
Net9nHVsd8gXOadB5r41VQ14+OSf0ELGgplrR6nKUmdt02jbmAkQ0BMYfrhjQKey0GM4MTFgou8U
YvOJMFwaSNzaMRanNh8K7sElDzvZj39F4/g2GNgvSeAUjBcFiwLfAVLyaIZwW0he/JbVL+MWa/Tt
NqnZqUZT0RnhGAd9C37JqMsRwZhOkW4LPj9B3KdtEwFeIuOiyEYB4JQOANwRchTXcZGoBhXwJQ05
JnQ9MwwAJC7OZwfBWLTFVj7tjKayoqtN0P1TUgexaq2LWbO2yY/zS/Fsiem4afzP7yCWyqGh+Jk2
L34HOiHXdcAUQBw20WAWqBpk5Ps5SzNLMJ7zkKL1ftBVtn8WUdGjl+9Nuzef1N/TFa0lVb2zON6u
HxwVgeKZQGhOGwIOWyxxBvokKvuZXaTTxma8HHXxOgb29gyxI3MNR4ARSqeeGLZqiOVFjZqCDGfh
1NdSQoUWEjaUsro7jYKAhRLcFnFNuaCFR8DJTemoyJAyxDyJ+l8dscrPi1902RRi/k7e3oSuFKOR
pORzjD4efeWGl417P0XD9Qz/DciQJG/4IXFu9esmjf96upX+9/A9tOxF8+c2DbkFucfej5rETBCk
fLoLx8ZFvhRxuHNeGnZr+r96nqrucH0XNBiWMn8byOzcAYgY9uCLoTbKquvDF0t+O+yebD/EI/0Z
TuC+7xJVuWTCNlO3eVYGdm4Sub33bGJp22eDgwDMcbNwJlX1yHvQpOgo0qwrpdNgTPJ27pdrcRzj
g5/56JkY3oMZcvqMqu8s68mQj2VSALOQhDhAiwYKbiZvGBLfKOBU0TNqPc5t1rvW8tzzf6b0fEDD
K/nbIaUQztPY8hZ5oJw4CwPhbKR13K5bnb/8ny8Ny8FgU6qf/Wu2hnkK2QrRschk7IGX5MR1PT4O
WXDRHJ2dr2qCmS0cZ3g0/O0dZbXu/QcZU7DUb88egdvgnp+1l78xdZaeUVuLOJ2ft/XHFm6vU3Or
YOfJollhUQH4OJ9UnHLKDAiJQGEruQ/fiOd8loPz1I97g7wCqpLBEQVr+IASOUoPhs1AsDhUu3K+
D1sWvjdTBQ++WUwT/5vTJBnwvbtdmox7QlttQJn+0y4yQSJ0lk7KECVKWWEpKEd2cNwdWbOUypKi
ShdHcbHzP8b7u8XeUZHFA1YTkdTiq7n0GAfHz5xwbVo/ZB5i68uS+IrjdMqEsQ6AprO/pzmETKgC
xqQce6CBHozMvv6e9S1t+U575Ns/8yLSHJYjPttCnCqPwhVW4HkYjvgy9KLET+lB8ifynqtNTSah
eLwuUZ9jz1voeOYXcbPeBPe2U0dAe2tGTplmyU6dvFNC8OYwpn9w9NrdCpkp4K6J07NQ7+vxQWjq
JfHaEqu0mlmE1+X8+xli4j09D7AvcPS0SuNiWql6kjN6cQOJSLy72+gpdKJ22q2qUvZs0fPOilQk
pZvJMzNFqdIGFWQbPmPbpOnbvqmxKrqdJPSORE1dmJBFVerN6rTxjvptHIyuXVqvAGw+U/lmmwQb
FyhUIJrq6S0CaWg73IyBgWk0QO5/aTIqSTfYR4U6Ozl5wks/cAPBA4abZjdu4lwTT4TsP89X8J3t
2Iq+BV5HuXaDLWL1ug7svwY97cSZ8ZyHFaej/ky1O0X08u2qo6+WQ0jZpYpBz8KEYMA9ezjdhzQQ
D5Qkiob2gHtEz4y6H1fJcpqECqghwBXGSNcX6sKbAtQLybYZC5X+1oXX48e/c+Kp8PZ8wrdW91J6
UwuXsYBd7tYAgbF6fVKSJYXatJ9sMyuAkzCvEaG1YUak+hRz12ezxsfdHZWSCIdxTqBa4DTtnZAp
QchovgV9BdHeF5D1g7fkmP9S2asVZQ7GbsB9Xsm8sxCljlFKhRi8xvkiS9bIUQDaX2ledQD5EFa1
tS5PQCRV6LTOdZE5rDrLOgDtEwHwsvNa7KJAmWe/To6uDvhkrLy1u7GRvFSTqE+fR7gApSRP5UCE
tYc3TdKWUoxhCK4vGjZqUQgcclMvMLkR0JVIYaDoy5Ky6S9VrWBi/6yrh4PLMmfHVRtDVVdDo8cK
xHbCpuwNeVtnN8qYff/204yW/WuL8+gPHoa2yxZupy0dsEd4JkD3Bw0V3SI2UX9jpF9CSMcx9dPL
qtYA1Zja4KdvCRBuXmZvBwgDDEOzzvsuZ84kAQldKICYJPSsjNRqmY8pW5NF/j1bSXFEWXSjiLF/
uvPljoKjGHqQhQMHqrIiwtvT4XdnVvSflVuflUsLXBg8/vtSvNJE2DbyEbmZoNGGzwYtyNkdkt/P
L/WfdN6OWM3a/16wGqxix1iA6tkkolZ3S5lO0B/Vtn4CfQveHT8jIetVSuth7anlcrTVJlIq38m8
QRPULLIqLzwCZBpCighTiKHf2ZuPlEjl0b06THYXWiGtyZPaBJrBuZcdfNdI5TEJf+LVwz6TVKFI
uyvrrRB/7O7A75i3TC7xGqmJeZIwtkV7oA42Fo1o3iCQS+3UUSsa3o7QZr1WrXp7CcW+szbZHdY7
S45T3dDJ1uGzXskz/VuDn3zdXCua5fB0hlTu75dhSB5Pe0avkqDleYiYf1A4n7llNWlu0qot1MdA
SFZVQ693+UFBagSjMB/oIY/L1ncLUXz846fgYJ1gnTQtErcDxLlDVYXhyuF9EjUpfQhVxToG6htD
hK8j9l7R7EVHAuoB8ZyXhqD+OjaVo6xx7UP6E3xVfZ9QJt/Zc++XAxPA0SFMhXEOO7uQMqZXVnRC
Ue6lA3Asu/XAQHRMfJOBP8MRqn4ejSWSE2jhzqhfiNP6Bb0f+kUHImdPxC9GCMxnWIkER+Y305ZT
yPYQQiFv7ygZhn/OoJGToAztfO7yFlB8u/+EfgbDgiIf8XCMuzrLOT3nWpbXJodASZ7NmXq4grrm
/mNuwOkgiYZtzdBie70G3uy0eQas1xeU345O1A2gM/RAP3WUZRMGhc94YAmgWzk6sfkD5H2GXs5g
UHL6ni4SvYra3ny2lYpE+/8MD1RBqEgPTdE43huqs7aF6W0aPj3WWVu5Fs5zGXzrr2Il/2XllO3R
xOiURUIwsIIMCL2F+OIKl/bNfMAIe3M+viEDbB3kfJ5GYTnMT+mHxvG5ddN/K9PXlPE4DOsAOmMS
+hRklhQ8JXa5vVkJG/fcoVs0obOkLJEtMMcK09B9Dpz6uv/HgLj4djqb4Q4VaHROj3taYPSBG3wf
kdhyo5mjOXK8Zo2qo0CzZ9eLuqaTRfZv7qLyOxaQg4/xZHWiWX5YazKz5Kcsj2t8GuoIWAijAT7L
RPPqXB7OXeD/DJunq9haS28Mhkv1uK6HQ30jXNc8DYXA/9CGrr3h/R/oXPA3P4QVxGgfTLa3xn2B
gwnarSKR8rdtgkMULkaJVlcvxrgoGsDyqUbgrbKpGDAcVBE4xn1kMCZ+3lWfioMrW58JJFQy3/wb
k7a1+QHqaJojhMjl1gPRnZWpuTNfBjans53cEXkUHmn7gmupUfCkvV51BMzbs/ZTkjAw6NrCU2E7
2k+O/PyDsUokx0IiAJ8VoDQ9R540wweODSqpT8T1kPKdbPCS5g0NEStESDNc/GSUyIkz90xbrhaG
n7NAw2ptQW+wRxWgZiIwGmjKv1xxrWL5P984txZ2Qc9qDH53PsaWwwpCsiPHa+sen4d/RuYgXGOa
8e/gch3/YhKICLZBatIxbmxHOAeHp+/8ZSOOoRI/JN55c4Oi4wbdRvjvkw6kwhkJJvBjZIZ+ERjc
31sI9/zkGSV7la1NHs8RgXSJtplX5nuQ0HZRsoaJlDCka5kIJll1Njpvr4GEkeKMD39W6w4pjr+6
FWxfZozLmNRdBWN+Bfl/NsqwCT9V4kQOHDUVgUH0uj6ygO6KPBAHeeWOjgpB5tZzzpz/qx6useiV
4H77w3qZvjhNwDzSxs3mSFSdyQj7n1qsg8Pr11PwiPBAbgB97sgxc4BieTIOKrBeK25JITYkoI9T
4BSQ2yklZC4oGAJq3KqVRHBUmc4K5fa7H1EHUbOZ7Fi3v0fwlx1qOwqHi++pk2z5Yf/v+e47rbRr
iTJv8HjFfpwMkIMppZJ2enPKiHzVCNNbXeU/BPniSd5j2Kt78gSjvFF6kGYIq47xXLNp54Wt7foI
ew1zW5jpfUCnUV+izjU6ASqOwmoHtuEnUOf0IfhkQ1gDzgnmiGngWNs9qxfLOEuV7qP4QpDcTXAf
6egjmYqAekplc542RBPe4+ZpT01TpaT9YT4dZtH555D2MIfWxk5LGAYu/+1tNOM9T4dgpOcp6OA2
1WUXEqg+E5B9JB5V3NRAEGVbxGRXWaX9So2pOkR6riGtQVzoFDQKclLPW5RWbwhp1MPIpzHf/lhF
kNENzozhyvhsLTs/g8uHUySWBp30HT3TsprtOX3AZ6YaBB42ms4bIJBnSwgu7/9z0w8cS5emwHXu
C+ZqYLIvxk4rAr05+CO3VtxBBG5mwTOO03Wp8pivojvDOfIqUnprblKPxalEReOb4nvQUT61suuV
JU4ZBIrLX3Yekj8YX5pKnHxwvbnt7nhDX3d06HHR8iOzllwFugrgov7yVzvL3ggy8oQrtXrR+LIX
XQ39zKojO5O+kyWbdtryc3JC/2qFIf3ZqI1ockR9L+YBCp0c13gyJZsOeX/tVSjGrHmsnB2bmeAD
6xztw/oOU5fq/OJhMpQW8AXZRf2SInMYEdrWhxuLrzswBD+nN4DBr2x8YWHu566r4djjPZNXQpRF
U9FfGabFhaL+XMTlJrnXSWADZPyDo6mKLI8pIHbQqMYiBWkNHXIc+dYWh2ZeEg486sL1neH4lhqI
E3qDuFP91HPS+B3r9qXdzRsMFXz8PsJsZmWxLceWL4T9UaLLyBzBjt5HtYbkZqzsncCV/3nB77XM
+jfqDC/yXep9dKH6D59j9KgYGvUSMlENI9UN7z0dcbL8+G2fLF/1yWSGq7I71/2ORUGPa2j0zw0E
Wk+ITaUCvSEI1daOKlU4xqoTY6+TB2C47FaGPaSp2GiSw/F9ngdYaGXHAx2GvndWMyvotBigVYaj
YwTwYpMPt/W7rs+WadVZ3TmbaXvxX8yQLeGJxc0+moysE1FnTFIXJ6b233QrD1Ui0QdYFEcx89Rq
30LUCmE9DnJRHBg7gAjKPmKz8ZPl+PFrzzkaXNAxN8CbPERxWAc1yIWHvodWRi74FwrMvlFghe3V
CgU4JPtP1tkDJiOvRqXfg5L4wbVHWHADFy9bR0siXhsjkt2jbE7OBl8CoiSnyg9y0VHv07IQoWWp
JvB+/uPpO+xAVU75OJAIZ9/oHYf7Jnt3KUThhLbA8Zoue30+43Cu1wLe5dM7voPjFUfG/7bdmINv
Vhe9GZg8N5AXgYR6i+H02tb3DwhwLhacEWbSMJxS6Pw5+VwhKP+91YQm3UJciovzreRCUC4kDeNU
W+u7flzjeb+zHxx2GNpTCTEbinIvTXDYy/STYK1yK4eCHfKQeQ9tglQCDyQvei1K6PtJZ5i4NcLN
5WDG9IBJWl/WnrbP2gtuY1AriDFHzOlgKJDeM8CnB2f4R9jxbMl9QbxHBTMdSGt7V5++Ar6xcp/l
+sRB+F+R2BTyDdDQ1HWXcz+GlZjwNCfxdQhre3uIHjSdJfkL73lXJY89j9L7stCh0mW6+xl3whNI
9g99fWVEkx0lslr1lAMMEkaThRiF0VWS2VUwyW0YbZnPQMKZplZpUHb2Kf4zgAHq4WMCtX3hjro7
n3vwZ8jc6/YDvd5wFqLsgMHGPA21U/m8StFNcxu6IN+wNjMdBCmS8oTnzZkOyhf0rg5PH2QhlENA
qBb/yy30N2lvqQkC+QUhA1Fq5GZlcXM4txmXrKblmSIH73U59qfGCg/byPlovqRqKJBjouTmzljz
R5sBeDcEMt2++ggb6G1pPMN9c3h8u2FvSP+eiJJEUqZl1/mAL72bHlq2OEKS2LePuwhlcR2ALYQh
OOjChbdpn/1QKeWjDkbVXYyFMM0eBpx0AHTK8HDNH2GdTXlnunoRLdkxTFvo7Q9e+lS1cMy2KeL9
SswIul7PL5+ig836L4O2VS0SMd4u90brLVKaPD2Wdh1EQW8hJygQ5ZireSxiEahnIaE0T03JdFBy
GtheM19AOqW7pRKrkKzdIaMGJJImKFa+dMttWra+SKjZA4Jf+oLm8N7jpOZhicWxc/Oolw7YDqpF
MW4WsJvsA4+Rpo3fhE/nONKwBs9Wuwu0djyZxNknE1eAiKR6b3S3NaqdkyXTgKqBlWvx62XaZT47
CauFVFAsS9r1oJergvqb5UPPs+QdhSYdmrziZRaCVx+4OqRva52jxkVH/CeUMYQy6mAdVRomZ+F4
csw5E4zK4jPEd3aN2Rz1M4J04vbDMCcjTzyMdcBhjbkv9BPDGpn8hrKPwzSGi9DTh23dDYxbNlzv
1LhvbtQLs6At6Av3WR1PoGLE9TPPPSBNwX5NAH0vSjpkocutcqne2m3QJyd2d8eWwXe4wgyQ9BTG
gG1ioerXMGifeyyc77nXjMnIe9/+Qi1Wtd8inqGrkpkK0eRdj90sKOiOrzsOSY/NrzmprGnnGZns
msf6wDRsaEJoLtagLWCcQIcgblWOn6DfSxWOnR/Tem5YM3/f5jjKBXvQSPcXHQhV8jNSwH5n0F+V
tZXxVnVDE0luWQpnjVE+rPGlEYWW0WUm3XMD82qZKlbV/NILHaKejC6KExKXlVVZRdp2EFfcPNr6
NPVhNAQc2UwsWOgTthSgbp30t0aJ8v3+feZ4XW/OOuZoSJnZdperzzVYqBheW4CWcZRdn/XByAd6
tPicUmq5x1T1VL+T9sABnUYr+5vLVJcCGC/64ZuH44ASwn5R5Ogimx9URKASXQPe3e8fv2jCxOdD
PAt1JRXU9nINhKUwSMpA15ygREE81hAnRuIvmCE5iT+xCW3EiL3TXpqGMBv6HdVpC9kG2knUiuZf
m4VqWJSDzDCylO2KSfracLGxOAFU7Wp2Dg1o84UhQT3is8zmu/EBTpsQMXZhCOZ2rE+gprvVf9d9
45v+rKrpWHzTNIQl0HrupSY0XOWZQDuUFiyz76NKzIUwUY2kRqEtnzEzuEkLa/GvxinyVCleanXC
o6gAqkJApm65OK4YtF1SDWrCgVes25E1zz9kvhzcmBeuNGLCR+jScULPm+A2azkiWIuu9axM8XTj
pW3dV8toPSbrBNVr2895FTMJ3lUfr6BMZ1+u9tQSEV932mIM2k3vXMnxuyWoL2afTFhXrqxfTNX+
JI6qCf5Zcv8pcaNRShZ6NNgAGHJmf8M40Y0XnfeaL4wjYZqQTe/+UTSrQdAGzN4NM9pQC4NsuLWy
R9d366hxZiRR6vfkNJzo0EwrKRMC9DTJSkDtPqhZ/YviNrUXehnM34BvPXzgWn+xaiBSUxgsOXlR
tIrp09iwcKrsFrIoFvKc6Bf6zMvtUuD23AZa5kuhs0sXuzWoBfna5cvCd/uPS8zfmbFM6XTFWKeR
vPKam1kBAU4zoiyRLzh9JcaJ45YKKBaW9hAhpjTE7q8B0KG7/27fJg0cqyV09FXyEj0B0UG3C6M3
B6HJs/wxSPwpnVIK2kystF5bQouS7kgzCkybi0li4dn/tDLg+Lp7D9rEtJ28K6BlZI8n+rHewKan
a4JKfWJen8mGQg6Ejge5JRXXzGyjNwmQvvEI2fLKzedo4Z1vFnPtUu3yUZBbKanG/5C3x5V2fJhm
v3ww7kPqXOzxnQ2p7Exw/FoeBrl+zN13jrFCGMMps3K7SSqWkYNEMl77qr/J+NHdMPdhxje4UMZV
ruJtCmdnT0+YLpjXf9SNH1r+mMFvC+74pO3XnQnfv0bSzYdZaUfjNrmw6E2CqFejs6GXgt/lI2Hg
onVW3MX/6UUigJ7wLdhZ6mgWeoHlGCUfzSUgeCM3jIqQ019nqX3jU2jok23P1ouqcCcCub4RggHu
Sqj/4sKI0xmgnMYagiFyKnc6L57ypFsBK58rgQV5waCMKV5gUQCWL3B8skq+2uQwOyrrEq2mV2Fi
B8bwvNDrtqax5qhYP6Uuuogz72krEOjTH50GA1SSHS5aVi4idia+NRKpldyzzoV1Y6xSXtTOXUI4
mhT5VoHCxW2x6m2Kr7jtYge3REXSAzwvn96dU/skh8mHzt24d1BrQVnf2CI0J0i0PAcvMoeDlCt6
DsDyuz5OiioZe1yXKsC1Vq4THZHYN+dhHrgjSGIN30y7jSCKhQzRdJYU2PgXHx1ZxA19f0ASqchc
oS7p5C3JS1JXE8tAmRXryhrArMBNwuDeVNEpIw68NE5C+z4TAd+QxJIYNrvSvD3u721cBYcE7fcg
LZy6oUP9W09/RGIEm+8htHVLWl7VFBWF50FqFrH42ClHTV8g1KXPwYX+09E6lebIFYWaJuXVb5vj
PlngcFFF7e0My886oNnG8HFCTEpaxobqkz4G/vHL1YFxX/F9OiqPQlbQT+0UayaD5EdagXmb3EAq
s/0HBLDOne8Eqdv++0cpdFqecXBL5bmmhadwqQ+4SxsIIEy532odsRFtuLJaMFKyU8dhyoL27HJM
YkT9C5RpYb6s93D5Zd1f47R5Z1r8pmZ5vWzwIG9cXrUuE1BKHDJm8dlaAMpmrBZABALu0RE2PH3o
kd9BMOFp+lAjojGkx4MSNisb6tv1cy7/C2BV8diOZB0BKHY+fow3YqMd5BwrlN6hRLdmPbW99aSm
znMfKXU0vFe7EcfvvmHgdqXrV3p+hfI0SF1nU67smcJqsznMN2JVTBo7Vi1Q6CntjPJGYtfArg9n
Jj1OdUQIzyph4hnWdg3zECREhiuod44AvhjQ2aaFrJRRkss3HjAVjfRnCu1w3ipHji8exi17hVnP
XRZuIXUirwklF7nY5se9xarMzZ7uhcVQzxdoYMBBrE7olO7wbX2X8rf7PtgACGqealbB5v8yqXrE
/sTslaQExREcv/Veb4cVoS4zf+Y/xVXzXUM6k9lNAPwUGw22CX5o3MWG/DkSqoGRGYgZAarZwBix
jfZt+OGaUTNkTN6rE1CKBiVdclvrD9ASeAoMRu2F9YqcaUiqa3ktd4T5pEkeZtIuTi2dgu3yET2r
mzqRRXf9EYhMsNuDqwNAjAEL8gz5OjTlesy/TJ+f0AoI7NKjQmX93Wzm8hZns7CoJvQbomqyee8f
YAG3wpiEPLFWgBXjYZLkRVZT0vR8nlUTePth9fvkpczqEb9RjGR1o/o69Nu2j8tiT0AHxcVwKCEc
9YW4xaoTVTrB6uUajdAYIIwftJNQq0LC7UUqzE1Tuplai6etU0mUJv3s6cUn2wBbK5v1bavtK0oE
H/d8aZzYmIXPOw2eKr/hfinaMRL0DvVOOgA/lkUeIWH+jzFa8XlXjK8aE/sxIqyQuya9d8YcFcCQ
DmzCcsH9z/y0aZiQ3M32xkSZB64PxwBBbSMcxVyq+w82X5VRNi5s4xjhSNf/3Be7qay4fGjY9vok
4NZd72RGEcdcUwf844qElCuXuDTuWnobpdlsj7Njp8gZd9gF3REshb+bMUT9VYe1RzZ8v/uPtamD
jXhoDNDHcz5WQXlUwqwdRGni5f7oDKsNmLGKC2Iz4foO78DuGCLdiYwIoKlzI/nfXbqqmzQX8RVX
beV1tX/kVr7aTMfZhCS6crXkuSPDZ5U7RF6m2KE+34noxIOFus/u1pVWIF0Y+gj6bouwE916WTyE
e/Y8qJ8iCQa4bcjbkJjkvke4ojShnQrLbivsiF8FAUmL5tKNkMAspZe/8ZNCHWIZPF1aghHNxxge
SHQjUT94qyaDQK6KjxH8VsBWoRwFkf9zh0K6Nh5Eh/2zObKG/fPFgoPGHdg+B3XD+cSm6nLZggbo
1ZoyTI2NoSVZgBatxoGqi2RmYoaJzuoKnueXrYmNyaCBTLl8JAaCOa7innujhu4XoiXtfk0W9gtD
3tJyxMolL5ue5KeKXTbmLWSccpaXJkZ5ItVpny92eZFSmHff8Pbnol/E0Qz7nIRoKily6oQlDsi3
4ds9r2fp6fBsSIFibB+xnkl7phtBYG9jOhb+G9+0McJZMMNq7Q0p6sk7c9VB3mry+anNVpWxkWJB
3vdEcV3gxf41NQ8R/sdPcz0cPjafbKnyg2+pvQg12WChgTZDHB4yUhkUWkF+I+XSizuR+xmBlcTh
3/XDkkPVBhvTwIq1CdF2umiQJtH4D7NX36JDWNaKalwDBLKuU1QCI+avPtqseWiiSIZyUXQ/xoYM
sZCSiTd71FYpY6oEuStP1xrWQ0BucBV6iNHJJzZkiJr0Pk7twy8VlNMEjDK7scP4Kf1QSMLZh7X7
IKFeS3YMlk3xXiao8I1hXXKCTa7Jy/zhduzfVnhpyOlIqY7WcGPUTB29OdLkOawiHgIa/Bt3shq3
dE1esAnjviQgJ/Ivz3GdmqGEr4sNtfUSsr6pvZAKmgVGx6skoDd4uvPk4eTOuFCDNQn1SeztOQ8b
b1yLA8uEn0cVPrbSqEoetWZ41k9f6l0cExYJvgi4tpdsva3mNBOBRrsuBQ6D6VdS8Z8vB18opcSd
+26cP1W4mT3t1q4ntkw64ep9cdSxqHnrofrSwgfxIL+N9LW7PP7QxjdOjYisdsLEufGsKZBZjkI0
G+u9OFaEtpPg/MtUnynsngTvcghtsRGvP3+64lYC5yq/9Msj7HL8HgDFHzCqfnj+nXluO8qEMVY8
Y8CfVvk5y4v1niJ/TGwksZuN5YqzAFwrHTfedABWYj2acvGI+QSbH7cjH5/exsZkYHTVPbh2Ru2N
UUkZBzVSmCqQ/7w3DhNTa1ObP9FQs2ikT14RVDE0Ym7lF5Q4/SFvhdTtftw/ii4DImcP2uO36yAE
VcFB+6rdo5qEVW/T8vfzGpTvWNbXU6of0gl346U+xS/JjEhI3g6abssYtalq+8maQY8CEEDIqbSj
TZyB2SJCaPIqv9EtfOpsBd9eU/vmbk+XLj9pR+ulJj9yGXlWVQETp8yLfw4w1ICxrgkcc3LOqXXW
Xi7j1wWU7xMUjBfcNeQA55tEXDWrnaNY5AGefR+RXzU89K3GlqptE2JSYDXE/8TS/hOeeVp5qQD4
h2Mu56z/96XsPEevFDg9+2JZTrh7K1rpEBPy2quLDnPpOIlFwLJ0jMPfCPjq8ZFZKbBame/JowOo
4y5HASdDom9j2i1ww+h4Q5RMbBL7OD7pBcF2SGpY3r0n6EP7w8iSuZpClnkUdT/MHlHdeDerV/HA
moBt8wDB/CvwznGNFukuEvYe85mhKqdLTfGgxJ3Fh3g9BFa7Bdy4mNGQ6kaIV3mbPdMAZt27fxLe
CvhQ8nQp3+VhNWltTo+hEk8jdSuJoXBrfxEbcpDet/Ju4ToymMpodOYwHh6f1OpnUFJBwa/wbogS
fMsuSDUocm/n/BzqOk3YzJiPlfWVfFil0YBCliXoov62VQybG54QzOpiNc5gK9RzzFzSUZq4eNc0
HBtUW2gbj5TVjzmednqkSxIoZ0ggTsug3agS508TiLspZSggjxiznx8l1+lJfAOelN6FM/FYhvIG
vp4tGW1Yct2LbCGWQj6BuxGtmVJyIplNGyzK2tXUnP/nWi1sp8SHIGFzbdNQSgUeDFgEzOZpMfCM
DcCisJAAVkb3Psrv5ftvqBRsRE95yvVin1CBIMQRWPDoBYIn+ty+kvPQc+utjtFqUyEtuBnhZAZf
oIjeqT2zrCykAUles5aLjwZ0QqVCBSsByaUX3+KKWz9eIKPB61Z8jQv5BnU4jko09JS1qSl6axge
peFF6EjNndPJciBaW85lp1BuF/foaDoXj8dazUs7NncwOATW2fxRvyvj3/6HaJNe9j90QP8sR3ZR
EEshAuY8AgX9Rf5vC5E2KNJ/ZcB+/LF9Ud9uLsrAIo91Z4AruZ14TrX7O/duP7UVEf4Rzpi7m5/E
0JGeGdB4jR7FwclX5do8NPHmTI6HwFp4dZ830+vMjB0N3OSg00XkOjJ3vKSSweyGDB7TLaD1hkDN
FZLmzdp9hB0kibN1NgThfN8z2oRVL/jqE9Xo//V9Evfjjy0tuVy6nuKsyTfhMfhxWIjXZKFm+NLG
V4sQJrWymBDzlERI3a9CePPBz160R5eciLDupy04dF7uYYmp3JYlwFJ6tLVsLhIfNbGXAAT0KLYa
cXdzVo2dBab3hi5GjS2KuLDF6I60uopo1ESEHY4aR39jy6e0n5bQgghrfRI5ven4mUghGXqPzI+m
mF2XJ84lo7F9gfiZAUqsCrA3spdMcWKgg8Zfms1Xs6kCkDB1HjnykPuTqNcLdK9iCD5SUaxMKn6b
1/fdx4E4ZSYumyZgHt9CjxOchd7nYE1tCz0Hg5O2h8VJ6yji+rMKVCAaRMY4yHKJYQwwQAtdbYwf
9zNa5/xIB9cQssQVaEoybQDdVcSPp2jkgopr+rWtXg2OGDQD7LfEJgcwyM8xOZJ5ruimuXilC2Yr
UEdDEXu4qMWld0fMMFccxTGaemMH8s8Q69UH+ktOAiCIMAKgBc1voPrLCE7mPOVOil81HO2FICUv
u36l0M1EamE74DLkvWHlmCTjnF7/6jnOWcMHgWrRXABDOLbRZEdtNcm3kCKjB7bmiEJHk2jzJWjR
MAfZpEHnmflzLdwI72iryNkZ3N5CW3ubsol9XzHyx55m36SkBrr2bEpyZMQGiSkqDcD6i2vJhXZl
oEOAug8BrPARbYv2PkZmGiBBhj7ASzQ8TG9ic4/VPIGCqavbv2eN9+fOEnpw/bONByj1Q/HugIwf
NH/q3G4ykXSKzpa7A8sWnO28vM6t5vQ7qavl7Cy7ss7q656jSZUa6pN28R4IOhvoqjdUBwAfeWMJ
qVhty17Ihax9lNojAH2bHlhKKIgsHZrGZrU/Qbzto0+LMHtMFVKPL61VAVuYLUnsYBQdZvN9fDu/
E0sYp33CykC9yYaSdn81nTE1dS5divpSrfpNIqvYz+rWng2hULxn6Ysa/BSx0PNcBIl65KkZ7K6Q
oV/qRWwVIc0YPUUJW0eax3mqmx35cdEHp/WT/FlKfE1e2MwGHVR8o2HBh3Yd5N+wczS5QLN8/YQh
FhN6CxTgoulJhl/hOe8a99sk8uWw33kEObII6ITSY2C9WqwDlSjgLPE8Xt/YWRgfXylAU5L242aL
UfkIKz6vyed2m6o3IlWa/aO5vQUqAmirkil20uewzFYThfll4+TiGWPhJs7cUsv7Z78ezQx0tMuT
GTf00HC5NtQFqFbFWT9JX7z9lFQVEegizoF5NFlHdtOP67c1WnDHtkWhDPE4xB45bSTzKmt6SOZS
UJGJ0uRzy9gr1ZRp+lrNCPQD/KkW/8H5RDefiYyktzlwP0me8+nUqKrZlhRlCxHmOJQ0uRxp6nnA
78WAD/056OYgu8tBDfTy6a9UIJGBSkacZug/I9XdTNiMDDC+uGdaw9XOS3H1OBH3TaONQi5lzF11
ucDiVMPcC+DhDPAWjzaa3MixWZc2UGnlhyM2ovZVRnDpcwuiYq1AaH4vYozW55pcvYp+kaA9VdAP
NHjI0gr3j+Z5cGtPCEUNa+Ruo1oydGpPR9teWrXg+3WG7/zyCS9YpOaK20P8Cz/U0S02ZxsKP/G0
gvSpo9XsM42nOLk8K5ycS06VbVJn7NPEQOS3CwcwTdwmo4n2gjK5xU9qBkq5f9qmTYOf0l3Ebb0p
IhiRcqV5hN1+ZwWWzv7yqDuwHxYxXyGIvWQsDF6EEw+TozH8NtLckhePm1e2+Mgw3EcPuSS24MGA
FRnydxEcbhjUWRmm7v/mtLwU98mpHPflTzoga84+Nz7F+V1YgH9yYmzc/kqLdL70FV2K+IRT1DFv
1j70lftyBP22NVfaGKSeZdc/mXeyLYtxHamK+yP+WM/P18t586w+sF4YPU/jsoP0TFC0pkloWHrH
e0p8Nt6xWZUayWQYGd6pvT34G7GjrkviAp0pbM8PEN8iQGf0d7eb6RAtndqOVaczXR536oWwlzYS
wKwRze6B580hdO2nibgpkeO/jHz01nroMT73twY9a2SPxhptaZiMxt88jvvog15GESYYxFtZZm4C
b4uzz+ejOAxv1ltG4dvWc+mCdhVW7d931YQufxlILCplrFeSZJLBf7xvKR2C+k6p2xPOMaozI2bp
3vWFciV3EZRyii37HNraEsxpIomrLCYmagvPGb98kM1sbxfSV+rn4E+nwQqMDm94gM6o4zACeQOf
LmqTxUj1GIA6jRJtIUrvBAAC6L4RL3U4eptqNYlmaUCxIf6PfY3X+4Zo5CulRjb4GCVzXY+iCO/y
+lhnnPyqmGn/bi8MpOX2PbqOzRWYd6Ccpyh2Dwt5xYDL3oOyshe22VCxSsNPhBc94JziKNwayNPF
koM/GQCEDiKHi/aGSU68uBnPkj9yKtsQPXDSMA344rGw24+MEqkj2hMqaqUMA/qyw4VhucpB2DK6
aMpzJQnHAs9FEUxCtKaD0rtFr9Kp1kSuSuLNWgj1qxmexszDGfJwmu5ddkA6o6oNEexSfG7xEsl/
H5HjHuG5p5QZkU+fpb6ZmGPGfNcF/FZBlOVLFPcg8qqVXaESC3z8kLZyBslPcA0Y/P4lOx3/2krD
r645b8y+02jce5IwtE6K9GA00zUb4WYs3vICV9ycaZQXZ0JphP/3vyVF0p6Ob3FkgZXEDV9zxk08
M8xAvlCn6+N2LVmeEcgsyZGRDUhD0AdD1+eVv7I6cPTky6osBu0RdBNEy6da8qsp8TyhAbRmQA1d
lujtAh727JzqtYG2VpCliEgdjZErb3/2HRn3k1UxAJvLij2qQSrIzVj5VwOktKLgi5hQuMhG/kJr
hdWFx1HDf6lRhT/5oq3/beSOoNRNYjmcrKNRtzpkqWbSqb7bD3yV+rm31A04xV7viuCw+WAhEqpc
jonmN6lXDWn5DLvxmxCRV5tXi9f7quMCBYdPNfo1+Is1/lowj50QwrSJotEvnuGw9BCEQ3uTS4S2
2I7NTlar/bBcM/VFWTqS4rt3CXPJyT5YTVtoqcDuW6QaZk4Nmx0RYIED0KyLhJltk+Fz7c0SWxCN
yOU/hesVjJY+lKufS5FksfYz9rVoS8kFs0oskhoEGTD5U7py0PbCS/qLMvbEivwcj0bBnZVyEYrp
4TP7MbIhyswBLs1X7wWZorKvbWj9YnMBNND4UQZ9cii97O8S1soU3rn8YVAOwwP734UbnhWWCS3f
6oj+gqNukwvAe5CjDIPkxIgUCIKBd3PXhOycpJxl9ITUJmA9X0XXhbdXDkzReU543hIcTjusg6hT
CHK8qjH3MvR1tgFj3vywhYV6qd26FNJKUQqes4+rDdZjWQG5SUFG23jlD7/g2xGIjl+ssofMDNUd
FnviRhYpNr/QHvfjFArDw87QCME9G6bql6U8rnIrPLbrYvnoXtRKJF6S/+n45DeDEpGbJ08jvtJh
x0kmKm/ZczbLfe6DD0QnsvasODHVoqHlGfVTYhP+9xoHAwUagmstbrwiZgXXYi45BTGe7WW+2iaq
I7udw8VDLm0U8OdedycaK02d/LJrn356Ir9c59Ks+U9D6+nIgqzFBHBzok/LrRBKBewHP86mJz4i
PS3w/F+H9nYUEzsTAWFHhIzsvS9hKknRnxdxurn9hpq0eR1pFB4e+KE6Vm16c2qEcS4EhAwzEKoG
tAm21cqqIbbDeA3yhi3+Rqrl29Z9V+EZIEOAumw3v3b/O8slT12GkeQbN2bgpUgl7e+oHOpTNE4n
bh10V30H0S5NlUxB3JywteI29m6HlZEzXJritw8g9zAIifXKBMVXy5Y31pbEczE895EdXB2o8T13
ajy0aD9naqPzeDx26OITrzwjm0sfaZ6OS3yOMO5dKq2UH4YWAF2zjH3P1jvqScVWs0EPMXj+x68X
4bquYylUdQ8LaKF/Yq1gm3ONA0jQBXw/9Ax6mUAl8CeRSp0POe6x7pNhGKx9MleT+x659WW53HCR
vZnFrUkFSieaREiiOChQD8g0qW7/QZ2Bsbp3PxFYMZYFHHm8vVuSYTdJhzVDIzKvcSt/TA289xBG
3FNl5oAl4q78PV5Slrmr+iL3+IcStT51jRtmY/LhTzdTKdEVTTNipBsO9brHpIqI9F+GGYL2rQsS
/h/+3Sj+lE2FRDLFDq+4tBhcpAE5m+d7CRfLebTGZcR2c5bjB5hxkFwNLd75AyMLdjub1/KnPno4
TqFRr7xsGnqSZ3UMQs3A1H9mEQBxHp1Smrc+s6VQyyTN28qh8V1i7sFAvUYu+0Fbonq+lbDfedAI
mUMFjwIidokjbl9IRrijLtDsKU8V3lFGb2csa+PWUq6TymvXp53P10hfW79zGEFD5hwI7pNpgumN
k/AOT3XhdpZpbuDW0DQ4MK27+tbODtiujnofRbX+PCVIgm2D7ipnGaiALOBzVzApCooLnEXj3iAs
PEOMDdiqK3P2/Q4ViAR5mYNV9Rzp9baE7Ay4WWiPpLBN8nw9tL2mdtmbTcxKs7qaWp8FnkPuCkiB
CgTCHmsqD1bI8ZxO1LufzfsjPi9Pvz34OjUHJuACSvbUO5/5SeCbUI57EbMxDWSDNsoxcZ0o6e8I
rRs8hIFQm1a1pQl4m33MitJKwOOC9t61fQ6dB9gFeXdc94TcSPbmsoJs45b4g4x+MSBxt07dCdYl
o4aEWRr+TwoORcS0KMZ1GeB3Jb1mLAcE8J8xZbkMVNoHRZzcIWbeX397+hADtIbVimqF4RlZoLAv
HmV2emfHerU5u1p6TTnbc6I1QVEsDUkZqPX51IiP9RWUmWBBL6OjjLYj5s+ijXE8u1B6YxaEItPm
FrXiAwrfArXn2Xe8Nxu6BMZwDud+zwoekpqADaqnCQ2ulBesCUx5CFP0oPgbv9UJWALyxtxWSSwQ
RyjVBdYwPCH9k0YOtKWOMbRUV3TqcP2zF67Xxz7mPZLDDzEboRrKA4xNp9ktXZ4vXDaZV07KeiYM
EEaEDdWEDos64OvAI593wwHg7tQgapy+B1C3ImRq9tUq2ZfKMdJbzyjyh8v5FvmxRnRGRB+1zn0X
IvTAVQoFQOyauhek96JNuImAI3kNVJv9O9gEN2Ii2heu8lXUI1x/ZbAQdvVRlCOexVkzrSTUVN6M
spW7EBvvY+NjDuPIE8EFG0l3OqWBPOnujgfi20sJtTHmBYKh3Vx0lP/G9BBIq2aI6cSc5kgTOUxs
21/MkUpXekmL9BZmsu3XqXfbZs+FXcCpz3iOez3yo0KTZaq2otcOU1ycdpYq9TyuoXYePMcNjxdf
gW2a0yk2zqWpCg22d37PnFk/Aae2qcxDchwi4BfeNSsiJRvMqtFInO9IF8mJqBX+xW8qhXlb383Q
iwyx0ppcCZDd3Pcszs0cwySa5FiCEerAO9nDm3HR+PJm1AKcMlZPSm8ykvv7jAVNGpaSVjp0dxJX
Tg6s1wwFjXWdS/xVhCDZyhD+AbxG++BAvZZEY2kzedoH4MIh8XhoGbbNPWFQQwXvDwLXDBv/V6jn
NuFOOYq6T38vnBhu8COh6Uor9ggly+JpcMW0M3aF2P9WcvALiBtXHtq+1cMzy9PlER2AdNIV5hAU
soE0t9WzXZC5xTES7ewFMU1QFWLehEgtn8DKQQrwG8q7HRR1ioW2uzw3z6SpH4IW8S1iuecUDEEK
ohDbp30GggSv4fTRB8JErjmmQh5JyUzR1IRqs+Q01VJFaMrWNLvC+wOg6S1w2+QLoS7FdjJromZG
h/k6ycrF5RTmtutrrpgKOM0BIGRpv8Czsv08NYJR77e7OO643b904povUxrroNDUo/yph75vsLEY
k48mGlDOxbIg/nlkcBI7hpLajZccNk497PcK74NqtZW5x/t47tAgZ5y81VI4Tno0fsTxCHaiR583
To4wC3QbljNeJoPsahXclOrsWQKekBYmlXMGfRtY5++VNZxfSQ8OXjk0PeKp9gWnqOsk9Y0HgdRH
AUpo3LDse+qvGluYrx3d5T/wb2Mvwk/CQjqD+bA+2LlXW9/lTx4nWlvguIdTeZHqccBfjF1rWpbk
Gj5IFCvF3QF3wnjpRMjNtiVFRCayETxytroSX7iXvhW2jiFMtTP5LbeNtS8YVXNo8Q8v1G7QVZOP
gUug88PvOKLUfeYvmXyONjIz6vyBtMoaRDtk+Yx2ZYoFajQnTWObXe31fszli7zKMPTcNhRX350i
eKeBBr1qDftbNh7DryG4BKBiK61qJVxQJF6gOlHQ9GrHFMRq2r7P7KATzn0Zi3eO5d/jvyfuOT5j
qCLCQmxEWhkPKyGvv0B21PgksVDWsdlE8ZauPC8aO8XeIVezO5I61TA9xXQV+y7VOZst/kvduv27
/xv0Wit2csKsBs+veUvxKhUCDRQOhBc24qEuBZadaeBkeazGjc4ybcZvaZ+dRZF163epuptIT/PL
5KBPRl0JdjJjCIzYeP3kvBQbHdczcKL0yQT6717dtoRefZxg/KFiCo12NL2/X7H9CWlMqqAdAWp9
pyuM4AV9H7NoTSqxA8IKMdUyQmFm/P0EGgzUJmtqGaF86EVIWH8BSGT1FPzOq6meVaEdErbecVv4
Xu/uZB75VqMcEL8GRDbDnomwAEJzIj/D/z3zgm5u7Cj0TpdjeHHFnWeb3Sic6XH4avpkXGrFIYss
crm0USIM4RvqjfK30K+ZfspTBTO5b2O5iC50fX2d4PDco6Io5zG1TVgi05ByVTwaaX5pN/8fgVlr
Icp/eKsnvYqMgNVCN8p/HhBa2PRPsN+bGxPZQ4zQYZn5fZcgeVSJOPxn/P1DMELo7lp+cGkrSC0/
E1c04NMff/QE9UAF4/4DUrSGcETqhlFuaVI3OM84nav5NTHKlcQbebiiqRC6nh6wrSUGE/y4vwhe
Ab5ae7FsMY8dMmjpSLtv4uYgD69DBizW9e3EQ2psJCyHE6OPejZrsCV7N+Y83Rj7TGV4GwXZLinq
C2trgSGpX+j8zBKjfxafud275ltP0zv6ULCkYUNKcUmg5BPCjclAT8pwv8lpnI1IK2zk3P3Ua5rW
arRP1s3bYE1WR9utGZwWRLC1aSgU6g+eQBhIvFJ0VIDvbEkJlXKWGQaHCrKQ6KDoi+6OeI8bLJAE
NTL9cW5n8XQK6ULxkhE+Ji8ja7spDRxxEkoZqhomzNWUEUEBA8vf/izXMcDSwy0nZhgGReGzkDsn
To2PHMVJrG7mYVb8jNV+UwrSxu19w6uIRNpIFS2zeTHr/j9EFnUW3ohoVqU7QBMx8AW6enfDnQyZ
vlEkZaGdwQX2onwj66bi2NZNRzv65pZmz4NH/XUNiscIs+ur+4VOwY4BLS8fjLZuTPH6AaYCHoyg
KwOHq3taXll/8Q7X9Fw5E8FOwLnCbLeRiDFgEcVqujlkAwcoaONe8MBJpl76kyzODz0+pmY1rEVo
mEOrk1EJHnNMYv97/n0lYbJeU11gN0xe9kUmPz9oalgG95mwRve/2D29akBiqIfbUwDCDVsurD72
sroxLcGpWzLbRZwbAUqCHF7lJiLagfvNGjdiIWX9o/jOJsatMtcUU/0V1DRbkgj69uckaOJznoQK
jLrVm34EAs2WoD83c1xAsHCXyIp5p/wb8Omma3B1/ezCmCQ2NVb4mG4CJNLJ2sPH16BiZggXItLQ
bInpJsyvQ/lUibqjLp8UiUoBVGPLk+TD6vXmn62nvAPaDxAeNrx2z1j6SDt4NJkhvXu97lhO81I1
m7f8gML6p/MgTcQN3OSnm21MToCkVjf3yr8sTwW38BCi+ISRlrHxODzorGH5/KYrLGTbj7cdJekr
suG+pTsHAM5fFUOCzxaPlcxiGXEcIn2dknmW/vQ1iqZB7Kv5opKWCML7Qmi/zCh09AEpec+LMOHu
jbNKW38MauGTRQDYfZ5gR5zA7/q84abdJ1IILhzFCHdk/uWza9635Qyukq/D+V+VecIhIquZWCYF
u8QSPwYf2OLU4rVmFc4dCyLEo5pjlH/bqPo5iovY0lBt3DYzyvZ//9vwAZ9hMYern9EZpSBtu7tG
UwXdc+sEEYaJ72huHpoYtl9N+i7wEFrzmd4T3b3DuitP7DKqApI6BgUlzK4UlfDigiiYcIEaiPFK
NMQGWGskEt7FyLbmJZW6x/8qVuF4hrLTY1oBg+HkYHUA14IJbofx/2Nq0B0R1nTC1w01oK9TQTgG
2qw4KDeJu5hNij1cdX0CHAsQyroIDTTJiFTbpmZaLXsIvxinljtVTZjJOZVXeQeH/63/KWlFjfhR
TS4HAf1s78ePloJOsGO/TwfpVdNz1sbs3x7EIno4PTVs32xTJTbsdfHaBlt9H4Sc3mIHZVJmjHad
nR8EY//gCfB0FWAK1WwxuvPkFRY0FmZF84gOWlq6yQmfHOwr1HlOURLN1YDmwQmUyow6sQb5Nd6M
euNOuhq5tba3Zd/IzjtwfuVEIskqvYZyfv8BFGLzID6US8sFarvPbQ1TsJhYJsu/yl078EIdOKwW
atBXIopITqB3UFAUwe/R6wV5acUDeVSyNVxZPXzI1X5MCB6VyBkoc/uIj09jzMPW3jeg5HW/A0YP
ndxJiplSpSzkCYDV8GVtUXkR1qG8puTTNTwjJ2lhziDNAb5i9Yx2rmthp/A1LklyaNEraYswMytg
c/b6I2OSBlcTcpwrWxw4QHwUNNJ8IhktA6nbKbUBb0P49TC9HOZQLp2c96lbpytX1YZHzEL3Knjz
INsqZ7LjFj5u6d894The4c6j7UAzQyF4Y9IcOVNbVYP8kBqFidkUKQW/IX3AJsILODIvVZT9Mtvz
0ZVT+Jl5BTqvRJmVJp7+UWXvB7mR6R2rf+qBXrzR/XEf4MC9/7mSbN6BuBnYXK7a8EMXzWOPntQC
tJXLUw0Fv2LYPfEVAg1b46cb4oTJOIRQ7C5YImfRuqo0S4tCQxlxuo3smL5r2SgqOTxN2asXHSsI
xAFUzvavtdZ8r72kyIWYuHkHt4oqjFWDEjqudnxUdZevTMjFI3Nr0s6cVP6Z1LJT2Rld+YcSzimO
4ZV0QWFc7+XgXWRd2DoOLDu6JHuTwzYRmGGsHqT3G5vb+59glEbyVos38wXHgERt1eH5kFiAO2xO
hmzZbuDPY16NcoTzamwDehJwmjGoK6M1VgMVjbOXM6oCvC57vCB6zdsIvRFcFwzCgLGjIfPnN5Z0
f87Eh9F7N/gec6Va7832vL5+toIKDRQsBw2X84ITJfmYMPxukZR5azHZ9ypFNRkxTpFJG+orS3hu
BQE9HufpTdLERXNsPGoOmzdhNwobHqTOxgd69N43cS4gP+sVlzCOsEUoMpnc14ALqwCMWq/btNyo
7MAE+6aFRsaa04Bzx7GsF6f1HnuhHPJ60vdpGgzD6J9f0l3zv+aQT1k8G1jMJebfDHvFAa9jMdD5
dO1QlxL3GzYiyBzfRzTQCsZ7pSK48y+Nw8v8d1RLfWfFeQgjsr+5YvHImztjdb0rW9pqctL3ZyGJ
Hwv/AJxdA+n1movMH4oltR6cy3nSXjn/e9yvprGXEUXn/9QN+smwMy3dUNeM7pYW6hleJBGcQB9V
sWEKJhWzB6M33mDZIe2mJ8uQFbFJTfg8J68zqxlM6NwwYGyTnD6bySzl1X8W1cHv5wrnrfkmrTzv
UAefofjAYNIm7Cr1uLKIcCWKdwH/bipzUKRZ3TmFwHklESEtqs+8ly/hgldEbXrTgpK0CiojieyE
65eqlb4lu5M+W4bm5BYDPRHmLF27zRld9RldDg7KHPDsr3/+FtVm1EedIhmHvqsWIicU13YqSr/S
ZoEf8ZEit4aX6i5mflQUc+Hy0ks1liwN/geFHlXHGXBtp5GxPKfY8eFIDhOLO5Gn6NMVDPfb79mx
oKi1sEEI6TJJJsrA8kkfd77HfdQGTwL4I5KqhmXdSx1RDFRDgsa3ShTh3TyMV4EVJNQLZCwEy0Jm
4N1PCsxV3kxTKYvyfaSIdViODkaxYXWI964OXdYlMIFlUL3rhWAtXr9+AG0I5Zew1dZe2dKn5qf8
2SBCGSHJKmZnZpQcwxVW4+HYgYMzcVMJqJK070Bq3+sibCNg56wxC4zRAGRJWE9mQRXLc0C0Hz4w
rCyqcgVn4MzJ5SgUuQ0dhvgIruvL4ScbuuMY77UX70PhBWHOVhWSEEMa/5UUo0mH2z07/ppT0zUK
+TqaPR7ZVXCe4bFM9HsmvCdwkyDNgUn8Z5dX3rB72EI7/n2kqn6eYDxnGc7rSKcMrWWTKRrtuB0s
4Q2ma0nW+XonHaaeQMmVRZc52dr+D2c8BpZxWNdLcv8bFE8kN+Au8K/fdTpPI1QSsLEV/o3+TTGQ
EZm0iJEFXWJZEvpBWhSnhIAGX6FOa6qlGRrf38824z9N2fAoGTrRqB9ebAws18p45b5zzwr9khhk
WwH+o2Z90evKYhxoe1fcwZMClLEJ5AKa+Bca9vBMAT4GNskBfmfS/HKQespHZiukHAslM84FIhgi
ZcFOtFVPilx950v/pex9zZGIieokR0ea/5EHmUIfvN/tIgo+0uxYS9v+zWcIY1/aGOvT/1NT9/x0
m1NxayoAukDdyj1SxR9JqsrIk0TYR4E+ObrJnZqluvDRkjPrUz6Cebasp5hWRlO1Iq4PcN6EWMiL
RpAgy4Tzczt9Q8vypJR0R9ywXKJ6llN5XVH9VNvULhf9fZaOU/5DmLOKwbmZak9+Lj/VVv+fQu6a
fNn5+eOb7LF/CJuFX5N20htEbBETVcEhu+9Ou41Jw1VN/hXT14CzfiDk/hNHUyxdEWmn+j1zhw87
TCBko74EKH1SPHg1sy1YHFw1O9iffiXhsKTG8bDqv12iT6WZ6RyvOylBMfAobonY1jVZw51y+FLP
YvJP7rdryiL3KLXbGZYroydDouq9+Yr9Wu/OOB/r+wAM+40WL1O/a5Cd7arQ3YZB3e1hgwVxWxY4
7p2yN6CtUnNs+WvnKpVkd6ludxFI8PgD0dCM+BCXkVvp9nydDflVi3qTG1eWzaOeVNzODIVpIYnS
4e6I1lzqobNMpPH+NpBwFsigHfL8BH7OKoLaG7LaESMBm+7S2lUO304uha6TU7EKX+9PEqwI+OXZ
xsLnaiAuJ10gVuR0MHrf22m0kxc4+qRFdNxxGoy4JvYKI01Uh9yui4M1oKnrzidIb4/R7aHHIKEu
NniUtvP3ZF5C9VoFaQOi1Hb+jqnU6ccfExPdVicUOJp74q2g7aB0CmE1s7MRq7ozTFOzWT+41t8l
K0nBkYZjknSrHd+6w6VLpXmMh9UQNJIpArSgqxKB9qqt3tNnNtFBzeWP7eHz37MSBp5bOrlHSk9n
XaGp6LiRxeX5g7Pk9E3NGPLBQzdeHBz/GjCzW9jb5bYO3Brsq+a59f1SWCjrfuHQGfkYG4BnYTw8
tFmvgWHXkRGmbXNFtFzZbyfU50Ey0bmDdNqV5ayPvItPrXTRk/Ppg3w+CcAY06UqimaPOihAtZbh
QEj2TXEdj1ykunHMN5AuiToKootnN1mj61YFR0CxoV6DJoPHUjAhhccmN9dJx4+PnvcKAMC2wzQQ
dEByQw5gmls9ROWsgB4Bf2PM0/gxm0TN9ncwwuZ6jF4lSsS0gThteN9ybSh8/XpLFXBQ8CbFPAmo
YxTFtE/QPPQ3XR5iXCJ7S7k4LvWiLQ0l3LMPrZfwYgiRIQHEKKa8qgqVVHE00RkPkbTu9rdPpsvZ
aqVxY2UjVRjpRx34AjUMRQH09ILmAeuSddgnqDofYrP0RjHIjiJkXGCNhPHyeqK6FuwF/mC9iWI3
ZQtReNk77szG0fQm5DbEDwJXaiG9ZZJ05/XBrzzx3mQdmbsA1MA2pFm/XEVLmUpSGV44wkqHWx8B
lyCl66cl60ONGuyagkpZIhMWFCRDR0K1EIlyLFjbMXo5KFg1UrW/mfArfLGFMr3f4KD3p6jAlMmy
W1g1Yzfg01oykJZiD2UzdF+mWUhgL5y12rwNpKTF3obAqjez1OPMFpYr/Z69AmfJoyHZEYME3DmI
d4tO9ti4YQnQ1eK+5RdxyfEa3nhn/a9X4sm8QsxkoFLHABBNeZttQkMB1w/BiwpUGurRzqUSlKSD
pVIWJ1jW6J+wQHAgeO+Tup12/4ORdpUsb6n1nJQ17itV3T+BC5l7FWUKjecK0jsXaRWJL90MUjkM
d3UCSnlHvy1MoBB8LQha6+OSeYcJzSFtFTyTZsSOzqydls8fvuzluIxlljIF8bM/ffDz7qbhwxHy
tqHr2/v7j4MPt5kVJgLdl7INnNzJ3EXH1ABrklerL3jSWmAnbvGlR5Vf1pmqOvh6r0MpPk1JUijP
L3lz27fRinT/6kguXqoa4IM+kVFIVw2DzpBtZ75yGHOn9qKiqgpK8R+CPQnHyV0lfR3LR0CraJk/
ayr5MILufiwZnD5gT+6B3n8iXrPnUyf9h3q/Pxi9z9UIzhl8U49NcEq2yRpzXSex7l0nnXwpJcQZ
K3tBN7xa7LFR8pVARQhlfU4XDybAX+uScNLN6M26nrMPQsj8NxJNmzv0ETVLW6MBJmlvKWdJJkPq
SMJa0Jxor9bdFt3GtGaMgRoO7mUuWhhcy+W1H++iU/YQ3JxDYYQGYttBUZGRdo7Lu+efkzwzKAQ6
TEerVtoE65TYjRbwMVAAzoz4fsbPKVcelAMk2tglcuYQ3cKuN4ozdAqidamHkWcUacJpsywQ3tfS
EgogzIf+5lKQbjFZPVh4Gr+aszU7p1n9fpALcJYGRLj/cCi8CQcRPKoCzlot2bIe18rv7AUTBe++
imARMQQ5LQ7CYFQBkqp4K1i9eEAxOoSCeD260USuul90NP/w0XzGQMYNYQZwRRF61HImLj/w/fgb
JUCHQMVXtu2y6GTN3u6hGqfTpxFOC3Jrg27fP+2egG1VTcrDF14W17Q/nzQRSt1rJ1xldkWgU2CO
1S1WyaODZRRxiBSI3KPDt+256tA0SPNL5tyOZAsM/HsRCKP0ByCr9Al4dTR8QaNTYJYh4hbzNcXz
sHVlo5RSI/PABQJI/AEgYNZLDRt027UiHDZ0A5WYHT/49u1AJ+49Q/XIamc8B/LCi/CxEBLNxcsl
Dzml7U8dEZTu0K/LSioGBlt2RMXaMKxCt8VM8E6NlMap7ZIqSfucB8R3JUy02UdU2O+Tsvby0nA2
sWPFMGASh9Lg54ExMinSx89Pc9vMJhkDPGsc8MptSKwuSoSM5gKxCliBrktCq4CiP9eOO7y8J2wQ
SUKQ03TdVa4VPQQfU6HgbS81GWtayMcw27kagGKwTEfARn0GDDxQjQNxE/gtzFBpXV/DEAfEoikc
xY7k8hZ2di8fAWziKcpbN5roDBcgXE2VkhNx39Lv1Vpb3qDt7AhRyxcjFIu5xbQYjicFq8I/Egom
MmY7BYa2opT0foec9EcuMf5Qcgc8XxOHf297CHsuPvIKBXHCX/CGKcJbuehCFRz0eYf7evvvbpzi
v/L8U6vax30O0Lua0Gqrjm6fmt1OllMoznsIFwrVSaKOSGcf0lF+HDUOY1WXDHGQkFeZknoKzqHZ
yNIz7YbNL+09oblcu+U8+04Xy2WgQvEhLklX5A7/DD3jIc9Ei1g4IA3gtTIsvjB4vxHdscp6dH9Y
96dWgXdOibMwr566TpfnCajiA3sBZjqULDML5mAaVk58w7HiRSV498lWXiRYuG48tw5dk1uNk27V
j+ODixr1OtHWFWAT196uTRtbyqwC221ne6HWEgmSeAQrVKVxbkJLt4EKSGJR1OfsCvALI9AaMuLI
dHTjltcqZbjPx5+1cEvu4RIokc5sJchQ6fByHSg7XlI0WMfL3zIU0skHS9PIHlBsC1PWxEunMLfF
emR5mz8GI4Cvkpeco6OeDMfzl7mhdXphFjCJ87W/5PFPlwhgOBinaMiOMI75pt0K7Li271/6/8bC
lBunRKU3GRjgInmNRAoZJByQb2R9M8y5n9xhXzbYLlKdoEgCEvCyzojKxXmYVt2xkBXpbE/Jq6qC
YkfrjJd4ANt0JvwlkjSDu8aixFs1FdY7XBa3NYMlz6J8eVyGIOBOMu6YMWA6sXfZQMowYv82UgS3
IbiZAR85MZchb8zYLl+kqd+UZcYXjLHScW4jskb7Zx1n13aGpT0b0LKn0MTdx4BPM1/Donu1/x9K
7Rmrhcbp+JwjiVrB5yzBbYr9N6wo2TzhsPFU+1M+7BcL6+HIAWzvCfxPNXtr17FXlEfRqDqzB/Dg
L3hT4sBXGuYin2OngNwkEgtTF+Ki5fgD8HL/YAfhJh9gXWQRCcq4D/gz/sI9GO11H7Qe0OJv2iO3
qcz+rJ9AwXdkgGdV5MMUbmBm8flm1xyUYaeswFw7vrPFy/qezCj7Bm5mCt/rnQ7n+1pW5WwJeauv
Md9B7aaWCKHlQQDpc2DOGYSgXt7nLqiZND7HUINFmalgjQWBT6+ag5c+pcFTPUrtL75zcYI7LhVq
pTtapXkfSqHVuSTNXdyKURzfRt/HuYOvBFO02URRQ8iejD7u90IkUE+vmrzarsdhVZvAKzNaiu2l
LWtNVMFMxlY4OApRU/w+zgSDGYdTrk01BLkPlcAkAGNFDKcbXTA27Ob93V9Wk3pUfdwZNUwc/dYe
2EMah6JyITyFpL6XIEBe3BDKJYeaOU63F4tk+aDirrohzcA4+fzENJblAiV099XRi19FOqqaw5GG
DlHVEOHmmWOrXCYw8CXdTKpt58Hyf3BBe02IXob7JBWYJqaRF57+qS+zqDJznL26vLZtoBYu7cge
HVwvGT4OMDvXvoHFJGKzONYo+45gp5I+eBp7cujehFZCMg/XoDxbabiUCkUvmFkaCkXgR6VVnyI+
GfFA48UJNQ1ENSWTx83GzY9zP67bQMgR8F/+QRr0rOWg/K3vvakpo4LZnseJqTiIzhpVa4UfR733
fi8oXCyii4toxVqMI514DeUlf6MsxeCDTC5uiIn2MRz++oxfZbPiQ+Dhwfnx6RvOM1Y7SzPSZ/18
vS5atyf/imuDudBaVNX2vd1kTlt3kRnimUJcH65Fb1jptqQIaFkm1KXOKfpb41OF8Dbzv4XTEBrt
I/bPYxjyroqqPY67tHCnuYaax96Qmg09aSiulOyaD3T8M/nCQWqsnTPFxKrZx8Bt0ae27brv6pBj
4D41mBcnoJD9/w2D5QcZTUpYT1giW0I1atQcxLCQSsAXj9X4r5Tl+zQnXjqF/QPU+f+LRKVu5tW8
0hDZ2tjIqPRs47twOlh73Xp59g344DMvg2xrzlgOYhlczD9FhgG7TR0srU2urbhdsEdJMUZiP2Ej
DH2cTklJ35T86mSPldyaPWrgkihxO98Ma9fnv9NnZC1upCw+Yt7HXEMmWNTPqmWaC8hScKO1p5Mx
a9Ad+9BA8gSfWwIGJsqJ+4lf8MFUmKS7svQ/qWozWmO7CkqqA3FuvQ4xByEQPLjSUvkPLY6RBumA
TC8zM5k7TKT7uaavpycXScrQDkHHSKkdHNkwcviyJ4RbANiaMdYRjE2tdjs1o1XtLslhtexRGn27
w6jg2n412Scyiu8mMTUvkJf2RQyxAmrYRcRkRgapQAK5itESLj1dpSc+kS+t+StLpv5Fn32PJf7c
W2Rr2sLNmrfXPJuAdMJt0JVg+N++m+S04ePsOzQAzX7dRcRAIPlgs+jmBU4pH7xJgxCUQi0oIxjy
Li45q9iYDnSU8rc/aFxG+wzGsWRUm1gpdMibXv8PENpFtMPbmRgGXfCa+ctV+WVEcn+i+s/0E29A
Wg6TW1BkRV30o8bhCBQi4DoOb/4bdWs5d41z0hkmYzSRxXF3FNCmF/p54b4k/ka0NuVivlQRsn8t
3rlnFq9b0Sc/JffJYMy1ifgNU2WHMhVJqJWu+7vHtx4886DBO1rLUid5SCh7JGggzgzAEqmWy59y
Rb8H5p3zc+oZG7UbVX5p5Gq0pu5+RpZJ8O5O102QPRahFN0mQ8ZL0I4gsR5WH6Xdho7Ne5+TaNkX
Gw6SYFftgA6EGPiHhknoZY2KkIPVyCTlAPOP0vUNgI16THy94mJgk+cN+ro+7dSgIH9okV22EOCa
BdIkUCDZO7aQBLrsJoYFvk/fP0mKmuluxrRmJ8aGFtlmLBA75fVsaDfPpQPDRQGpnVk3SXyRXcnB
4wXxM/AgK8+fWu1C1lKelRaFx+rvIR7OAsnOy0eUjqPlk5CBHHnq+s2xE3GhDJd5tvJ7gl+dI/YS
L704IFL7DCiHbIHQfhablicW0rqHJpMDgwl21RoIxKKfb83QzRXfbZTcdXaljG9NQy21wr2ojhaT
fNMg9gzBQUqPMqnXjUGHmRRuF91Kse7HGjjVBTx5H8dJkKonhlBGdKjm6bGNM7ybLiM7oC1qjd5t
59z56sNtGB4yxKBYy2ZUgK9UttBGtdKXV61cfY1Edi2CTqU6mwo7BKXsd/1fmW6eTkxOQJKapwwf
GU2ZXwLBb5dQIV/yhVCSLJPZ7KvFXP9uu+AYcqv0ACGgKbZ8/I5BS1iaf/G16XL71j/NF+2OSnHw
GefJG3MPwaCJKTKLZrkstowYnN+RCJjfVb8pkWAi12pisWKebatHBzsf60THb6uaDCZW3n43AjSL
qsi8dmpCJuCCvN9TR8xzjCmuR9IbjUR0V9tBFgEu3UfCgBh0nTyC51wL0eEkjKjuOb4TQonnqzEd
G0Ozr4Aq6c17X2WElkHSzm+qdVTObdVtxvNx8bJMlpekiAlM89/RGS6eC50SYDQ2Ui16iIfoZoxy
o+cu8IlgE4S0ly4/tR6NAYoxErsQVXGG18OxD2QasWR5v/Wtme9TlMmj7JEIpkUpGeKkiMVonVqL
HVI0k9xXqisDtioT52eDHW71jQOrq2/8ArdBaznxthzSXRJd9aHH+7tulTurV+kqAUHrYHBqS3XS
7P6/5hrRBaoJ94mi4Z1ZhhkjOdvlqPxuXMAdulCxY0XBuCA7wI+3LxpU66x+Aw4ksFiAdIbV4BjA
leBf76rZ/5JGU6IKIdJnm+Z+L4VhkJiSwBS9gF7Pu0OCzXg/Hvib+hZReCJ+BP1ha0J/Ayge9b3+
Fo1zTT2Ccowg9UnDoBpFiYplpAg69+BJq8PWNbuJ4dDV/2DvS1+GVS+l85pNFcH4/bEPefkObZxc
2qBG0eec8kHa4K9uUT9/tf7MMwS/MBB55mNfebhXf/Gg/Yvi9PeuRv29HiA7WxNPaxt+GiGT0Evo
6qXhC3b9W0wBTX7ei2LaHTO2cdQPG2K+8Lzq+2lnY5dkeB57L+A+bMNYicTzkqSi2c2zXqYCxQVq
+Ue0sSzzTxqLL/KFrjd6M4uLGzT+TtCeG9bflm4rMhzWUfzd6XEIhwS66dKeOtc9FAEFlMSOEUBT
S2S4ZGAixbmatsKSBqZv7agSyvnWHhmoGun0wrDkCnPLqv7mdx0jQAoia5ifb7K/x1Pu7Q/ZH7cw
trx5raAG8QvF8ConHBfyYjF/W25J6EMVJDnRGSqAPiuT1Am2fBogvvbvFdqKkppbDjtoQGn+8zpH
uYpxIsFJQgOuJ4kS+F9aHAUxG3UyuCVKDyCXpYA/vvkMGeYRTzepcfb+FUY9A9jFWzfr+BGBzLKe
aMKpSt5qDFOdOUb6Mj+jL1lr0WKJMrelfAZgjzrTsWpbmym9wEoaypJRAKNjyvxcBcso67nYP8ZW
hBMa6/KGrQlMOM1oXDtUrcIGT00wShpVrzCCD22HGaOP5Oy2DZReaDYk/x+ztbrgzD3wwW0LUxFx
7dWaklJPWwzxvci1mPQrCWSiQUC8BlH0Y8m85gSyfponGtjbOuYW48cPF+2JSQi2cvsUZLOXtyGZ
uVaG6dNc8vtPh6iN9LoLEhqTb5HnB5FuSBkA0LnCu9fnm0TeuPhFru4Dmx7m1PeI3nl1PBUn5310
2EtGaymidqUnmXLtxeocWI0Xz+7FOwWmVLL4RTVDAcuy6x5Vx5lWM/Wf0Dz2cMcSmHlK75IeRPN5
bLpLWqyYbyUpfeWnqJX6fmocGIPgHrn/uP+sIyf8TpQ8KVS6+/iPHc1ZOjdpfi6jiLWBUNKHGY7g
pUWQzjt6gng4NU3aMmqVa9Rm4fs6Nq8tqWpwTHxqbKpI8owKIUkQqSpdqhhzegFnrQuceY+uxL3E
g0IHlMAmZUyEO/9jNIXBVjVtE3UI/02UW9GQpQX0wrAoY0gHZUqaDW6ua2/G5Kb7At3qWKfQiuun
c/DPofHp/C+sHkZMEdyFyxxai0ikj8aCsmbFwcgX8o9GjkiFsnUjHF5oppcJJHsy9ey+dvcIscoP
8kai5ORT3vRc3XV70Rq4NXT7k48xvvCEW1mm9BP9BWN11eRuZkHYZX0kdGBmyqIzsmMmSyhrmk5y
pSgUsAdahzZ9/HrY90RQjbJJKvHCwaJVIruEffDEU2BD7EPKxp95WrMRVqVG4tyaTQnisq7D7Jql
pNCbw66GD++bCb1fY+db/reBADGlnU4RdOKP9KWsbRo+SNrordZTWLl686p5kKljDpKq9SeY2sTB
O/9SNKQi//3Z3Vl9I6cnoD6dJjiaoBgKCWyurApz3n9JANGIJ9mkHLxUKxHm8ztPHfddhP1iMaVk
8dY0/C4pbr7cSUKiU3rVokR/E6X+wLIN5VVBxzvM40C2tEv736nh/CS/P6zE5Y5GAycUKYWujEgA
PzdByyXl9KFiYSd5FvJD1vHsHRKpZctYrd86RregLJBFKRIn4rX9g2OfDCdkkerKDOXjViWepIVt
DmC6KA3rI/f7qy5zgFUGvF3zWz3T31kUzXorNlLq6viyfb1ubvmO6kyPk0GGkoGE/YZnrJ9YeuHf
1NEUYMviDppn6jxzMGh0Pj8RswQHC2LC+1U8W1bhhDjuOmD11jhZvlNn2roTr6wA01KRYXh6j+2y
HYPkyZT4GA4zxroSi/egNyTpYUSwS/UsuSzLkQ9yXpiIAsxxqs0KlH+Epgr+pAXJo5x6jCkSk4RX
HoWJqc0JGFM33gMOorvorXVI6MTGcxFrgevsm6E/QCni/MZZv6VyrSuD8hSFObYY5btvmdoR8isj
1PANFTLa+iTZLdqn/tHsb/L8XWlondmaCUBo7G6UK5K39H3D1HOvKAcu/KcbrgvBWUmcz3xOPJtw
EnSD9G/vlAg9CRi56YXjWdKGVXaXSPMsevC5e88k4oik5PPfFK5U9qpcFc3AM4YZHRZpxUm9ELqE
pbJszel10/lQDNkCg1z9bUVWDHInu9RTFyM9Jd/1RypthkdQXMSUrUwLFCm/lmZZQY76utPmbVqP
3e5X9aaGpefQPHq4d97W4hoMMijSqZZ8MAo0kYVeacAiKFedPBiV35yFIRCY9LJoKEhYnH4hv2eQ
AuZNiTRedVcyASE8/pfUm3kgGr6RuxrKmDEO6Zdk5251wBPiYA2PdZrkbnHmkQpXB2vEJfSk7fCU
dkxX0we+ZrVWdeACJ0elMLzg4LUJ6u+d6KaOLXMImVOOUvjD9tAfxV2Uh4EfTDHbh0GZI0bh7v6Q
1fWGoBj39OSg8B5js5xXUTPeZq7eksuJ7HuJFlY7LT7XCaKM/kisyj61ZWjI0vCaNPq0k3umkrR0
KZbrI/C5wrNNO12EazbKd8TetBPMngFY4zGGgaZKx13U0utYlpLXjnPc5BgHZ73+bq7W2Jtg7QiA
wzS0fvIwwCIeu79uJI1bXksXP11nbbNdSc8aa44udVSIiiGKIK/JeBt5gGfuYQ3UhgzEIU+TOeLk
v1lX/AellSir0o9d4MrPDPcyWe0jUgjI5V6ynSjczrep6usXXlx4hTHhfN2LKy3d2EXyoGpgNfS+
+srGcVehfjjYaLzveee4xiV1xRrGebyRtyQ37ahqW4+qst3FepX5raUp8//SFDf5IJkfzwR7H+D3
3ZsJEfvIE0uLk+sgHZuQmzJKOqzpjM4uH2r9UoNwYvpLPqr9USr6IjfyXQmZwRxMTAD+I+T3vpZW
tGTua4kvPrNu1kz92XuHu1Np10xweCMm9yPCajOU6mhylgduyyDvhURn+LXNLWOYjWexFG2AEgRG
nw9smhBbqnWypIRqHmrat1K073YIodEU/oHx2nWf/71mRkAtjS86y/JsSJJ7+nMBTN9gr/m5oMwV
2ypdirMIOKR4jl/+JGD9I9q/0pmyB67Ouf0FIohuwa0B/VKtG2dZp0CYjKuCy/N/z6HzYOFnXhNX
vPNik/3W9Z2XTQKW0iXYv/KtpOPqnyX75epGUgJoEu4+wrDHsagkmXWDO4GTMGHFeezpmgns8IOd
xzeFzXI9PHctCYusc4hDiBUXU3LUAKeTtSr8b5EZ3EW14GWjUMjDhXL/YBhfd8YtxdVOQh7kzbZL
o3Z8ccpPMfPTrUd3TiPzuWEkP7mOGHB29xyA2H2wrrXH2LTRv0OWYcJ3pHHX3pnJZR+7EvInHv5Y
ockcVfA3wVkAmol9hMz3VNC3bYnTnyeuAKNF3uSXoK04hiC1sXy+bWm+n/7iObv/B1bacYgLs2b2
YNWihowQPezGwiksgH0L26YRnfRT3eeF2M2bKShliiFK+Iqa/QhffV2uhN31kDYe3wP6m3TLnrjE
swMcAzL06BteHeHbJ6fz285YVWKDDO9tkjXY3YjVI+vRe015FUjtdW97MtUnw+bya+P9IIYpwPaZ
PyJU+9H17ODAdpS554qAw28IWCzper93Wyp/sgvR7A+sH4MM7Wz/S+z2E1rJA3y/Ci6UaJ/AurCD
Gk2lQ87VzA0tbw7r9PutBvpqeJRkJybrMCATQ3Q7U4JzyvuinRFHhmwfC8aeXQto6U3lkU1kgdcb
dOEUPRUOcQ/lmGhn6AkkAE9whsH7XFfZ9p2e9FuBMBVcZuQFvRMh77TZF5y0eraoQx6Ujm2ZYPIq
ImgWH49RFNAY3pvLD6y5HlVEHGnlHZg9xSELybBA/MhjLrY0/UCApFAFfyus3XcdGArbAq5ycLVr
6LPQMVbiIbFo3fp8Vj792jX0/Y15U5J5b3n/i2oTp8sfCGKhNoNwXca/D8cgxG7/h2q0SA860Vkp
pDiNEYTgbbLhDk4y8wWjmEFeP4YnlQr6gehNBGR3cj9YJ7ltQOGwXVjnTMpo9+qsXEAZCw1Uysg3
9OOCQUJF1cWuv+A7TM3bM1THtyhD3ik9CpZ2eTdpQq/mnHQxNlkufBXj36qH3lXhxctyEHFJbHzJ
nHUJli97IR95ZbQaG4LF3e2YIKXcKBXMAgWmuXt7X8Vo0s/FEkm+wa/K5tvQ+s8B2JuurGiRcGdj
/USOTlVTbSCFtvkO7UvMzQ0qjXgDULrzKxspuYzkBT9DmFE13Todqc8oF61AoAmnXy9T/3qC6I5O
TKDZtMh77dmyqjIjAbx2QdLW49c22z0ZHjR9I1fSxkN3RSVWgzuc1yRCTJV/LfZpRkP6RTDYgCck
mQJ3lsv9Fd0Jb5We3sqwTLkJ5QP79uoJfBUW7wkrXsYP77ZWKBRjNr7jGzF2KpXO+0ydQxV0hwUR
qJz+MJbKuGx6wBdGLNtu+Nd1txOSdhXbzgp0paKgnDXxGn34aoTl/gA99foMe0Q/zrcKvgAnWgsB
cuRHLG5YPLyR26pDTQoE/UC8YVaSXgk2e0CRWUm0a4Tef/aQ+p/IrbUZawocyUqYZtTvyDEKxQKT
GODPngPIs6kxEmd6cucu1+PGy6iZs8583FXjp2V0/nyKA28scQo+mASu8xbWqg/S2vRLZm5kd6oP
sXYQt86JIlhr0+f7qe0VrzcbiOEbo1aEoLdodZ4QNBiJdmtN2aoXYYfeOj0Xdf/VAZFWuam3/4CM
wv9sh4NxNMlxXi1hUj8RUQkznB6m3h/Y8Lsqib05zYMSbOjNLQC9zI2RkEaFMoENDb2Vl291qdZq
2YrgYc1m/ZTUr+NzOB8XYLSvAKFkCI9AVmvQlLmOi1QTc7+jrVtV4zT9kRhbq4KgGu6j5Uay9NgH
GbRnxJ17zlelnEf8bGnE8Y/jsB2KlR5UX3iQmV/Bx9t2YlY0I1+jubK/ODip8vguGr/hqvUaOFL2
eQ+owJZYXAIHqpMur4rQ/x36Jtce7HBNNKlygNKFN2Ohq+bgWG08Kn08yCfzT9cO/RvqrrextW98
ay3HcwRyIgIHUgUjcXkg5qFZFclLQeDDwxstAFZ9SYcDIM5WMDJ/rWdo/Hz4EBQYKXOxz8hA+1Ij
HC/IpUW1i7HPWSceayhkeh8rKB41kdxqA1rIYDUwdnBRnVpVjZa5t56EMXGyQow/yCrQ9KlLiibV
a6E1UisoAgOf7AOddgjrRt0GSnLL5UG54pz6QSKZ2aSnmW2KBG4170be8SfqJEWcpkN1x9IwBRUU
E/F9WJEqdJrw8SDZQsLxsjliLRory4f50L09EKcrwakEUDFOXH0CFYlDhDQqFp2V/DRvUdcrGiji
eiVvWZsGZbnK5rhVib92rodap9wCZkZTRDmLAq7gg3BlcUSqiqMHmyza8UqGUqYw01lrRG4mgr4P
nRuNk2N+MUnaFon6AnAQBS+UvmARmwvlP/rtNRaw079AHqzc97hTkpBEgvlsAsAYukYi385XAw7c
lKpTjjjPXwTalb/kMqaP/vnl02CqbpbFtlB+gYaFsyR2/h1vVaLilyP6QCGp8uc3arKk32DZ98Yi
RYmsfJ+5NhD8qbB5zstVhgcpyfu3vyQtJJlUBcltSG4Z38LuVSsuUkOzCQFsmZv/xKuDy5IJvg3V
R3Rdb75xPzFVKpX8cf0liP2QlP/LbIdBBQ0bkCLE4ppry1K0BV8oqipKpzV6ZG/1IJNEZFpdFnj1
7rFZU+Y5YJGSSSuaSKQ8eyznLVvYxB2issz9+As/Bh1PmUcxMQEoujQvosIzs/iXlKR48fgOPKoa
hVUJGPrjeLKNnvabcGcuUJayCNh5zirKwpug/R0VlXIJJVWIJgFfV4H6ciAuvBo6EhfGnjqSt49L
zC0ylhIYhjEOCyJebuisATgPj3En7wKn5pw14gY3K56jXKnf06tFn/49mlaAJ14r99rGnZEgm758
xQc6IQofqbCiH0aOZ9+fMstlRL/69zogZoH6neQyF9oPrkXkGH7RY14PunpDpkrA9P5mYhFlzjnA
CNnuvNBzTxX+kXVtnWDI+FQR5AeLJCdzkyjLkRUxoD+KnmPQi9l9UPWthgfn5Z8r8FOmamfC4Z4E
3g5V0G6kFaZ+uPei2GIoagDiuxM4hMTi4gIvp1ZZVV34Js3R6rtt4IbNJ6XqepnewFv3XItSXKdK
GxAjg1tJ5ABrkTqZgNhJkKZeZ6tmKutaUOQojBcPffoHgDGkrrdezVg7Ok7UxGblakKv1E7S1Shx
qQG8i07XtIW1N2kHgZBukoZPgbDeb/uc4dSjUKseAW/WsyToFjINdshCv7TxVbml3RPo5CUPmTKB
BilvjPfrjKDbpIMWzGGXcu/WrXS/A8+B41TEEk1kh0TfHD6TNy3NiuXKga36XIyxFPcRGVSFdsR8
mOYYTM6WGtzyCXQSwRK2+g4RXm5HyDgyo/tujaaEj1B5XBb9WzlTcOmY8v9rSmmeWFY4RCgWgsCA
DkYuRsA88fF5y0buxMeJTBf3GlcXImMZse/sD7Ot/CQbvRVh07xxQ8Fu5Kg0kzvD/2Juw/IZt4Jp
IlqVc5CZnZXvUvnCDLtYUkAPFxcQSwyU9PTddoiPL5Co9dpMADzohi9+K9p8Dqf5u5C90EYg0JB/
24M+CdxJF4Si+obbsjz/HpIJOOHxZbELr9oXFdnmIymFSz9FWcDT1umibeP2ulGTHdW2WIIUzo7I
wYib6I4jUno6eQW1X3vtGjGCwG9AVhR3+SGfl/gFhCrj3LpGmylOl7AXtibNpVNILD78PGvM1FFE
Qq4G3PBlEDlodhvVax1iG5poVlDVw1k+WVfaXjQ55sfdG6LVvgq+mBGuaqP5vpXItJPO/4+xu4Ae
f5mzZctxkeBfiuP2Kt479tBKw6sk0AQXWtOj0raifx9mVO65ohoxqZtCRIaOVREdtEIf4Snh5Xs2
vuVtoOvKE3vReMeTI97623RfMT1FCf8XxhnG+j76EG5zqndgi3UZaYXwvLHG4+q1qunevCzsa8Lv
M72Iml/CQ1UhPAAN4Sw+QfiQHv/9xZot/fOGdhJB8n0xLjJmQd3tSXwQBRlVZ4OtJRZ4uLjXKcbr
BCji1nXda5CNc8q8sQkDIcucG7HmiljtIOmEhr0LFu245bhf/6UyJuop6W5znkmVJhPD2iZoYc5d
4agFBsQ9qC1jzBfTFmLvVL7Xb9WRqxvolJNeGr5xPIoM9RVvvau6uIabB+LTOWqRo21IxGG2+c87
dwyAlVgctrvMcVzZe4MREvA7I8I5wmSiGPiOtcwijg+BekGPnldeQygQqkqfbZucrZbYodVYXp1Q
Z0nfJexydNbYcaNegT/MVmnD5Zrxau2iewjw8CaGl8ejPnQHuZz7V/pedFrM1clZtYRhvJEHfLDv
7C5KKPeQOkJYugSG6PBDYSsJ5iG7DnHxvrGkT9DqIIsxmOZkzt6g87AqZ93a6rZK3rrcUTyAG9yU
XWUTqMacaJA6+eREGGUzPR5MMOfFaNv34eQ5odUWh/sQJwPhLS7k8u5l8dYa44Duf6zWPpB4uB42
/WHAl8uMyhrWOqd0fXuKJ+oVabvtK/rPYN+B8Pz5V7XR+5hkjRDAeJT/MsFI8GYndx6Tl+dRMHgv
7VHdAUNxxBNKtNlN4WSP2Xk8QLbF5HSSLsccRRnEYcAvO8nWUpZzD57XMhl/EnOwiSWrS1lIjeB6
Pw78Isjkh6vT9732p/KUr9tRC3hTt5BF95a/55yp7jIVzKQpfcMD2xh7UV15+JjAnSSDXBaX84Mw
gRLJ8pWqqp88WQ1zdreYoRe9bb0Pp8P4YrV262U2xKF8ZWTzXIARZmCkjjfwr6FwMnwtmb2na84s
XdlYvib5IJ2iJ3jzEr7i+rbviMVGdi76hekS7BWKG84cWTFwl+Gmv7dTR3/au91gW8FWH2etLDjZ
AC3aqDTzMTYkkO9A5uzjqYJGgGO4YikAp0HUreq1IDnsWDuSE4dMYAniLQH37YSkHN7hjYQbLNvz
dkTCLvYQ1YCM5Abk9HWLiSxeQx6twHbKvDLTdbrq/dGPfeO6YfFtvf3ehbHUA3AB3q6a9Eim7BgA
BZc1TDWA8lAfenGbxySo80BQ88C0zJDXHJRZC0AG5NIntHe9+vVUgxHQ1TB3O+0Y2ajFljIfcD+o
ompFLb3+9kGTdZy1VDgHJmuYFyTEmHPOFpuTQf5R8grb9YumO+92XI9wpa54drwbTmKh5JMj7mqW
h5G2l/XijTYD/ajJHIYCY48xCM+PvZnIlcgwGabN55J1eLDctwpa94zfvZ4kr62CfJBw3QcLtVEL
7BvCYu5zbBftv1AnmUiPhIEcokMjsO3evVO3I4xe2vyI4QlsERZ0CQ8krymz08emuYf4fLRRXC89
qEJAx2YxKg82Ml/m/u1ssmYzUBkzqLm6QOHS3FgREcrfzQYkxkvTU0/yiVRraFeiMtZd1EQLdJ4G
51/W7OxzJ3bZ7fS5Y60eBJ1SVvvNur851omwYN3KYKM/zE8z9jISRisYbUyfIFwW5ot99b9F24TD
wRO8TrQG+/KbiauPGLpvPbT90ETj4Vwkg8/McUiQVE05guPpbNZzwTnljPa8lnBez+HjhReTL9U/
0gpDiq/DFgWO9M1HkGk00ZpUorvgYwRVoUEGBjsOjKpUx3RDNnC9CUEr/YHwYJhs1eisT8UXvEWL
jvCSB2afvSlMF12GQx5bq5ufJeRHGE2CWbXwqsJHxofgDzfUkKi+ILfK3qTyODe3NTo0g6pACe9V
P3rglC0yhL2Pf78jr8Vmw33RXgJXro/4olblcK3vTN8L8qIFb9uluW/J9ErWQw7A0KcBKCKWbomE
SfbSzPxefDwOiVqnFhDKZeQtHz8voZ+Z6r1OSR+4JIla5wlE/zEF/TZDu9lZltq6f9kVHRdsPNPy
Yoz1vCx5nrSfo1kBN7fpljc9VIaKKl/Ms/nc1sIlG4AQuSqO0nqmi3JPwc97WYZ8kEKg0pDIEyN3
q/WOjbcBjBSpoVKh0aaiu99RVhCVFp7cYaC10A4PQlFadSrmvSSzWu3OAfUBSTzZebDbyAKej6Ty
TfEWNDFi6iQ9yU7g68inMbO016mM7wS7yzQEuQX9tRsJFP4MRS6R8Y1EdNFFuZmlTd7vi3BP0lWL
lq0DrpmZlXymRBOd1Gj0RWzrNwcrLHiSA+ujKaDV+F/MJCIOZ7nL4n9BsERVjcxNHXws5ZKimXyS
xJttEvbFLIwMjZTdawQIdITuCBGg0ODeajjfKyvAct8wu+BqlF7p4GBR3G6iyiZ+D0tIdRmb5O+G
vLtq4TlrjXaQUWXCEgyPzUYxOcmdZCahqil5chb6AnNRFHIo0ZZ30Cz6ifyAd3lYDKUWIZGXU1d+
OG6YZXk6dn+XEIQg4z/GSPWRDPvGe2dHQZW2lkbPPmcF3b1OwUCamUFPmA3cyHmie72kR/odeGi/
W1Hrs9AI+WP34br+BiZ8RMsrNnMB3qaUqPTd9JUdraYcAzWWAUxAFd7zImwsD+h/l0uVskpcSVmU
6efHmuEoE9aMTEjpRRiQXZSzoURbraEE6ljUuh0VTlgqZJ5h8heHL31X8NsUVIbBST8bwRuLgDSy
bv/U/lU7cHXHL9tduvPtO57qopeYS5cbfUsFyQo2FdErFWAghgvzUAfvCoxa5i59v8ZU9KDhsqpw
+0Jx78TGchiQ/1CPtui/dvae033jlgUZYCdQrIH68uw53BET/ohpZuSWBoPqjPQ/KsfyoP0CjHZu
nLEAtwYlY53Q8+saS2DfFYiLEXWgyG9664E6c87fiS3Ih+rcTrKXW6YzsT2BWHMEoEYsY/kpdjSU
ha5rrYdibztZ6RKAJoot2Y78jrIwZJl67NChRYbp502le+4wt6MUzbfRTmtyNg40VLce5hAaZNSS
XIVNPq+DwVfdUSroO/G6/luerkP2yYmhzfDPDo/QHYHPrsEff5IFN2mlUZbvX00xYeXwUj7Hh85w
iubtIyfzGBsQBrtFrafQ7D7CuI5hayopmC+ez+txldGNaM26y32HgM4fEqQlgkjC0hLk7ouGLBY1
UETWZgRbkGoItYciGVGl+K9+2PUsy+kqZvHg+a0t53mtgzfIrhEy2+JOshOr22Bkk0bvwXXDealM
SMsFOLm0pWbiCaVGAI7KiVhaTK0xU/P4ePGGddT/c5MXTxBXyRpjfMLiZj20YZZrzQfjULNJwFQO
4Ce1WdddNd/TlHKeaeKZPYprBE3RCuiUhdr0JzKmwqbgFxN9/fGHGL1h7ObRjcD6ZkP/d7KcO7Km
zH8b2ogWrQ3WPj9YRycQRdyx1T1H7RjyKjD81pJjJ4kzry5Rot8ULQKRkVdbuyfQd50eG0eIroER
kElygV7Kz1Xub3RyZfbHFE3z4HPPnm7CA0GUXz20Rfha3iQrfiPxoXXOAwCEXN4JdXcOcKudCXW1
tK7aDUI1teOksQojFJn0BPtbhYvO3oAZ+Cr8dlPmGGJueQx90GE/NbV27Btwl9yS2+EJBttcNuqz
qr5qUrrFIIb6v4cD8PzvsUr1wvrzVwYgrhXvttEIln9tEmzACH6ltqlD8HEReRpZA/CNeoOTCuqb
+HlxzliPHAmejmNzlShJBGtTY9km+qH+oU3E0Ro00kUWvXkVvRAepkA5GcCbbyzZeCJT8QMRlqN5
l/vqP2Orwkz/N1Woy4CKBsXWqg6n0cKkyZfw+Hb+peAZKnCK4fe0wdT6RTJ0Tj1y5pxdf1ve4lae
aAbrV1ej+Di3+TXUTE8ZLUdguw5ip3E5tEKZBTOzKW0auYNruEp3efUvW57UcRkHCNgx2WNKfeQI
BkcwapHjiCVM2NleE7eitpneVd18yIWoyF76cXuJWZ4mLJjy4LNKH3toUgILRKeHEVp0r9VxRIEi
zxP24+LET3TIQBk7CmBzeAyPrYKiAI5yr/+JQrG+gOC/BY29J0NBUdQ5FkHa6hAerYThJ+iWdbOp
UKwpM7SJZzDUcCEey9YNBlInmV2B6TZVLgv4Bi1tHJLwP6z0IDd+DxyIseZKUVDKg/lnJ/pg2xp6
05l9xQ8S94lvKcwP5oYTqz5uDcFX8KnEwhdUsqk038Ppsyh9lVAN5APsv/fXvue8mHU0MU2knUPz
1idaG6lpWSMZpJ5VMpnDJIAVu0JawYKZgED3W7QuLkLS98FFw3iEGGRMDPn4f3PYz54d0iAHtqgf
AQlRkl82mtIuowvm77Yv6rply80R/MJgQ63yFEs/SqtB2xHuFDQJ72TUMHVL2AtDY0/++cR5Jm+6
IqXAN4/IEoId4Zfr7RQXfv8TUxemkTUlqPSKjjavHL8zZfamC89oNTV0EJ4fLylw6lNXYrZe727A
NCJdQtVQHaTeQDhYnWqCaMu/4VIUvIpHCOmx4wz04I0+lU5CrWT2doz4i5YU5L+xLUjOYNhyTDE5
NafC09SYcZ4KBGPE8sa5xav2a/SHHX04fxnkWTfVHZve3wGmnXoiTYolXLNC2P3iLNhXYZ/YMgLo
mTQMYNwau82M1nQUo2LnNK9m2gSvBM7RXHt90+ZDyvncNGxi/pJAiNAka7iQc9UhBt98fSuN4yr5
XCzp8Cw4/wxMttlqsvEn6sxREsjgK99amvPUsqbV8OSw8nnt3k1eFGXwFoq5MMcY+RtKa2HI8QfN
vzZF/VCE8IUO5fTso1p8Mc4sFK/YoW/x/otUKanni0hxWzn8tecJWlCW2734tCNC1f+uWSq/Aqbp
QkBDTHGaVoDcCgoIO8LpsGQhC2molhdw3XrA/VaUY16uZYVM3grn/y9KUC5MRz8N0UmEQgpM0cwS
+mBu6ToTdfM10JEByUcH/0haa2JSjvK5HsKWNyVu4tOELAJi6psrS+ppzxcNcuxHIy3w2aObxPaG
CWBDZ6aFWxjDizAWIzwVqam3Y9nQ8WspOnYa7MhskXfAgFxbzmUWl/j67Iy+E3JR+NzLZ9uW5n1U
qKl8kFbe8gLwWb5utVsio/ku64MMj4F2VJjxUu2MR7IGSZVSFrMtHL1aH7V+N7Oi0FM5tlceff3g
e7ldopxeHnoWliQYib0d1K6b/lmrAy+T3/LeYhAnG/uEU2LKoub6d08+wEcu3CyONlBZNYau5RZg
TSMPjjCWUT39LwqvlmzEYV3qgFQZvQqDMJlaDwIqOmLB1kSRBPPDb1P+/3iaoJUVCO0vwVtjj64E
2QP9pYWMoOmrZBDi56/nMmTBBMstlPd3Z/e1lQxKY2e9pE2xuYXewbJXAPU6cbwjVJdm5ESUR5CY
e18ryY0JSIpy7U+aTas0sIxtxRVaTZjpTbNVztzMz8RJLeEIDxe1UL0BeSbqboH2LAKqy0UdwXzC
b3HTJNPYF5onf9ns/OWfErFa838h7FdTjPGoNCtVhlI/bafyq4DU0ABrDjlmyX9hyWLRUm2fLJzu
xmaATVNaUEVEgFx1SwfKKOoKeOZSpAdUengpn91JpQfJwjZvBdgKQgzPmXi/rr7IFebTRqzNEoIq
wrerS9rtNDFdSPC5U1Ffws2UYYHj6nhZogW2CI/r4cng/8oRxVMRky/WcD1OhP75nX7PtZBRLGRN
QGBdo7k3YJRHjx8N7UIBMbshPswE2+jvV3ELqPiQ2Wczp4FC89Zosdm01XVi3hp1NoWcpcDa8H0K
fUbVK2tAjarW4XCwJ82ZqoBrUMeOKr8W5WvEBdhjMGiq25W5l1NORLMc9KTgePwOiWmzv29kNBjC
i2htnGkT5FBcbjr3IWoynq7vCkgswGLAsfiPqpkHTfVrF0i8Sn8i2zCCHsaVj1pWbvbsirnd0uvU
5FDVvLCgCw+HbLlX1GrAw+eogqKIfjNbROSp49FU1v1M1WxD9reyhxZRC1M2ZeNWDXVelasazunO
pOi0EBvlREpY6du0VBIeV07LRsRvsoD9o25D7An5plyI7obXhdPT7a3EquIjMXbiv6ucovuPTidm
Cv/gWlZCCwoe7eDdOEZRMAkhWA5iotUBYyCV/xyp26sbdhvNb0S+I/9//oRJrXNy6X1cgTu0vYGY
caWsvnFtPLbmpIfeDzFurVCeXmfoENpp4XJYNDCoy8OitdOWulxeQeiYLhjaZxkvFFr3ZLxMS+e8
Z368UAXb5sWSGWKJGu3szLVINopPpEsZlrCqc5pgtxnvdsIWrzMMX0iFobDOS4KueaPhu/Vb445L
ZvVdH9pZ262uyZM9e+DtG+85sXy7g7jd+lFJ1aMhfP9uXN7iDugERosbjvVLWgT550pg5LT7uUBN
CEJ3Fo1zQ+WMJUkKCV2FuDYNiQFh59w3gevIUkKoxdsSXZWw/CZCvR/IKbDgDn/9rtwgJT6Dr8Sw
d2fM0Dar5ybc1FPHIG0lLH3e8MQbKPm7XRhoZnOVEMPlh+Qux4w/XjxJf/4SocnPtTkU4VYR/K2F
j5yH8qM4X24ARVi7hUicYClgSOztyGqgqKbbOQm+nnZESkfLYZHMYdba/IoIx1tdj3nkxXIHxu4Q
WiDqlCTlvD2K3WBk3eoZ/B2L/p2E4jSDoo6gT9JBCvEXqQW43uhqn+kqYjGZCpvkhGqFP2l8ssWS
OHZyIixWQUg8JS854xjqpJPb13Uq/0I/I9qE7/oED/Z5Azj5vjwxrZ1fV4ALkbhWxWgH35yN38Qz
MzppBlIjCxVt7E4W0Ihj1A2TdG9SObWNV4/26MKtjIedq6fXyxdEQI97NKamrIDoScI5P1FprQOP
fqD+IVh6ElsyZgHcSOfoexzqNbT764FDr5YyBASdk4JuT23zwrVS6nQeU1dFNhPcw/VYLtkLgWpx
Rxwc5r70OutPzBezyia6H20PALoIXWHDJByuDQBjF1uMbgWYhgRJKRcnxx7ZwoAtr/ySJi/HJLLa
UNxtGsVUlbWzl1Mfx3JBTo6RpB7+CNkD2qZe0KicBgAeml0PhELRamvqa6opH7KTUXWSunEtqg5d
KHZD2+TkX9BDyMkobU4u2e0lgQaGXukgMzzEDrQZOkew22QZ8u16VyVwUyu0JAzyyzYsZDXMf79D
BlnvXwnx67Ail7mo15T8iL8pnnWwNSM2uF6oLB6Xl1KdvJwYQm8GtvS/gNsgh93J2aSrULE+zX75
ti5ZZcH2EkMDCXyjPo2hcQu3MZq7FQabgNhGTr5zkG1gaaJhillz4uymkNhgAh3YQqmzEkCH4EA0
aAXJWBtVKUyzkSWvqJoSanaVAossguIJ9PfxYCe3hnf8i8C5ms0cyJ8lIx3/yjNCMP+8J3bBDG2D
IBXVLZT8go1QOdo6j+3IKQRSytLx0XtEMd/7RQZ4H54j+ghTapLTg8QCRFAANT5kC6PunB46ZY1D
kNpRyS5FNbE9aWBKpKJgk71So6AalSLyRXn21v6UCNZZQjKGLc/LEORoGDP5ia4t8R+cBkNHjUhP
+qeuYH140y8xZzAUCIitE4tlYXdNx/MazxWWaFHLSCKV74So/jB7rWVPbcoA8sMFfwp48KXL7ejh
fviyGrzogYuLSLbtLUQcfXtPTcRExBAznTpNOHOvFoJYEpD5M0qyegDGm8tyXUHH67eHAoq8/vJv
03msrAL9l4FGOmlyXZsUrNojeD5ZfU8l3FQe01yKuYy3Auw14v/G1oEusjhJIITvECtstYJtnJn0
VqScI/Rbap5wn7XIq34n7s6A5HeWMfLeV6EuPhTCXKfAwioqJCuvGwOYj03gCwB87r5W+InLuIdf
1vFSfyrt86IRPyKIIGl6k7SI/G0biqvHPQFKoudaGL5Qr90mPUzXiCU4l6ttqBqrg3EKc0Vuo42w
zwd5/qiW06s+wm+ljm+elSemsXRowzd1p7invkff5kox4aj8TAjC3U0Js9phrJ55YwujpzqOXzGz
WypYI8d7pDKfifVmBo474gMNzVB5g7dpJtTsz814MObspdpk96ge2tBOo1RnjMGlivNhVTLfsMyQ
GG+EaPbgkfSNoDj9/IoxAFQqAffjnrRaqu/emPbO4Igni6x0LbCOFHHeGPdWkSFSi6ao3uZDADFU
wdJg8uIDg4Fk9WyMrtwHj9nS1Mida7cf+TX++T1rKCyecX8brTtD5+3d/EM2mCCkPCLigxU/bjQJ
ri+S8mIXL6nDMZMt7CCTV1d/kWsuito8MM0ke4qotUYLZA34szNij4Lka8SBBkiIHwQgr+8+ENBk
IA5+MfZzVRq4a8BvIo/Lhh7nZ0T7EL4E/jgAEYBCoJuqJPtytVLUvy8XbwGcYBNktnBu1iAGzs0o
kxt9Qz9yKYGbARYDXZIRwuNqN+TJZuWOtmbkXArrjCCLqPc/JBfiNgpSCgxfOUzPPh9Z1MEOjVcX
fHHTvMVo+0/4r99xiow6BSy0WyP62IK2MuqxnzMVNzLWz3M7s8oi5ygxxDGtUDfc7Adi2tpcOBAf
9mkHMSWrLtRcsArRJ28q/IsYjowOyAzgoLlHuQCGW7i18yJcwoE+mLpfVwGvmbocUdA8zBuNWdG5
9VHn6ut5Oq2d4rpSb254rnpv6hNF7Dh10Twx9xEPQfBARTSqfptWwrInHyu5D4SLfeMtcMUu0Z9D
ifKEv5YMUGnfwfw7ujveMo2TqgJQxDvINBXAPbwGP7WMHhkAfRwh3s/egHl6pZxeqidJi76leBMO
0qC3M228nE3/4kbXgrXvl6d74xeMEvThUqWSSz9qq/LQ23tMIxzFM5OlpCCtr9G/ZzYy96WQBbAO
A+6VTy3Qem4uk9zZXFpjVbGwbRR55yP7rroGQ2vTp9vufUMHGGUldh4pcKiyCYJFBdCfgMD3/2jy
xp7Qz7dKWo2C33mjy1D204gP88rUr3D7iW60EHchXG85bGZZyvBzXpE6bK7PDVTunNYQeyDl0ea+
lj+lIcNTdWmsJhjWp1wxAL5z5t2aV7omi7tgiyLeKQS03xgO2hQOmiHF9/UyT6addsI5xSJ3vws7
+/1wXhtSbp/dgfatZiHfkXSROm4ASb7BZHDd+ThUGx3QJVNmqBTXASp0cXP8CeejQTRusqq9zbwv
AYcz+gzjNTUi7TjXHFkB1U5Zlkva0w1Gdb68kwBZ10HtE6kHwwarYXqYFwZb3e6fRA6/Ut+/eUsS
nICKy4wma8f0/Efwi9vNKODIUXTrAc2swqOCeU9hBjmHfjPIQM556vI2cVc5pXbnYl0tWB55lMs8
2s7y8KRhBPPvbnZnMfpS7uYyrr/bif6iIA7diPZiIdMmr/uPf+TrN2Rcgclb47ls2ZI5GRhldiD6
XvvISWG4q304/3vEtUVU90QWY/5Bvu1VXgSgTI0/5L8OR+itD31f7FNp47C8yMuxVR4yBZfh007n
1OAWCor/+0gq42Sfc/ZHSDlFT0XVdok/WoRigf7uhsnYggZ3eIX6evRNvdoCzCBaL62sflTDmaSK
GuJBMqvfjn862IUKxNv+yAfXAQZUqgztD+AbcAh6RAl/uT0kM2n08nmy7o3AkC+jk9XtRnldb/xT
ueJ8tedZwWBzr0X+XVvjUSb+xCldD6G+fzx0DFfZI5nyaAWh6AZPv4bY8reCV9W+ukUxm3x7V0+b
BGwT98aq2wVXjvgTbjPM0SqouU8hoJmx3gj4wzF+0BE28Vc4ZtsG2S+k7YbWTkYdLf41sAEo3B1x
ePUO6ZrUeSs8eq2kKGB2emRq816GtEvswbUnb2i3ma6hpLlFTVJGaJlhexFbvez/g8c5ZjnAzOWy
7bwAnsNJTI8qAKBDMaqUbMXTZod4lUEe8M+TiwujNKG5ZMB4jyRWqrZAcvPcvASDohG3LRTtRqiM
Z3NHxAilo8zs17xYHlXd5edqxOsWulamAlug0IIF9K37c3TQTbeGT2dG6s9KIsha78v4RtQ30L7N
wnSDWYITvFvyfW7XRgcs/yOAkC2Qxk4Tj0L2j18SMYIpq0H2oblq/Qf41G8S3bhxYE52xggPMqNQ
bbofhLNRnAyUHtkFARrb63X7kYkvhTWiv1dBG1xiNVL8Iq1FLDDHBn1m2eER2iWgJ0CRjY3vXAjs
y1ZM6Py+q3YbCPBOKxGmQ8tt7mcR3+9lTPikQjA+AWwHbkx6C/A/I28frDyBDX+7RtfbPIcK4hYU
ACWNH8FtB3Oued0rr6E73hw2upBziKy2H1rVydhAzgrDJ7jOOl6m+eOnbZO+HWce25CDESouqW6x
ePeYlZGOI20s+qvIcCafTZi4zgdq43zBDGEghyUPEofYW7pj3OCEi8KaUul/tr4Jpy/RaUwUdt62
asySquDJx6E7hYXx3waOU3vSCM0KlbjWEBgDL1Gb71Tps2/KnlCtwkcznIAGldscJTqPC8xN4cSR
yknMF7cE1Sijh82kkBZoetsEc/gvLpPuNKlj8uR00XM2wM4IUZ8Lll5P6+02sQn3rbl2w9w0Kxo3
/2T8uxkXmHtlGr00afmhDC61kE4weiluCYsDREHyWoG91tDIyG8S6bhFPOnp9VInzY0pVMC4md/m
Kr0NYL/+ALGFO7fdwMkvt11iaXuwbyoKy/Bx494z+ciJB2V41Gd/llDQLr5DEwwfHTkHYc9bilFR
rILvWcFRQAIkOWigdG7YnlLszEny4fUJ47vJWpvYGoxWVv47b1gtQfU/NrHLNfsVhG547MrFtLO6
ninTkrI8gQFnIdPz+RWsNa3AIiNl7Z+53/RE0TXpE6jhRVVgBlHpkLSeZkJ5QTzSHvIhhkdiwjPR
QJ5ji9EP71l3bw0htXeYUT5lOSBZc1PG8NVha5BhCPTCJwN3xoVLAnVmcuEc4uh8RAGOmyXb48qF
i8u+qPFaPTMtITPYnkuBsUosSr4xmpMCnw67gzSkzs6gcqwhB0zEMfU/pqumyLxLRAWFVyaOtE4V
SAY/NRQjB5O0Seu7vnWE0FBz7f8nv0sgLZHmF2EH5CglnBEWrE9RCqMwGaSoGcZke6YEOxb9Wo2X
BEQeH8UwD7r7aviY2K7pDyH8FuhofsbPfjmupPxgyCMOdE5P8guBpxfceacTFP6IEiMnR3Ev0Mkv
F6vVHMd7wRMVbjfAVnAqWcxYwpHgHn+fMr++j3GWanOjlxfBHm9Gg7SZN3bFf4/ArY6CClQmP4/P
uIyvPIlpkbaO4bjnQgVjsdMc+R6z/C2VMq/8Rm1u4OrJc9mOXIBxbxftObCic60yh3bzboR1AOW6
j6x5+UPmtln5gnZr0VO/1ThQd7WY5GLPTJ/xR3XWJrRxXHTzNGHSabYjQr8eWg4OUyEfur2DpcOW
QXKKdGvVL1NqiMiaOZzIMe1Au6AuLC8LKx3AcMTN+y/46gyVzOI4lioKtfJtPc00Ukiif3ANznMo
rH90AdFo/gnQWRW5IMqX9NAkjBI7eudiAmNor+U2mUtFjHPRjhGectFIwIraH2t5a5zFUT1Fknb+
xF5UOzZpZaJ8GXIoQ9abiXb31+K9nnMkSzkZ8NA0n6j7QyO0qpnGd34hbPWzO9BBIrzM9B6iv8ez
ReDiq3P3t5FkZO4JHL/sxyT/1Obr+qVjHjXAs6/RGRiN9YXp7SYxNTe2P9f7+tkHlWkFIA0LkL2W
CeoinQkHjr1Wrm1vrtB6DRRUooYZ6a+EEVzcM84MkvGIOQOGxwvvYRGJyAodYXK3RBM3/jI0C5eq
VsVQ3eL0GiJGlpN1W18y8sW/HRbq/6R1gux6Ega7uq0e/8RxYNeH0GcVS4kh9D7wPUD4+Ywy8fO0
ob+gTv6PgOQSntPTlFXBOMMmQS5kkOx+8hjU3G3kVzKjl1b8aTsQo/NlqBzZCNUQ/eLkJhDPFJFW
+Hg2s0xE1oo+nzj9BwZ4LVkSoQI0qbZN0+CjAkNlMvamTkuheC51Q3BJ4t77xp+i+aVceYPZKA8f
T5WN+i429Hs5OWiGQfygeXd4v1rKiJSLd9IVUGfgFYaXcaN3dMTjZB/qoByAqk/HZOPp6FAwCtJ/
3qK5vGNAuS5rHQ5IqT8RQwMW2scO05z5CsrbpuYsf3Jx7OOapfKexVXWHq8EvvimhQbrKF+peGBE
1VKpFZC856mnJZFA3fG6vD0DmzY2ZDo56yxVRoF4Q3rajyrRNDxccCuT40FJaeY1usx4vdAWgH2/
C/PdBpf18zz3n+GW1jqXHTe9G3yt4mN8dMh6IRyUapkUuWsplyS51IVsFYqyDl5kg4T/Y0LC8tlp
lTvZjJhq552ZQSq/RqvcN3gCqYBLsYcLAkf38oGORYkPtJLtV6Csy4/h3PU10ghDN5rsAbKQVTI1
arSbMpbjuA9vlkO6Ru5SxvOsDCqkMquC8HeF7Gee1zYeEJWQYZS/oIvgk/g6aHYZeVeJ6NOEzirs
5kwE+Saqmsg6HqZYTlFM+xlbucBNPPxo5vvrY++Zcf31Eo9wSiuq80oU37FCE3yRQuzt3+cxPP4a
Xw+7xG8ihZXOnnThTgvlughxaDF/hptmAX9Ua9Jntoz7MAUzADgbZhMWrSmB9sLQ0rK1AnyCS6wq
rUEA2HCOgKWYjXEmaMYHVi/jfCZnkGaWmKqQ6e1V/PbA/SJeFiOd5UduvyDIjl+yg+Kvwa1KeSSD
oR05JLRIBoayU1t8ZbZEd26affomKYyYcWABrVirH8Dds4ib1yhZ5KPkB/Hn403M7fmSyb126zfx
YGUgMmCzBUyXzIn+JbpvTiT1BkQZyn2yE3HApT2q0lBX4nVpGSWElojjdg4ernPMptNsAIPv6/Nj
zfNXclYw8tGAvwmf5wDY5hbGUsp8ZLbogMk5oK9d/ns2M0UURN9F1QQf3Y7VEfBZl3adQYzSmcJR
8xEyK84i3WP7GFmY5+1xir3ijxQf7hQ/lrs09oGKI3hRvb870H+wEV3J2dBP+O8MnE6X6LhtOZaE
KLszhKeREHupM5LpqssZUAKyxirbkAVxJfS3r6zAHuqvMHbz2x3hs4LEkE1K4cHI3/S47oHVlbX1
+LkTRw5twEu/79g7kj58I5EwqigGbm5DTqshrwvVtzdl2K5pG9vSYdTvS0UMQPJTN98Om6LJeykU
jgjOcXnzyWm4i6STji8vs7fpilIvz5JcQwsuRTC4s1vAm6F53ZMfkn+eaACZ47Z5HKYeuKEoEMzt
lq0Ckf3jSOZrjOZAPuXPBw5WyYcdH2ca1Tt3WhJq+iX2GyMfzip4h0RaW6KJBIyhqH3wLDTTJKod
Yr/x7GKfpC0lSFNkfSZdwzQBOUDKPWUXMU4PN9JJUQ61DyJgHJvb1DRyKQuq85PoseYuWP7X//ap
nJq2jKlvs4p5wYsGlM+XN3L5sYDrs5k5ec7253JpHs795Dm+vwt8LSyuAnYcaVwgLpH1kBa7RIJ9
Y0WKWhbRfYeBJNcBHu91la42swM2FCKob2xw85V6WsjGMHWfG/Ikxar2BvDgCUCmObcMBfVaR8Bm
WE5LP76ZzV1ClZEFV1otr97KKC9jGiw6CMelsHvqKwRE4e7M8NycpO77580cxpL2a8rrsDxmfxgA
UEJUESgKPfzLdMPNiB56kSCdSUrfhprKcQgKvD1dRXn3hL1KS8GRvz6l8D8HtYwEhd8twB5Eov2J
V8piD05Y/8xGz8ORiA/2Rqis3IdQLJ8XZ0EVyskH9NHovF6kM4dM8QSxezLwJ+v+hxSchIhJDUmw
g2fTsM+6G1hLqD0xhEkvkEAUCzbF4TRdCvkPMrK9Z31DEzwBDnqFD7kpd1/SnUqVfzUYi84rf5UO
qUarBqMyWXpY5+3XoePLO5iR4QzqUusoYPMW4UA8S8gBUWLjmxJeSda8O5kUzCCE76WN9DyuPhBM
vmVsRv20YmFOs00bii3hdqPYBFj6MxpGmRNKLfp4Wv44wSxb4q6We8ZirKb+2dH9a1YlqRvdJXlX
kWQ7Il5onn/TN472vS/fxtAoYzi6MbrhsTWj5V30PCKHjhd21u8EhLYvpFoYXpxE4gH6j9clkHZS
eAVF2yVGcGYbUG7lJcegJajNpiLcBOHPgghcKr4746GIOr5qSZwdXbZDIVKXdeafcNDUdiAXsxjP
vo5UQGYCASBBz1yuCICb0V7JEMAD6Uz2QJRRGm12nYfBdjqaFsKv2E376i9OvIV4GAS9Bqfmjpzx
czP7tQpxBqVNPEwZznyelgPKnkNjoFibFFP0RCijARjGlykNicSIaLHrt8Elae73KStYnlcBWgO8
w0Mzx20QQfBzbrxKXeN8MkGLUk5R9n74YxrxFs+Cy7B/97TjBWcejZR2s70AT4Rw+3Ia9Rxz4CPK
xrVE24DR8mlGLgZQrKuqgqbhvtmlw7tdDEFbkKHvUOxMwWeSVt9fkJzUBlPQF45W3RRFceb0oN0a
0G0z32XPgJAXcUXj25Aw/KDv0ZZ5wFa7zZjpcMg3FIWO3A28VPuyhTJNnxjGlZZw4rWzvhk4FWT8
92cBQ4dQxeXgUzVjbsIAvb0E8dVCg98JCk8WsN1lTTAc9rP6aopbJ7St4XIfic9/zx7IUiUPmJ2y
zXRlC6Pq6RyJOqN7NgbKbPeSdNqknS9b2zplpjBeiU4XEWrEHSJY6bljL5OOryuRcGSxBVbK1SBY
8O/RVKnH++oQXRoIFj+oZm8mD5PjK6XrHad1xiuG9s/SN1X/C6chsEEaFy4khVHC86j3PZfJHjNk
Uz7h8KScThcA2KXX7IuG/U+4Lo7Iz1qFLYdnqpxX1/Fl3XqiPh25vmZwUIAV6Oq1d6MkIHFc6K5v
Hb5vIR9GPjobVCdlIjKc95LnAzOUV8Di1Aeck3jhsoTa9z5h54ouqa4f21MqFQ7TpGVkpzXfMow9
n+cvkwvirzXjKT/kNiMtHkbUsuA89i8m/OR5Pw5Ncf+US7OxNBx88DhrBrZRQ6U0+sY4uSFGLWhK
QDOT9y8JGI8ljJvUdYVZgglsT2pIE8VumLdOLIiZUaPRUnV0dKnfykmQ+bZ1NXycN4QNk36g15qD
3/R9m9RJ1PgnAtZ2A4QyBPUZu2fiEWnGALyy/XcNbMWTnR11xozGhj8A+/1G80+xusCgi1vawyTQ
yRXiN67ozGZTcA0qwGEU4Bc/HFYBbadHbYEaI953TahNs4B1tu9beg7Kjhiu0PG4bA07KeyEeO7k
6PPzSwOHISMTJ/m+SsowQdIPNjH2whwOIeUlJc58GLneexcpKOtP4iZXT5DJNSh9b4Kg/VmE09YZ
XMNJ6G38sRBY3t9ANJjI6IYpR8qEV6vb4QnEo6PqdUqkCS63VUe4o6aZfP7Wrba+7TH7M2ynAlHQ
nwlFDg8pWLbxVS4SWZHWDLi+u4Cl2gy21LZ17knlasevpj3K/8rhX1Ya+slPTfc3ebV1ztYeVCCg
3/c0Y/vw4/c3dmPG3yYsx3qEiOeOazP8IDCEtdv8cr7GNmgI86KNOXLlnGt1aaoLwwK4jTvkf9AP
m4WbbOlt0+aG7zJOw37spHXCi1Qxwke/MozeRahXql0stScYCzYVrpR3blbr0dlO8WeP8++Eg/et
uxIpJOWUj0JiEPnOCIiR4aUl1+Frk0QwlcZDeA8jlQ8GneO7v/zJ3D+0vCYGyZELByHfuKVzjEFQ
lTbJKx9wwE9xlZcu7Aquvckj05ndb/LL3xzQSQOGoQxeMocRaO5Ru+CZ8i7u+2VPdcnoBqGYcWZn
lwGE+FMmVfWVTDsSiwcIpVeZGKwCoLMBgr6q3xre2aSkoSWX99rDrfYrpjPR9M6XiLBx6U6QGI8q
VhUyYskous9sjggj8IBM/PuU0USq4V8vPTgGq+AeDbR5RcBRXItzB/C5ewR6AchvxH/tF/5OeDgU
zdsFxsXH6wVx7BoW5WbzY6su42qsmiNBJpgiRIW7SeTEeRW6NiLBNgyRz7H53i8zZL2XnlgSRyrB
8swm+Q16m23o2pbG5cxFtIOdio0zHaqJaT3T6heVUUoigStxSfulgsSGHDCSKICDobfEtXkHE35w
pGEOBVPQGNUpyjZI9oMTIUmjpCw+TIRCe03IzetgwVsL7Gt+94i5SJtiJvKsf+eHgx83h6iInCL5
o4xUZJwC07LHNzV1O8YRyGSs1rIuCIwNd8pBf1oX4+Wp+Rstc0g68REisetZ2IGo6zUO+74VOw0U
wVPsc1CBhx4blCwnbhp6jQtwRYQ9y901SoCw4SlTA9n/LaApsC8i7SLrAgDjLZ0CgumqPJrzTE07
jdcXujPUGLfOL2pWb9oGL95utHHWaf55ERezSvoQLHzAvoZSQSRkwlS55ZjowVaXqpXMq6ugutri
Ngw1aHI1eychSc8QuEoDYUrOyMxwBeLDBUe59EEmFtcDN3jfjJWZTAi0Y+29XZni/D9HkzMCEdvj
ApD+y8t6RghVyNoYJJGwJY8lwxh9xUXaSIAsPdJDtTw3/ozPy0mLpN6VZ9s36aX5KyXofcap+tvT
urTTf9TsXWHaw70Ibng27VNatFntnxRoURgivMmXH2KMuH2adzLU0DaMzW7T+O9Lcq5boUZFE7as
w6WLkaeA4Dt5Iygk+xVrB+u1s0hPgfyMyfOg8C3uQqzElXyaapS2VgAimTNKntiHfFqLivpa0x9i
pfMvAknQ6NPyZnnHWbZNlpCyAczDmTLRdqpj/45XIp2OhFoTQyCnsju4x/DgpkGUBTJthVniC98H
A90/x8IsyrMoUePqEmFylSFMycwiqunueSeaX05V+q0SwkuphzZI+7eAiHduDcx4qLGmY4j4AbsX
xmxjblvgIkaDxgqG7YJiPq8QIPRF6+GPPEg0HbOI4xeWwEIYzDmEXDMq87gfgUPbPMU/YbPKQo47
pW6QEOAhw6SEmO6cVyHfEDEzFar8L9eS1/NlZTALR1J2JhGSVB9cSyNKxWhjQZcOVp/NUIraH4lY
j4mhVC7vC1hO4G4ySoRZs7Ha5P7Q3O8LYRd6i4SFTEwsRtGKakFbVbuhtB7kODUdifz4fqgYwwfo
jpi+fI7YnjwyAsKmBa+rXl3cntHIBbOxkvEx1VGg01RK2tlT8UtQukB3jkD/uDvp7kfrqw1v6u1b
TiYowNAkK3DoU9PPZR+g8S3FTOeuUsACxCobHilvwzRsAufXv1as+VEe12eBy/tfOiHCp2YQcT7m
cQ6rSGo60gv4dtV9HnYPJz/u8mS++aUOrIGdH/suiGYdkuWPFDqVl18L1Ueuk/fg38KEckClYuvm
8A7WhYQmIC13TXPb6+LDRsnylp1PdJ7+O+I8dEg9YIid1qfQmRE9kczz8ix8yGHCW0EET3CMCyNI
R3QJaZlkRUCchTSOZrYNyl61C0aLO8ZnGLsw46FI+lVw0aOnMP8Nood1yC9pkPoEZU1UU8vkGLNu
e47RdoJ8A/6k3op89+681APSPKa5K3pvqKiYhIgNYCsaAAS74MaflHRP3q9gitaogRfgYTeOhhae
Ulfsx3xOnlSlAIwFSunwuTGV60T+MUPWh4dvaOXKGTaUQBRskEFUTktDJaGsC1Wcwua+e8AhQ1eq
klfhjEHH+M+F3MdhhenyQMR69Yn5UqIgnWu13obRkYDsdK+jfShMfwln5IUxmWcPZe6r7AwG7FOy
QpmgWQJAHsCIFT3B0R3ZHHifg3mTAWz6obR0J6OnYi/g+meTHAeTPdE/fFao+GucdguzcFsVSdIv
m1fdD54n5iwJORD55jGWU6wixTONifS9bZ26ff8A8o/v699KJkG1E1em+eNECN991jlSi1oFim20
W78nJtn7di0TRTDegAj9VuyqYCRnOLtuyokt2HHmgpkITDxdOFst02Z+T+MvafN0O+xE675Xf1I0
uNW87Fx6PF5w20N9oRylBMrprtxxju4hr5F0aOMphPR2u92h7R2ZfiyGbRPtaLTFOiZZPVGbNzU3
g3m8CQF93P729IiEP9jl2PgQ35Gbft5SlPLlY7NPVWLsF4PJ6P3Nvg3eBS3ik3QIbWiLQHUS1Shm
PgZ4xX2omiYy6xJZdDUzhKkfmRokV3krzikHdrOB2afCWBXkhk33f9SS3Gpwk9l95yfKpsuhqcEC
PVbFcU7HCSFFZrHkclilvgevdWKRat/OqdJ8Fi4weNWs6Au7sdAgIxkXeN8hDh+hvWQNntQjDmIh
D50oetWJ6fmmidZcPW2cceYkt/1ozC30tFNfkS1OXdz+WDj5XwuU0jcF/0obKWxzyOSCQ2MRoInC
8sdHXod2yTt4ARxgUXqodAj8jz3iA3+mIJaqY/pK0BA3xMFa6S8Bliej/KDVl/vyb29A/S6ZuOVR
1BM2llddKHHdViNeIhfqfjQemYBR8vQDJ4MA+dl0OaN707GWimflTHB1iaiZ2V06UJ8Gf7lN5/CF
w49i3/w4RqnlwHZkIebvFiZ6RaND+pWch/rrUuIlgsyc7k+YFDZe2/PE+3qE8tlGUQcXyD+d9vz7
c5fuhvU95sN2pkrf/g2vWSr8GEVy5m0WWMjUUaoe6d+fLq5bR4PiwvxDEGbYaDBEsgn4b3jJ93Fl
9kxAXJdWus7704S84xcwNdFWfS4CzUMJQuPGWCVv0aoSLiNeu+vM10hUukIG5lxC+8aH5UEz+kud
J17OHMbc9hsH9kHefC6qXJZ4Be1xwA0pigij21rzK4m6U6Eaj5nDIxRqSrynAwT8hDjKZI9Wpb2O
xdRL+cmdUg5u1B6Sz4jGU2ajwtUgVtJ2KUL+vmlWImqxa+rT/ae6WNUhGyW3wNgxZQz3N//7y+Cf
s2FhnO17kPuoCaretR722epvhvhni4h0v8aij2MF3BR7yVOqqb6Toa5lUW/pHzocyip/fe15QUXc
4TNKRgIXzdGXYoW5m7986Kdg9FVD8WADLOOFxw90Ga34Ez0yGbmLIowOjt/kqPQ9Q4eoVvgP+Xio
X/5NKixYmouYEjMHD1gD+ObVHRFN/hrSZSrbFZah+naVvpwjL1lwAIRhcks9aAmwnJ9f+mY3fXjM
OeUT2TcaaOFZIOEnK+pFO3PhYxWUUQJ9KiFK78Gyd39ftIfvwq0Fd/sx5SV+4HL8EvK70TBPN2qC
SbLTDt1Emu32RWxjpPZ0Sk16UOTiTvU3NN1YaQq5ylpA1eE1GE/loMK05h/OKsQ5jJfgjWIsHPRL
96LIPgXGj8Fqo8XAEEbHCnEiuiXiKA7KDF/7INJTr1gABUrSjBxC6hRHrN5jZyM5lxuhCtyv8VmE
pVDSzH7kn4k+aHVhzf8YiIiTWP++nC0GVyguzMwdvkGHi02q7FA7s46jh3B6Up3zUZaLHrxy6PT2
yIqREjT+3SCOV7wbwIGkMbjAaCHtH5p1VezmPpyPQ0UI+jN705whGTvwHQ1xYeS1Yp3BhQWeonVv
Dqg75Fp1f2h2GiHV4D2G4zxoPWhomyVLeMjB67i1givsh1PoVsejiKv2il90v34LVGok4SauAYkJ
7HBncez0/RdHeZQWoZd3d0tY5vCXwQnx9cI8QHYXWl5mBrdH5ZEFk2Kg6x0Z3zgjXuORicgYTRVb
DKJyx4gc31SKD3D7oMZrJRuzCXjMoWMMuwv9g6qn3vIjzEr+vzLR/Vc+c1kemNzyHY2sWNfphyYx
sI+Etp2wscu5B3STie5FWi+kly4Fpl6dtthXxNsKeza+3Dv3k4k/vaEBh+I/XYqSq+FROg6xC6qE
ONg33M8Wg46f2EjhgwNfbxIdp5CBnjywnNKecC+gXWO+NP0wo24pLGEJyif865kQM4TeNStmiqmM
epJvrsJTQjeN07ESroYA9rzZMYDjPVf9Leoj14FCvRtZY875k9pBArNdKtBUzhZ1UgInlpRlGcg0
7EgUBK2QGQ9cRqv7dYGQ1LTCMIcNl9sakouLjKXJs3PNVXIwzbmh5hYE+OqfmaFGpHtB5Mbv9or9
qAd8ajQceSEcjWEuvDpM7874cjQPFBXvrL3Y7lebHh8IP3+n9dXeM3gJEHko6g5FX4Q3Ev5YO/N6
MKAij45BwM8E9TLC0Kr7xvR/FsdcVrzqPd3Hc5TXMJjw+3OKP0r8d8EeK2ND2kluyco9IpQiZfpo
jvEBrEY/s+kIgsd45qlt/IXMFd34plnDvXsewoUHkEBEvI8F2OeODeCzJbYVsb7+XcRgxFwpLk04
5bk26jYzYCSFOmf5S4vZAU+7v0PJzyW/OqEUSXWFrHzwmaqLAFRzsLgwaDQEtxAUhLcD/2c2skl/
zD9IQE4aImJV73CXK4r7oY57PxyjBMIlul/5bg1Ltwe4llkbOBblEN7sXeYoaMq5nT4xbi29np6d
fxFq8h4tqApT7u/i9ANsnqlqDN9dtUeJDRZiVHfFvvykg00739zubs3ITBiFIrXBYqbmlJNm66z7
6XzR/CTjFXcVD2FLbtHs9TlpHvdvXPjA7zF0gwAz0JQS5cgFKJmMd0U+SkHPkl8vld8uEYpgFJcy
gPv7cIRiArueG3jl6PhJk1okZz0owTJWgOR13O5K57sxYp+6Trf7NBp0Ngujg7KdJTjoYN247N2z
Af4EgDhzLxUucm1lC5GAKwBMDp4y0IsU7c8PWiYKjq9H4BCdqRtcldTzLiTqacY0kvBivZUwxedV
3osDWvjnWhOHVlRDGru9dnD41r0J2Z75aDC/e8E9lcuRZvP+rkeotyHaWI2g2NA0vvy/7Qs632TV
o8b9KDczWTyRZKjEOGqKUa/Furluyvj8qyEz4pE5t5K4hr62+DfN+ELAvWt5OMNpeqbmJ0vUjj8W
lGvuYiwZSRI97/mmcM+eBN8sG8vDVC6YYAXRRZ3nDzZRp9hbjownMqSvJaQbD9y0mC7NBvCAfozJ
GqzQZR8ybXR65NNsQRuBRV9SroJ6bQsEVDHwRZIJptNJl+nq9mx98lH0RGxyn853jl5F7jfuHa/m
CL34jU1F+Al46rAIfV73i0309fGGu/II4pZJ/NyciMmlxW+h2Mj/Q1BFb4jgtVFKt/ZrO8mnxPyz
A7oriJ6dh6t9uPE9VP6OVcuSLxkzEqQU49QfXsT8ZtwMRQPeWj93hSzgZcbiVtjzPK9wTW/L7GKk
Ge1BQn7j7YbrJnJhjUD0sWztZWwu57lUz56PW2MTUeY2dqdbr5ZMQsjtTO+Cv2HETrT91VBTBUSk
F9ySYIVwLbyQ+gMRFkrj20V+JHmUQl8Sw8SxPfM3FMTqHSM8ioYLOrHqVnSZiJ5T8yv41RY9rmTW
cbIMWM8IdSDKYIDht08KruWWPsR+AmPJMUzlkMc34/DDCBmtNGmhEFp/UYpNxlzRBheYlrORIwv9
k7hWhqYYtm5BjplMRM2Khdmr5+Qxn9zFU4MsQVZ7n+7sUWQ6BWe+HzvMjWdzs4R6PgNS5YAdzTuB
tK+LFVzqU/MNsG07QHEDDxSF3uOHOZBAQn1MXvupic+oeePtebvbYlQAcgH6WnmjclifYhAR6MVM
AGss3Tqm9T2La/GhmMLBSV4H46UNOwsoQSLlHuQpRknrkQVxn0bw0Su1fXuJvIk02xLp/Y2QesO4
LXaPG8w37taIwQsYH9QTAPOS5RkECXgdWZgzaawUxVo2KYR03wVvEzdyk1A+GlNFfxat3M+PpHf0
3DDZj1nNiF1YKQNx4Kau4dAa9Ky6eZcB2C06wREgiGA4IpsWnsGP4mreyB5jOq17lcTSGdqXYNCC
Qo+CoS681U/euu02SaZlenX6o9uzp43Fv6b6Qd4yOMzmJkSDjB43KWyNuFEC6DUt546B+JtjaWWa
02kZiBHEP6PXqUMofmn6gsx266NXdymxS453QhHON5TDwryyHo1joruS66fMH5XVPnnNuKZpjfs0
ggKJF6SaOOA1IaVgboa6eb/T85BlUdSAPa7ZxM71e/KcEZLauqdmliMLtcbg5eKGgMxp3SOU86g4
LAAfn1e26gNbtw7Xrach2JG1khzEorAsQ/l7dqUKW+t8JrynLAoBz79qwHStpSmwTAYHVRS/auwD
Xm2S+yuf1ggeE128ypjDxUrrEKULhGbMtBPpGGu6Ato2kSzC/oSbMWybqdafoDbwxYsf0FKWwBdB
NBbtHRN9MRMyp6KtAZ59irYNjDpOAs+agtk+6tsTGXeZoJe1HG/BPGVNk1ybSf51yWEPkL8OzQwh
A3gl36s4AFMHXXekU1M1+247UuCURMRdrb2UYemDVebWoAIZrI3LeVw1COLqLuxsqq56H2UGNRa5
FCxu9nQ0JV0fJov3/I03k1rHuQxO5ghPg9m7Yhr+pDGJbj7NIInFocbcTxJKlaSPXXXnrYE4Jnpc
SrbBPCIUvHs5Cdyqt4JDcp5ZngPRkKnHD3QPWXti0cTnYV9RVWqFcde9Q3TEWb1Kwzh9CpS/hoQv
kBQ9h77ckCkrFnrvZHnVTqa7jU8egPUmlqZjsN4JYVFvqsy756ZRtxPgnAXilkA+0NQsAWAVY4iE
nBzCHH6704hxzQjW5mmxz1rRpcQsslXPeh7W22zkFXkXXv2KRrnZAtErto/9HKrE59+k7sbDl9Jb
he/QXao+f3NiKXyRCcYWizEebNV8/+KOSynw+i6FNXK+HC8qGhvN3T7qm+Xvbbptt14+K8TLa5Zs
WZLV9gVLcegVGl9mdhy7Y6umDvpaHPA6gFxpMdWRClSp6/wMxg48xpv/Ji47tAxM3QbjkbbbovE8
7RgENWQ9+FL0gDDmQkagxxJ4B1o3lEyqBX9eIgIRurZXaM0E/+B1iwilNIMUHQQwZpIOutb0n/R1
eAU3KCdHjnAkNeDkl9VzZ90otFKNpGAVa7WjTHpU3ebvwNaVvbm1LIUljACz1IUcOQhqkBuA6HvU
26TAU+dCGyvwqxo9FFAVZx3r4ZUnVm+OEq7G7IXKoM+iGOKTJ4r1sHWLrTQ6PFsSh9AzVM69+yxr
o6CZnbARtAfB/Eq5uFbP21njCm7UMKkm4P1Mzycep2pVC1lpOYT4T71oeFrfBIMrAydY17jf19ZX
X7E/5+/NxVM86MAWNozgnf+BJb5LQzoQTwOF6wdGRRhkYsMCqNvHN0jjTh42L98dQOstrJa/MBuN
bv9QDmb5WbTikbZkin2o28oUp42OURhQFf9LnIrAeTUxrx8AxUXrcluCsGKhsd2btbM4dEo2Hbpr
pMWbevp/bqLRmAAsAO8jPd75mLoyPeetW7bx8fUhOfd+d1Eq9KYPIgoWsLpdt45A9soqOf9sLARS
/pE0imSdObSJ+m8qAxg/fWUR56LJwSypSrNjOoFnPJR6bNfQmbUnn2LgMLJlblJ2U/L8fNqOAY93
WVrmjkXzRXWj8ksu47ymwH0l/Nyktuyl7weZ6PahjyV8vtq314CaJ18qGPdpiaAYtwwtYNdPErSp
SZXgeWmcgd/OYUNklIjmi1aEWRgOl174mf+MYL2zFvVXs0MiB4Ln1UNEGWyBCOuQTgZ6OVtX4LYt
GHAr/nzXuOeJyD3RieQRUphTeswqzklLZInKq/BPOHF7l0JVygqQrIBgMJEft6kGLljoYqSzYQ15
cV8HTkepKUxrXtYDnf2lpMgOIK8qeh/IWTYSRIbPAKid4mbobHy5PGIJyUvYID7xjJm9PskaxIL0
T/1ziW/bkx3jgoXPwBuDvb7nNj1wT9u0rLsLq/V1unkFRlV9TIEWeSA6lUHtYrsRKLNRzTg0ct1y
oHu+y5RdnIwfCzz/weQUimQtfYhiokQA18MKSVFH7P+OuC95Tx5mZlGekskozuri6y0ONqB4k2mW
4NqMCYxmymwj8cnZbDdPDsIwBpf2BXaQlZmy5evK+7LzCb5sjaClB822dzu37wSVQw1znb+C1n9j
KZyykexILPDc4YO7AsX3d+coLjug4JLFo18RAWQO102gJKch1yW31/y8AYgnsYT+zBFWrzVnc9HC
mz9dWRspah0EOyGBSTjONCVkUEMLsD8WGVzu0n3O9cb/aK1q1WsMM0AyY1LAyZ5MLs5XHC17MNIE
nDEEcAV79Qp2iqF5ffJdBMuLTwpY1hO3AoKChX7YeIG77nRcrOcjQo+v8hY016c1iPraHXsPN8i5
6Gzka+Yt7+vXZ6jKa2qgdjlZj5KYKWJXPbPM3rK4+TzEz1ix5HkDIHGg9E/bSe4F8rj9jv8vyrql
094oFaa2ZCln7MxLYdVqwBqecRbLhC5o2ek1/qykzHBQRQ37/tJgvTklFVyeN1wQVNoHtztXuFS2
qYcVD8El1DtzgVjbRhdoX9+dPPAQ1nPf/MTmW0Zv9SyWzE86Bx+JfC1WdQxxQzq20k2FZGtJthVt
AtVccpVZDzFzQ+4gRwT/+wKm61ezLJVCcVchnzEo6leSzupdc7JDgga9ZlXs9w8xhWhA85LdtC10
YYxoFYiLzMkCzlB2a9Wfl/sVATKT8M6Z1nitLOSLWT/vgze2JigqkrJ7lhWPDLiRj5bZJe8W+679
/34QgktJlQkzx+9qNE807ZqF7spAVC/n9WQfPrbE8LIE4Zpg0yQU8wrSRRnEVu5bUQS9u/FcxaxZ
RxvnEYQYLNO7u53/IFRdsgdBJDoG0iPuw/9D+WpdkutZSLj5kKzs9pjJNTWbDztRXLJgXwqvNxbt
1oXCoz9+ytj0Ll5bYqpqPlwYCHvbZAyiEktZdshEMFwLLV6hp7PZMaRcGAOWWZatn6K4/tk8ko6n
a9FSfxYG4VFSSpeCi/TaJXey4O9ruml/eQf7FoADtCxBnJ1n3LvLKK4chtdMW4ZTAm8NYrars3j1
dH6P8MnFKqBCAr68wtOivd9yW5WTY/79kuKLO6yPmIsyBC6yQPljqoeL6mLY5mz8Um9JSmLG+KTZ
A+JdqMS4aN1r1rLxQumBxONl+M2FR3Ztwrw4QFJd+MPmTV7CEEAoLVXbLL9Dj7ltFtIU+w+pQeGZ
aL4OUEBOZR/lPrC/CylzmqT80slHzcdVR/LFrXyZ7bkKIsRvhzuS49l3k5j12G4JBc3hV/Bxl3Cl
2wuF+4F2c8cqbYeC5//HOgR17UxugrszGf/YAO2+Dol0T6ViPsQYMLm2QwqUgdR1MXUC0vzC9sdD
ALNSzrM4s4Pem8x5QstlpJVCapQMUWvHVL1uKad/+BXpijErc49lnG9alyuYXyFXbC+Ab9mugU+H
efH5tDfia/XgLjGwlgtb2KV5RdQ2AOoNdC1Q6LYOMulO9g4EIpuShUo22SMKLoYQVi/IBO+RltEX
354HmF3MuB+uUJzc3b0YmMGFhPjGtU++ejyQqpBh1b8JnUInIwJ/DBi2wKMzQX5+63RSWWxLZkKY
KnQGSJ5SwlMhBpaW3xYKxRRiO8mZFdRgV3+znEaSyS6q6r2Aeo7amgQvqNNIw2PSYCqmt0pcmQrN
tOOK5QLKJNyQcS9mVkRf7RWs2oibyVUfCA+bXe/N3YSokma5x9Fi8JG5TTRUD/n/PbS7HR8r4Xmj
K1y1zpSXCBX0E3WgRIChIPOkTikQCWHOBPrnOczXqIVQCfPMv1ws1tKEMPYKbyQ3yMbZIEyxbBPX
nUF3JW7dy+YqB7UFLcEJH38tsyiyNqL5tpdjOVnrcIcyaxu2wnzLPEwosQ9dbY8DVW3Gp7NLqymX
6/E/leumMS37xktjuITUpLJhu+Ecxg86en6GLfbd+Z9q17AwxlDbem+SFY1f6S1DkVeN/RNLeT/I
IKz19pN4F/YjXabwrIAFZUdc6ibUi04Zo80iMMEZtpVNvp7pq37kpGO7/gsbFiPrRY0VCPeZqdOf
oeyPZjOQoMe1BrUg66Uu0uOUzMogvTcrj3qC1GIy7r9MF5stUSooue9MnHy9i3XouLqFGY5xpLzz
wxSoCQB5NxeDTq4Ek5scib1UMlERggspz1/dNR+ZqDhefQFpZG1/9RefLh2T3lOIn/uluUDvnZ0K
Ej1E16+40elOg8wrlf46TDNn2LpRSUt9pZONymQQQoo87/OqXwE+vRlbXUxtEk29xeamn3tEayed
/JBn1wMxF94R0SOzz1/5eBdhumeEOO1vdWnaBJRke9izRcEzfOj+fKXQ2TwLrYHUB2c+p2Q3SaFk
uXL302P0Qs8kiGUTaBRb5/L5v/CohCgl3rujgMl3KbeaF5ylD+0hHBoyE3RxBfEEVttsnw3XYkaq
q5IpYhgd5aqNhzTqNwATT+7Af67JI+wd0Z+z9x8Pzufbc626+s17ll8OuHsjVX85rfHKXLj0ZF+e
lQnELMploQuEc3zH8fQ2jMmdjYdfJBfM6i1hewLR2gTBlXhcflpcaHahRlcLl+YWSQUwS6aO4RF0
TNY/Tc1N4/33gbN7hBtkltpE/WvMruWlePCgBmDNDd3z7/TKrcbV5kO+dtOfE0tq5fBn2dxeGPLY
Lpk+os/PaDm/QwP/nbCbSgoxCKo9ji4ZQpQTT5D7MADcGVG+cVEVBLzS3NFwQ0Y1/G69n5ddVOdy
8RYUIupMOP9kEZhKLFWJau8NM9Q4+I6p9UoR1g/qpHNPUAY7VHBzVH5z4oAqINk44bSLE68jQ8JC
xu63rMR0VY3OE4GzFfvw+blegmIeDRYX5bJ7X8IFQkIormUtg4nExoqE6radZ5mI6eeI4oYn1d7Q
KevSK6+ymsyIzKkIi9wSK/UnC6EufWzkGrGAJ2Qd3Rk7odk8RNT5VxOZztNgYgzsRuX+7VHYI6L/
5C1YTg3xumja+IfJyJ2HN3ghP6x1FgGKRGeyxwQjXjAMQ3ptkAZV4XSip20CR3kaRFn1LiCIE2rD
XhzAjXvknAiIdy6DqDvfSlp6W3LafSR7dt+IKDCqqH4RBCZWr9b0bRJy9NMeggOL80DTW1MdQ0WO
mjT5yxmXBZ9QS5vbme4AHRCYuc+gg9dDYjZkwqlompdd7SEskO1UoQjKEx3O8KsX7OQc/xHMnhjp
Bkd1jFICWHS7qi4e7UdS1YvTBZGeedLEIt5sPdYDvU3Mg030evnJe/GQQ10ZA4+L5Qh1YDr0H0b+
foPPiyDUsaP8+1DbzwPKpGyA01W9InPcCmtOcwHvr3UiYNgjAdkld0i1p2jRHXlUt3cg2Ft8IoHJ
sXe24P7fqQjXszvZ20N0bL3Myb0Rif+SexWJVq+nX/yHUlrmyORWnSErLqZA0nF8qSL72N+Dl+82
CZWOHEPtQnTy8tPdO+570dfUx84V24M9JXMtR9Z0C6Qf4ui/heG0XmH1Zup4eQv0itOONMsj2evR
CHWoD3svcDpBQxrz6gumWkH9Orn/dfMbA8cotRDIIkZpoSmFI0bkY3mh0gF/GoSWjp5N0VgBjHD7
qhec6THxfIysZ56f6Pj2d/UGzM+iuXAQyAk3LbyprMWLFjq0htFmb9A9yP9Baxhiod1Qs/Iy7niU
xx2yOrjplAzggwapLB09Y1//fNsdtYXclYu7JHbdVBhHWohCksYx/fk2+S7g8G9kLWZ+2oaBrcWh
Ao5iBsie4jaxFvKluE9AYDfC0ixYkJP3d7uUL6iLJouqVdRte6m1oCVL/Kd4nmKiJYuehSnUJrnm
j7qr2r9NNorLSrqUMteJridAne10iqjtMxe6Z8T0oTrD7zA5GVuPC7PlvJ9Bg0rfouIfMZqelitG
aYGPIlZIN8Zr3NEWl0t6iNReaEruiME8efJDElvPpK6c/yxI4W5Au89RXacVO30oXtA6pa4fjDtF
+PJMt3+O1StE28wlFiY7KKdqhBsMhoBunYmqO3sR01j0mlZJcN1T2yqdlXtLoJbYTPMVAKMQ+/nc
9wmH87DaT2GUCFOmGTVybq7Vu+C/nD9eV2yTDTlaThSyha1vEozeR8S3PgC9JgEjbMBzYqF2gFYS
hOWK46Z+YfFpvnK+lj+oo+18KAmIYUN8bQKsTrn8UZl5rXktz8CYTJIRiDq/NveBLSBAH8z4l4RP
Du00bTYhZszZk+xPsKZ6oc43eVB/awyLrbdUDUDlpeAVjTjTSOWTGr4P1Y/dNp9JDprZtZ9WXlMb
5SyD5aY15xsNoZsPpmxVKjaFdjEBZteBnq3L8aGkjy4S/35Pc5cQa7ZyVjPmHNqzXg590V/GQg7b
ZCbgWZTa1x728juMPNLLZnZzgcGQjGh3ovcLH0QgrfDPl74h5tyNRUqhMexEozxoela5kSe+XJgy
ANjC+6RuSqYZT+mWHx/s8h/wxro8Z7y+SCGK1k97j8UN3/LBznBKMhKIkruAcOD0Pr4UApF8K1J9
aFE7PLFOnO9BnHlY+TIvokyG0levpQlTVswWrygIvPAn9I6uiUs5AWod4hroCVt4J/onwaqqJVYw
9MHgnLjEoC3Zbann4ajcxarY1jemitF6L8vbhdr13WHK9Q3E5pOXiscVRH7kjMdrRjcxRpSxaywW
NPxeGsv4eIZpcOhd5890Ew5YcXXO6NIXDDETNyWLZeHUrL5ooDhfT+EYORvuRkmOqpDtPDWVsegt
/8N7aQoDf5gLbo7lbS6g/7tFmaIyibR7ls1VPyIAnqr1L9vfw8reNBWBxdoYMv4hzq+WCFDgY57p
ulyVnQnDKJmAAqfsVN+/LyHE7c1+lDvI9146KzRpdfiaAg2AcnPQWWdjdvH4VgiqUaIiKXVISjdE
N90RViuf5N/04nFkkep7+2oscvbuMrDW8rgRslWlwvftOYoRxl48jRY9xQ4x8v3a4Y4ov1/HaeZD
SuEocBIG3Qjn1F1BhJWwF6n+MCScFkA+iYgiKoXrRWC+2Yvhnpm0UqqmzzryoGIPd5EqwH3P9xUf
VKrIs4385eJYrb5piJVUWeB0YjOy5CZIHS8787tYxY+saecPeXNkJObsUbfuESuz7lNFrLOOt495
zY83XaDPtGhpxti/8OS6Ax0E1Kb5JLTOUmRECb91R6mV5DMv9HfEqXH4rOElgoNtFTqqDn87gxzg
ydIwnBIrcNeTDy+QFWCzRMGICujBRseXSPvaUrcISUO+kZNGnyOBttLO7rBEZYbTWPh6YD2u+jKZ
uc1gti0tSl+xWtvEPwxEM21SCxmnDy83vofcHbKW9GIuPQcM2eViV/VoEJyu6B7L8U8UyQwIXoqJ
B3F/3N1Lpcs+AbG3nqZlsG7J4yKYN1ib3SBukp3+GDvQgkx4VCKjU3TlQHPfUXlXST+fqlXFyRv0
IleFBpKBItFbGbvmpw0l2oj18bm7lv0+a3Q5POFYM6nRvtMc9HCwnUoApqUvE3ZHkCkmSKt37e11
qEXuIXWKF98HzluIYGf+scyeeNtawAVVH5kr8aF0IA0kt8MDSSEFGB9tu5WBCfsLtg0RhEp/uufA
viuCzfgLUCxxO9rNv86hFF1rNc+GOWgvy+WstW7cnul9wcFVgcsnnwIBwmf6GcbmTYnrgqaofuIZ
sLie+J46TY6KToRlxB/xT1BTQ/qCEenT9B+o3L9wp3ePKEJ+t2LltujakamKZy5rYMBYgQS2a7d/
bOwVb4GSvjH1siCMX0wYAWE/NJzcsQDBQcjpTDkTiKUCDyEck9J/7ZHxRO37Ihm5cSYQqFNLWhlH
B+Lrg7lVTg5H47qTtpKFRvm3ZKHeAqF6fqu43zUekuUxaLbkiCer4pTYn+++FVzH2YJ63YVmW/r+
Rsm8H7NqlXpxdnVdcHHYrwKu9fehyhO4QhXABoRPhlFhdlaHeTdtLCnDWA3YX/I/Ik5l3iWDp7pa
BUQliEHBs194ykwIZ1X4WZB97IyYt//pNCP4PzTml5+86E91Nn+98qHSXm52HeDcEKfO8p6g2XHd
HTw3moSP4MHWgWMJ8oCiyQy0WDlIqWdjVWrnlOPKuOmWxDKnq4egugQ6oqxkN0FeJUM8go7H9eJM
FPt6EvslHrjkqpRHuB+koghlPZk9q7pct81MuAXelkCwJP6gv/byIYLRDTOemhB8CB1TTKC7xdLC
MmBwNlbHQTe2IUNm6uH7b2E3ISmwMttoRzmR7662gVUGG/Z6UgKB2653vqKfpcTpDanCG1VlnVRf
taKfFnKxQsxjigf5BSSY3Opo6T8ENxlfNdxCxa7tHy4Jvfy1b+CIckqoju9fICHp45P2gZ/uMwTX
7Blb0YZRUs3hYgyXsqpKvKSnr34HexAcMKTYFkO5CK5aljyncQbJqoKwmEUX8JqouQBIhxshX7bO
N6FDMHc2CofW9mfXd/PuooeULQ9XR9GM9GsHbkTcdIW20JlAzTTqJCoMBzoyB2BLP+eBTdMnIKtB
M+ABaSbfQkczFvfwrfPFbo2Pukooy1sK9oz3h0hjTVclskjqgOuM+rqL9MvXbJ2fOw5+IUcvGQ3Y
bPBYg+6xj0wPGSOfcMrbT3NE2kzE2BIoJfahtEnWVWKgcjZk/iUCaniVdOO0jSiG/yHySQUbxY1H
op9XVElahOm7gDs40Xd6oVjL/nlzhAJiIKT0+Iw/TFkg7W2SkRSlVhuc2OS1syeD5/e24etLibWq
HLs4sPxOQ7byOfkB/e4jD3gqPdckoOG0KN5JcmuJKUL4rXVvhjDLK5jXYFiniOwxVqx96K9qbr/V
omLaWN/6Ffthuo5qc4wmA/VRygnlSuCbaKFYKUrXgXdoPzccbWXWYf9V9u0JTrgTxq4dmjlw3pSj
U8yZwXYpl0h4B2Bcxi4DRx1o2QdTRGE0YNEnIMoXAVLmyZ+kuV1yNj0KrWAx5N1P85vjLR2uYXhO
1sx/nHBGNja2VCOy8N5We3BbK2Qifci2Jta3JL82J4osxt8sPhHjJHq6nqs5cJke/px+MX/OtGj1
sFJUlIz1Ypgfl3qkjPZMiGD0mqHjsrr+mEeamjmJPK1HSzmnH3Hm1jAOpYyusEB1dFOEvUMvm0HJ
Z2e1CaiAuy0uc3p8RS5OxPYjbzqmwk4ylnO3EwpDEW1YXTFBHXfVR27AD9scULVAy4lR785Q8GPI
vdp6SebUFjZK5RgMM+9HjvPfV9r2L+YZF81W0aayDUtUDJWz67HVdUlfv3ID62MTbDwSrNJkamLx
kBBbDxqmloBt8pFC9mkZzK1RkREe2b2HmV+Xpk9Ih29M2Q5+ejESiEy9nFwOeWQw0VhlhYFpqOgx
3NS0G2dNO1ogSXNyjqaSqpnEwCkpk4YDgXr1DZH3EzxEzBYfnkuawRCby/mKpICw9BWNnEMySO00
SrZaf68f8+/cAFL5nx8ymFPEg3qt81ktDFj+3qHbYMa3Bp+M7DwCclq8b/pGSIy5kIyyXXHjxugn
eDgaBQGwrfE7kzBg959S2ZLj72yGqPcEgeUamAb5TtKIvFDTwUbxtADjptDTNhVwy1OsdOYtFJF+
w6VA4cUBREvlR2I7XX0Bq8fshxJ4HRoToRriemX9Gtv6b27HPc1RR/9E9X3QGB0U+tXFAQrW9ndy
NVq+In/jim3BWGKRCCRjKcdWQDU3e6WPz3fr2CY6rFlaNmNSAXjaZPQLicLFvitG3nPfy/ysUqC1
L06eLTOgKt1VLfl8sQnbVQhn9nmQC0cus0Qobwl+/w9RxIq46LSVjD0QK8vbC8Zuipt7iteOlrYm
ElXS1pZ+VJiEd/efe6bNE42UKOiwBIhNszDhyFplCIDkvjBLuN6+kQGFrxAuvHotrUHnixuw9xT9
T/YLD4+P9q/AR6Y+MF8uJN2ihBp0XiK8VFTURD1kjkHVCsZFGbUPnoUcIjK46CnAnogTk+UiX6mQ
LVpBHiZ18e6D9+qjWr/OexU3V8dk+2MW8pJOySJyhoiza30S8wc989Lrdb4U/vmFCQr/Nd2tSQ8L
ERe3i/fc/opwzC/fpcz2J3zB7F6+cYNcIdd1nivSl0bhO3xBosjPn6YE9zTGx9BB7PFJBJdd+DXS
pGloqiqmy9shB+vKuRJ/v7JVoRWsSUy22rijStAzlTwVvSe3+Y+5q65ycmYlb4l7+0i/WeIZXM38
HDJniLpYNIYQN9URZ3EVSqqxKjzjZaiPHHif0iaM5OMfmKSyeIMnWcHuh/nkZy2TbcXg3yVG58tF
/di7pWBICdYfi/5TF9IWMERwL3WQeHfSNAG+UhFUyJwaIRamFZzpl4RHOjSCCpSGSrQWxIIH8gCc
qHDncYRBLjmWc8r32ojErZKaHTK2xNJ2oKQyBfXpTFZIahgtTwuVtIdndLOJ5hxSVPUHlCZURHEF
YxVAxLGiOGjUqkncr8Bps/X84cO5Q+XPlWjSkh2xm3jdk/LdFleaeQbjrBjmZDrPhZx9I/7Nm1+l
FyImCa06/D5IoRNyhNZBGDdM3uaTvdroupZyZYdeB9sHB7fObhYIGN9MhhXYx+6I5X/7QHPBH1GQ
etTGTooFjhGjwOA2JeTPFVEePx+gER0kQD97AG+FP9NUx90Ztt1VZkFtTx8OpOq6t+HbNdlHXpqZ
IqeeDGdATMTxOhC/P2JPM4cdsAMpVrvCMuwsQTZBKqVteRoDm8aDgO71MxtgszZex+QUPAFOcTDC
ficCPa9Xr77DXcY5lIO5sl4G50VPWQmVRau5dRLKEF1dEVDIStrc3y+yZqEIvErI2iEwp4DXH3a7
tE5y1bkdqr7a6pygw9fRYJ6oDTtsCwWS7gTRcbvvc4EFIqBpD6pk/lP5OT2vL5f0O3bxqYx3UIID
/z4KXZtXAAA3kNA+G8qFlpL61qEH4wJwF/wUTWJrbw0rBvJwI8FYhkvZI3Am8WNaUS24ebMrxmwj
zAIiSCN96CVU5r22ufAaiwT17fPmVxDzj4ZcK1ShNU4srgcpPIeedpTsffvjNG5QK2T/0cYUOToD
Ucpxa1QRG9p8ilYVuYffRIxnVnPLwLtVuBOxrUheCvgxd52sX1URAk6VdYAOIPN8r5vzCdnluPQI
5AtB30W5azsXf1EhmPt24mt/21LZDj3Nr7pCxbozgxypactAYV/g2XkMu/NAhh8JmApB6EEog7nq
ffjZ8Lxt5dgZ0wj7luRO/OLXVANPzNT3RepIopACXTicAJ5GlnoFJGJQHY0TlflisgQPCtzP3cQg
BE/wDiVA4Vi/0DUNikJndjoJ20k5PejdSqtgpQW/YeRitdg0xKG3t7nBnGP9hgt2R32734OrIPSG
AeEZoIXcMqXWzQ4gtcBRSK1DT2cdswAKzgOrn77RL+oDYf6OhPl0jvGGkgqt6S99mlkD5op5s9lW
RYeMPBPUpRaVpqFFnAHu3+na78ToN4AgxhRY5athKmYyyNOJvwWO/EFiolNwOm1DXUURAOQRvqv5
/xIS/syU6ph3OjERJGDgutCrAoUNuk8mShgd+em7FhDrEJvk1HRYXnBfGLQjvoZ7QvnF12g9ebJd
ckOibZGf3zbPJgP6I1mBhddGYRj9+jzcUWmQFgVJ8Nr84Pdm2iESLkx5QcwnCt7bBln23PHQ/IdO
gix+VOMvBcIT/3GJpG/lo/v3/n9EunJJaSMkvOAAcIQKwy7MeXgLfEMeaQf+SbF8uIqUAZw0UBdY
oKL5FpVnR8BbUNAUlGQt9q7FnwQJtM8+c/XgUjetHckrl4V2CrTRDaEnzv01GGxX9ND0YWNhbHmS
e9oIOpYwCZZ5eC0HNOr/hyLuOxquT/rgIGv0OWFbjGeGB7aet8h+yEnIi7KSxYNyg1z2CwmkNFrG
EK9BZT7p/s4iRkuRXRg9SLZ0x83BH21AqUr3NKKEcvqpC5RAw246EmY2HQ6kO6oM1dzNj9Qdfzmg
QIoN+posegYInMCsTrm+DBEmrrkgGRw9/Y4s1/cVU7RVwCSBBrGSsol4YyZ/YFiHJHnraplhMLXv
hJhF+FcGm4NbpEozPj6RTOSxzXyHj9FFNk2tE9lIbEdLMt+vXh9GYZr/jS6iXLqgY7NL3MbVNnGD
KDuByD6z5DRThRZvFV/Aiwvhw5YoVQ6Ufi1lRpdQYq735bJjU506lK/s8TvfI+GJrNrbbow/FH2D
vbU20rHxK/pjghSyV6DhHr6LpqEcLRcI1A13HJNCfAcdXAOeW0Sdn8/fey/ofLEqj5pgLTRiqWWS
3/1OmVyzyyv2zaeLDngnA/E5xCQ7ZdssKKnwSCWq6dXHHyvIwvwGiIu4ppPlk2meIzrG7PVz3AEc
H6Yscf1u0gT6G7wEHbzr02CiwDxK/ppkY8d/3FIzxqjRDR0OeQ64KmZRO12vv80EM1+uYKeRJPDZ
eWcmnrO8eJN+DCoUlOLsVCueaF0UQhaqQG6Gf6h7Eu59JKQfLegkZdYE+QN3cp4DaxUjPgdiYaK6
GLlb/bUb0FlqAA90oiiG73bKAI4L9RWKmiKp1RKzSLF0ibBdLfqd7tc6wc/PHfC+Swdn46POSazL
ixwaRXvtKEdCyGTISyR6xcozqi4GsArGan3yaYPpGLKRPUTR1S3JJuGyYXsMFPVNqCDz9m2yeX/d
+lOZc6IPG7F7akn3Xk8TXo18f1DLgVbUW+YLnJZlfJcy94YXqY2b3rlB3GM5iLS4hj23q6xnyzTv
JYiCrotAY1HNNJl5GYnDFTVfhu5HkpgmPG/nnFKU5kvzLOERmRyfKaDA7nW6B/osYKq3nOpP2s4I
78OHjkAA+xlJmcVfMXQopH+w4ZqhrOFFQikPZU6CU/piYRfhqYXa9xow5/cNCfisZqSGWWYhLWvb
TODTHjKigmW3Qb6xuhCapnK8wtbHCQ0L4B7mAUBfYkJBZUMSLjf/FgP96XjOrZuDla5gpU7zVyAG
uIS2OVIyEJFhgoMU93RtCJccJSirYXTCudqJPu9iZPYeMTQmdOD+Rs7Av+KezvUOn4JjbLipkAVH
xZSjAqgFoybOBp+RYKA1hYVvpfNOLd6hRICYz+uqGxXgKHxAUt519cJRkXSJ4rojJAiR6/3kxTNK
Bs+jxvRUz+3rJW3yc2TUVqT13MigfZXPMLUQP5ASdS9v8MrhsbNSa9NOoofAmm8yZ1ZdefeIvtGd
bk/dYzOouH8nHtum6OMLuF9vUoopH8JfTPHsmbpKvYjdtSB9KAzz38dHijSC/WqGV16LHJeUyL4O
LeJO4hnEIZRI5Mv6V/NGKrqwgr4lE6wgQMW3/VCojIqFAadEzYEkMl1GcDfVgKE3fftErl53MKDj
FUfAlm0qBrMcQVpQOKEkMvNEXOYiw/yci3OD8Q319GIzXPk8D1eERKd+spxTSmbjh/gKUi2A+0BQ
brls2e0sZTE7zWO32DbkN1AvvVkEDFiJvAWl5LYPO4eZEjobmFZi5eb1wYRhn2/+NiCZN39XUpkK
kW4Xo7R/U6GXRS7Mrf+pEVmhcCmF55dy7otsCAzjaQ8xp8030ISqL6r38jfYYaB3WM638j+YexTj
JYNtq6XooF7QE4i1Nl3A7GaD4IDKyaPWEP33mScAIE/JG4F5/qmelvPSR34T9NGkoUCAFhBhM57J
RH12HZDmiTrKiQLmpXvHhVmYux+sNdffKbNC7aq8styIOvjCea0fpHB0Jv1halVqjHlSQeLlxojn
dMZgFDk2cMrPB+J15SJOqBCKc6/6EnMZqBR9UDfejzxguxoC9mdC9bT7aLH0ufRmebdLTYGa5QYL
aaPVCAysNYAYglhZg7vSV3sko2xdn6gpo3pgi2oiRcYRWfDouUswajS3qZj9oOUXkOAOWqyAUndR
B2HIhN0zWQb+zkbcqVSCG6M/xzKhF1jGYFJz0KXWwKqpwoVDPxwYdlzXiSTjCcJpgSevz+h/LxME
297e/On3xyBpbzga6elBICxKans4B7AkfKFygCaYUGQVyuWUL/8CvKbFKNy3Ro2CgWTfiQk4qs58
/jJ1gGDGMXjAUnNcLPraUEKqZ5DwOIfC0LywQuEDFP5ZaNIkQCuXJ9AN7ML3BsDg/joPb4Ll2TGT
ezK9/YKi6wyYERrAum/nbmra1kaPu9Op89DjTU4It3Y5CT5TufkFyh3xi+xmuw3VyfOhevq4IXAi
Tb72EBWj+3gsmrgJ8sBepU1VACCWoBipj/yyUPoTNSfUWiISJ/g4twnDCGlxnJ7oYsox0QoU8dtU
iMkcsgmY5TVA2iUGGVeFqfO8YZ3D8KmSfx+feJF7ADx8DmmL6QeIuBld2yJ8P+PyTScAXGcBsP9O
60LPeJ3e+5K6QYlP92pKUrrc5anv5lj0efwn7s/mpU37iqErFJ7sgzx4vQuJ/aYKjiuUznm3m2vt
WpQJFaKTAp6O780LyvzKfI/+A+1uedpv81tjwziyO/m1NfstsBKfLhC1LpV709Fd4u4md1FRqNX0
K3Rzh4cmZrHnlbYpLVWfTXi9/HFJbSWX3BUcSJTWgoj1WSwUHCwUqjbsQWBeo6cXx2II1+/v6++n
GmRfRFwOJa/600DaViVxECY7frVCItyyR2IdMTNtv6yNnOfzUbhZ4lF5rCR4Ga9ItoiDsS8dyKoN
sbL142rvoSw8OYvT8fi9Uh5YG0UHbuHPY3+qdPp1y6AuUB3zw5KQoQyFa2+n1bNrvEszTrY879lS
DDVXrWUxHsfCg5p3I0NWALime3IBBEf5tVE29Mo1lxqsfqqO4MMaWnLZDfY0hY9SitzSVpdB+Z07
HkQWVYd0DIZJHaAYW5kjRE3qqHKGqwJMq0t0dnWO1fNlWrrUaSn6wrwzHUZeCt/YimFkAadZJffb
EJk4U4ohDorbPlCQbHqsI8/xmweax0xEvG+bymuFCt6/3RTtMv26hfXw8V0YPL/+7by76tbyVrfM
VOBRipisaWwvL90rmm7C1If5HQlrQ0H1D338EFI+lIfQyvDrNlgx3eyM0pfe7WFUJxzN4WuBJhT0
CXdA9XW/cclPfaFSh/EXS8eHuG6pwsCwKhjlYL3LZkWJJ3G5l8gHLjXw+8S+348c/Hu7nmjeBSTn
Kkf299FmbrnCri1Mp8UewPdd4IJsj9EUITV1X3hOOlLk3JTj4ULZoxMQFgC74R8vI05dDVsyNBB2
asZup0m89AB+AO9Qgz9NOd/luBSL3tzzDIhKx3x67oi5vnp6+MXGC33fBPMZnOFwu30DFmo2vqdE
Mrf6AoqObHe/U7A1wGNTHgkQN1g5siRmkw6yhEn1q0mdI20gaLu7w29fI8uk2FJbhwzf6ywY5j+/
pyOmk/DRh5gug89a2cWwwVeoDCaZMtoEaLA1nrGA3Mqu7/uxjzuTWJiBGILA5F6YqrtwgCMxeJeP
CnbFXldPncfhPRFeTy8x+zUxPTACZ0uaLwsV5twxjKLFw11nadrK5M590RG/XPaOfzlNzT2Rj57M
2VJ6MxT7cfkUoEjrn0/htPTOlO1w25YK7V8w6I/XqVWikDRhqSMcoSkLsxkT4BNFOb+x8hgClE3k
srNzKfqgYzt/1BWLvaP5g6fXQI2zFKTdCccBqvv1C2YT/jcj4QXxTGYX1SVvLTl6NrmcPUMEZjo8
tQeWsNH4wtQE68+elIRpDU5Q5TGbKn/2gxN9Ztyj1ATu9A7nr/yErP3VATVA5x2iFXTB1O8+ZdAL
MzR7BAld3b/amZJSIdvpWtSzMlBN4HWDBq9BLwgBpOLbxHJADEBwn95OucvxObqaJfy7/X96jtPh
S2HSD64VM2pTA/gKkFSp3PDxTpkddsecEISG3+qU1ZvJ8z1VNbJpiOwyPqkVHBZMufrWhYS0vVY4
hrn/FmBBmSja+6/bDlc/Hcy++9oFwN2eG3Yywk7OlwBn1qMgCrnnq+bFtkJOdQHwWJp1apFjAqHd
nxokeVMmiMrtqtH0AAxeZNJ+KBjy6iEPgc3ingaPc7HeBi0kknQQbwJTHzEFyAGiPwqLRdpDeGbt
sC9EGgTvpQ6GsLZRZFfhobakzS49c/4BaeqEFbT+vBL4KEDzc+uqZD5ZXdM4R6OlzVKdJFMI5BaM
QLKF+Ksjssif345s8srFKZXkSFQKPsH4ReN8F9CyAc02cZ/cvatzkAhMOxRrg6dAnXjBIqVC6agb
9m9+SQlbyA7sg+xclf/W+V0y1YJ15P1F2fSn+GvgT0UAjEYX+Wnx9bUywSRXOMS8f6mq6rUscVgu
KFEV3/hozfb6jtSWpOYWItfiqJgYyRaOAYy8yqGcm7LKn9NxqSkUtu3/aBazZjtmjzm2xy7+ssPX
Wn7r1wFhs5skLfsQnaFc9EmL6MMYZly7N8yfWAJnOV4DELtGZaCFOB0UHcq7md2ooRY+hehSmXIU
N27D9NO1GSL62G+FQ1Irgp1gboLDwedIKY8VprXLCi6E95AN4SEx2nekHFuO8TxqTSdIPWnmCaaE
KLKHP3bIwyFMqA5p30WB2alkG5CVaV0QG6ijFjjwh5QnqjVUOh9dg6RHexqSWRCi2ojicEH5CjwN
G7ctl4G89GOY9MRL+rnfzpFm/NJhAHF1p5unOyvAdXkGp6wDkfffwoT1SAoHxiFYRplKX/uDIy1P
E4hX7OMknz/e9cOVXJ/ZzHQA8LVhgaci1Ms20l8Kw7oOartR8GZ1Zkj6tzBFcFLTdOtPEv67BBnY
tUoCwEetQirwnb+C4IrVQOmUizgARLnlUhwBZcuJBiqT5urx0MG0MBqUcQHsUbI5c/hCkhNZEQig
6W8GOvuv1JL5J8K8um0/7Q4Aq+C+GX1RpWolTNzn1H0At44YpZTed63zBVR22dhd1waAxkP28YPK
YDsNdiQNihEJU2ILjnmNGvMXGf97trjBWMTLfwJgENeNLNT7MiktaBVt+LhYltECJpyR32dQxJZG
XjXtQ114M0utLBf6Usek1y2weDgcX/wn4KMwtmV8B7VqVRgCTPJFvcfM0BQrAFk2GBEBRauyH1NN
3USOCiM26a2GojYqD5cPq7tGLL37npk4ZSxzHRrMrVyWI8eOFZGWU7IAQGEwp7Ih9U2/AdF2L7hk
AeX0ciK1G6/mq4ULmlZGBqxC0s6jhMa56awhGeLsw61XxSDQorDGB2k7/1bOeEYDOoR1qk6IHygP
GH5Pe3tyvEPp2vUZNv0C6JvXl+e2uDEVwNO681ieVS8QTbNvcDMNea7tU+C3pTwoFzQOxaml4e5b
iBv6aDnwoTzbfgdTgiiA+iWmxHPTlz92NlAGHyPHJv/uhC95A0HfPfHtja7Ogx19v52MtXvh/62F
YnQYaXzJsBy7AL+p88Vxg2PMc20kCEmLWUrhd4SIz2wKcKfUjfWdHKnvPb3ffGiTJqJ8CBaa/UIT
PpBroDD+59DanslJS5PQRCNxVLOh0K2qV9trGrLi95HKIMIB3id3eEr6LGB1zzSGI4glEEYC2nku
zAooHzb7h18jNmyQgYhDHVgiwxvmw+M0dFjaeKJw8+2CtYOSS/UuuAA3qw3214wye5amcS9GAZvw
TVF85y9DdJrdjL3FUFUMjZdxwckSc2dC8yP7jqSIRF8oSyq67YDeL0ryAaf1ISS2OdQZ6eU7w0Kt
pX+TPtlrYOLkdg0Rl0eTJ3IlVz7hTRmRdVaVPhDRVjfYXUNJEpUUfKg7PQYAVzdAZTA9W66tgg04
vP8yLWy/fRvc//buqXwgTfKmZPUvg2nW5APUP6VpZuNkfPiQptxRelCptwVNpC/tj/I8p64C+35S
vhjEwJ5zQbpW2CPtY4RcnMCtXAI4c7VXCU6gBq/fnar4bXgmyHCnrps7KWlVpHUIfRDsvJqLUkca
ARoHWDnuegQILi1vYxayN8BkPAnOwK6SMMMO8yAa/YXDVbx6BRqhjvr5aSAkrOmOo0yGINEO7CqF
NKXfN6d+V7nnCoswQRtFm/WOWEZzi3gsDELdRi3obFjEFf1rx6zKIpcFHEdcuVwCIhb3Wn41wzIn
uk71qeqPdOmvuKFHLBj1NW1qeT6Wmg1Sgbh8AyvE9DKLupVBJyJTtGwEzbK1jlkbToUd2V3OB2Te
27zuyW4KoKta+8T78d3DmFNfprFa7odK5yqthIS+yQXBd4laDR5mr+dPpSbfRSE74oG+Def0R8ov
yVcAPHvoqh3omT7ZjkBO6Be24sZBWejc5sBkSrfkVN/L5VEflOrEuY4APO1gAmbt049rIv0t6+qw
KWUoPGa1CRsToEA2yNnrvzAgRMWo49AASpuTFCAmfMpnl25s491PP+C7aT9kemBs6cONl28ss9CV
gZxZhjGaDqv5v/5IfOJHIaosIiW65oN1bD7xRre55EmUvBZrJXZ7YQ5WVXVW5iy4SzId5JgDRfLq
TxpaQiYbLZrZdgUg5C+oVYAyXrydNzTQmFsRbaJlHXESgViAVlCTAKUt2lm/PnSlAenusK4G/wR4
5Egq9yRFdFwXliDF+xgrVVMSoDbl2iIMxZY+J4zaXx77TlTiLIsK+S+DHxLovJCFcBqpU7fRUSFa
wn5N5+FBEn3Je58ZTV+lZtxvRa5crZRepm3lz9hy691gH9It384DUScvKYJO2Sk4TAFBIjDbjnoJ
stkO/J9fxlY1Qg3VDC59kRx7EWvJxBoyFIlqNhVomnaXonyBBBydKiMt7coT1JlI1Uy+p/cBcj0k
/qirOsqTNrjRvS3kjGq2ya+JSAuNjkd8akmRXVawfxsYeJjnmh7Ft3CxWjSkG0qihgvNcrk1br7G
uEuc06Dgx+h6ZGNzJCAJkgUjyo8J3fAQ/D/HX5CdUBcCQ3Rnko5biQw4Syn924xu9g==
`pragma protect end_protected
