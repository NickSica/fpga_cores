      output  [C_PROBE0_WIDTH-1:0]             probe0_out,
      output  [C_PROBE1_WIDTH-1:0]             probe1_out,
      output  [C_PROBE2_WIDTH-1:0]             probe2_out,
      output  [C_PROBE3_WIDTH-1:0]             probe3_out,
      output  [C_PROBE4_WIDTH-1:0]             probe4_out,
      output  [C_PROBE5_WIDTH-1:0]             probe5_out,
      output  [C_PROBE6_WIDTH-1:0]             probe6_out,
      output  [C_PROBE7_WIDTH-1:0]             probe7_out,
      output  [C_PROBE8_WIDTH-1:0]             probe8_out,
      output  [C_PROBE9_WIDTH-1:0]             probe9_out,
      output  [C_PROBE10_WIDTH-1:0]            probe10_out,
      output  [C_PROBE11_WIDTH-1:0]            probe11_out,
      output  [C_PROBE12_WIDTH-1:0]            probe12_out,
      output  [C_PROBE13_WIDTH-1:0]            probe13_out,
      output  [C_PROBE14_WIDTH-1:0]            probe14_out,
      output  [C_PROBE15_WIDTH-1:0]            probe15_out,
      output  [C_PROBE16_WIDTH-1:0]            probe16_out,
      output  [C_PROBE17_WIDTH-1:0]            probe17_out,
      output  [C_PROBE18_WIDTH-1:0]            probe18_out,
      output  [C_PROBE19_WIDTH-1:0]            probe19_out,
      output  [C_PROBE20_WIDTH-1:0]            probe20_out,
      output  [C_PROBE21_WIDTH-1:0]            probe21_out,
      output  [C_PROBE22_WIDTH-1:0]            probe22_out,
      output  [C_PROBE23_WIDTH-1:0]            probe23_out,
      output  [C_PROBE24_WIDTH-1:0]            probe24_out,
      output  [C_PROBE25_WIDTH-1:0]            probe25_out,
      output  [C_PROBE26_WIDTH-1:0]            probe26_out,
      output  [C_PROBE27_WIDTH-1:0]            probe27_out,
      output  [C_PROBE28_WIDTH-1:0]            probe28_out,
      output  [C_PROBE29_WIDTH-1:0]            probe29_out,
      output  [C_PROBE30_WIDTH-1:0]            probe30_out,
      output  [C_PROBE31_WIDTH-1:0]            probe31_out,
      output  [C_PROBE32_WIDTH-1:0]            probe32_out,
      output  [C_PROBE33_WIDTH-1:0]            probe33_out,
      output  [C_PROBE34_WIDTH-1:0]            probe34_out,
      output  [C_PROBE35_WIDTH-1:0]            probe35_out,
      output  [C_PROBE36_WIDTH-1:0]            probe36_out,
      output  [C_PROBE37_WIDTH-1:0]            probe37_out,
      output  [C_PROBE38_WIDTH-1:0]            probe38_out,
      output  [C_PROBE39_WIDTH-1:0]            probe39_out,
      output  [C_PROBE40_WIDTH-1:0]            probe40_out,
      output  [C_PROBE41_WIDTH-1:0]            probe41_out,
      output  [C_PROBE42_WIDTH-1:0]            probe42_out,
      output  [C_PROBE43_WIDTH-1:0]            probe43_out,
      output  [C_PROBE44_WIDTH-1:0]            probe44_out,
      output  [C_PROBE45_WIDTH-1:0]            probe45_out,
      output  [C_PROBE46_WIDTH-1:0]            probe46_out,
      output  [C_PROBE47_WIDTH-1:0]            probe47_out,
      output  [C_PROBE48_WIDTH-1:0]            probe48_out,
      output  [C_PROBE49_WIDTH-1:0]            probe49_out,
      output  [C_PROBE50_WIDTH-1:0]            probe50_out,
      output  [C_PROBE51_WIDTH-1:0]            probe51_out,
      output  [C_PROBE52_WIDTH-1:0]            probe52_out,
      output  [C_PROBE53_WIDTH-1:0]            probe53_out,
      output  [C_PROBE54_WIDTH-1:0]            probe54_out,
      output  [C_PROBE55_WIDTH-1:0]            probe55_out,
      output  [C_PROBE56_WIDTH-1:0]            probe56_out,
      output  [C_PROBE57_WIDTH-1:0]            probe57_out,
      output  [C_PROBE58_WIDTH-1:0]            probe58_out,
      output  [C_PROBE59_WIDTH-1:0]            probe59_out,
      output  [C_PROBE60_WIDTH-1:0]            probe60_out,
      output  [C_PROBE61_WIDTH-1:0]            probe61_out,
      output  [C_PROBE62_WIDTH-1:0]            probe62_out,
      output  [C_PROBE63_WIDTH-1:0]            probe63_out,
      output  [C_PROBE64_WIDTH-1:0]            probe64_out,
      output  [C_PROBE65_WIDTH-1:0]            probe65_out,
      output  [C_PROBE66_WIDTH-1:0]            probe66_out,
      output  [C_PROBE67_WIDTH-1:0]            probe67_out,
      output  [C_PROBE68_WIDTH-1:0]            probe68_out,
      output  [C_PROBE69_WIDTH-1:0]            probe69_out,
      output  [C_PROBE70_WIDTH-1:0]            probe70_out,
      output  [C_PROBE71_WIDTH-1:0]            probe71_out,
      output  [C_PROBE72_WIDTH-1:0]            probe72_out,
      output  [C_PROBE73_WIDTH-1:0]            probe73_out,
      output  [C_PROBE74_WIDTH-1:0]            probe74_out,
      output  [C_PROBE75_WIDTH-1:0]            probe75_out,
      output  [C_PROBE76_WIDTH-1:0]            probe76_out,
      output  [C_PROBE77_WIDTH-1:0]            probe77_out,
      output  [C_PROBE78_WIDTH-1:0]            probe78_out,
      output  [C_PROBE79_WIDTH-1:0]            probe79_out,
      output  [C_PROBE80_WIDTH-1:0]            probe80_out,
      output  [C_PROBE81_WIDTH-1:0]            probe81_out,
      output  [C_PROBE82_WIDTH-1:0]            probe82_out,
      output  [C_PROBE83_WIDTH-1:0]            probe83_out,
      output  [C_PROBE84_WIDTH-1:0]            probe84_out,
      output  [C_PROBE85_WIDTH-1:0]            probe85_out,
      output  [C_PROBE86_WIDTH-1:0]            probe86_out,
      output  [C_PROBE87_WIDTH-1:0]            probe87_out,
      output  [C_PROBE88_WIDTH-1:0]            probe88_out,
      output  [C_PROBE89_WIDTH-1:0]            probe89_out,
      output  [C_PROBE90_WIDTH-1:0]            probe90_out,
      output  [C_PROBE91_WIDTH-1:0]            probe91_out,
      output  [C_PROBE92_WIDTH-1:0]            probe92_out,
      output  [C_PROBE93_WIDTH-1:0]            probe93_out,
      output  [C_PROBE94_WIDTH-1:0]            probe94_out,
      output  [C_PROBE95_WIDTH-1:0]            probe95_out,
      output  [C_PROBE96_WIDTH-1:0]            probe96_out,
      output  [C_PROBE97_WIDTH-1:0]            probe97_out,
      output  [C_PROBE98_WIDTH-1:0]            probe98_out,
      output  [C_PROBE99_WIDTH-1:0]            probe99_out,
      output  [C_PROBE100_WIDTH-1:0]           probe100_out,
      output  [C_PROBE101_WIDTH-1:0]           probe101_out,
      output  [C_PROBE102_WIDTH-1:0]           probe102_out,
      output  [C_PROBE103_WIDTH-1:0]           probe103_out,
      output  [C_PROBE104_WIDTH-1:0]           probe104_out,
      output  [C_PROBE105_WIDTH-1:0]           probe105_out,
      output  [C_PROBE106_WIDTH-1:0]           probe106_out,
      output  [C_PROBE107_WIDTH-1:0]           probe107_out,
      output  [C_PROBE108_WIDTH-1:0]           probe108_out,
      output  [C_PROBE109_WIDTH-1:0]           probe109_out,
      output  [C_PROBE110_WIDTH-1:0]           probe110_out,
      output  [C_PROBE111_WIDTH-1:0]           probe111_out,
      output  [C_PROBE112_WIDTH-1:0]           probe112_out,
      output  [C_PROBE113_WIDTH-1:0]           probe113_out,
      output  [C_PROBE114_WIDTH-1:0]           probe114_out,
      output  [C_PROBE115_WIDTH-1:0]           probe115_out,
      output  [C_PROBE116_WIDTH-1:0]           probe116_out,
      output  [C_PROBE117_WIDTH-1:0]           probe117_out,
      output  [C_PROBE118_WIDTH-1:0]           probe118_out,
      output  [C_PROBE119_WIDTH-1:0]           probe119_out,
      output  [C_PROBE120_WIDTH-1:0]           probe120_out,
      output  [C_PROBE121_WIDTH-1:0]           probe121_out,
      output  [C_PROBE122_WIDTH-1:0]           probe122_out,
      output  [C_PROBE123_WIDTH-1:0]           probe123_out,
      output  [C_PROBE124_WIDTH-1:0]           probe124_out,
      output  [C_PROBE125_WIDTH-1:0]           probe125_out,
      output  [C_PROBE126_WIDTH-1:0]           probe126_out,
      output  [C_PROBE127_WIDTH-1:0]           probe127_out,
      output  [C_PROBE128_WIDTH-1:0]           probe128_out,
      output  [C_PROBE129_WIDTH-1:0]           probe129_out,
      output  [C_PROBE130_WIDTH-1:0]           probe130_out,
      output  [C_PROBE131_WIDTH-1:0]           probe131_out,
      output  [C_PROBE132_WIDTH-1:0]           probe132_out,
      output  [C_PROBE133_WIDTH-1:0]           probe133_out,
      output  [C_PROBE134_WIDTH-1:0]           probe134_out,
      output  [C_PROBE135_WIDTH-1:0]           probe135_out,
      output  [C_PROBE136_WIDTH-1:0]           probe136_out,
      output  [C_PROBE137_WIDTH-1:0]           probe137_out,
      output  [C_PROBE138_WIDTH-1:0]           probe138_out,
      output  [C_PROBE139_WIDTH-1:0]           probe139_out,
      output  [C_PROBE140_WIDTH-1:0]           probe140_out,
      output  [C_PROBE141_WIDTH-1:0]           probe141_out,
      output  [C_PROBE142_WIDTH-1:0]           probe142_out,
      output  [C_PROBE143_WIDTH-1:0]           probe143_out,
      output  [C_PROBE144_WIDTH-1:0]           probe144_out,
      output  [C_PROBE145_WIDTH-1:0]           probe145_out,
      output  [C_PROBE146_WIDTH-1:0]           probe146_out,
      output  [C_PROBE147_WIDTH-1:0]           probe147_out,
      output  [C_PROBE148_WIDTH-1:0]           probe148_out,
      output  [C_PROBE149_WIDTH-1:0]           probe149_out,
      output  [C_PROBE150_WIDTH-1:0]           probe150_out,
      output  [C_PROBE151_WIDTH-1:0]           probe151_out,
      output  [C_PROBE152_WIDTH-1:0]           probe152_out,
      output  [C_PROBE153_WIDTH-1:0]           probe153_out,
      output  [C_PROBE154_WIDTH-1:0]           probe154_out,
      output  [C_PROBE155_WIDTH-1:0]           probe155_out,
      output  [C_PROBE156_WIDTH-1:0]           probe156_out,
      output  [C_PROBE157_WIDTH-1:0]           probe157_out,
      output  [C_PROBE158_WIDTH-1:0]           probe158_out,
      output  [C_PROBE159_WIDTH-1:0]           probe159_out,
      output  [C_PROBE160_WIDTH-1:0]           probe160_out,
      output  [C_PROBE161_WIDTH-1:0]           probe161_out,
      output  [C_PROBE162_WIDTH-1:0]           probe162_out,
      output  [C_PROBE163_WIDTH-1:0]           probe163_out,
      output  [C_PROBE164_WIDTH-1:0]           probe164_out,
      output  [C_PROBE165_WIDTH-1:0]           probe165_out,
      output  [C_PROBE166_WIDTH-1:0]           probe166_out,
      output  [C_PROBE167_WIDTH-1:0]           probe167_out,
      output  [C_PROBE168_WIDTH-1:0]           probe168_out,
      output  [C_PROBE169_WIDTH-1:0]           probe169_out,
      output  [C_PROBE170_WIDTH-1:0]           probe170_out,
      output  [C_PROBE171_WIDTH-1:0]           probe171_out,
      output  [C_PROBE172_WIDTH-1:0]           probe172_out,
      output  [C_PROBE173_WIDTH-1:0]           probe173_out,
      output  [C_PROBE174_WIDTH-1:0]           probe174_out,
      output  [C_PROBE175_WIDTH-1:0]           probe175_out,
      output  [C_PROBE176_WIDTH-1:0]           probe176_out,
      output  [C_PROBE177_WIDTH-1:0]           probe177_out,
      output  [C_PROBE178_WIDTH-1:0]           probe178_out,
      output  [C_PROBE179_WIDTH-1:0]           probe179_out,
      output  [C_PROBE180_WIDTH-1:0]           probe180_out,
      output  [C_PROBE181_WIDTH-1:0]           probe181_out,
      output  [C_PROBE182_WIDTH-1:0]           probe182_out,
      output  [C_PROBE183_WIDTH-1:0]           probe183_out,
      output  [C_PROBE184_WIDTH-1:0]           probe184_out,
      output  [C_PROBE185_WIDTH-1:0]           probe185_out,
      output  [C_PROBE186_WIDTH-1:0]           probe186_out,
      output  [C_PROBE187_WIDTH-1:0]           probe187_out,
      output  [C_PROBE188_WIDTH-1:0]           probe188_out,
      output  [C_PROBE189_WIDTH-1:0]           probe189_out,
      output  [C_PROBE190_WIDTH-1:0]           probe190_out,
      output  [C_PROBE191_WIDTH-1:0]           probe191_out,
      output  [C_PROBE192_WIDTH-1:0]           probe192_out,
      output  [C_PROBE193_WIDTH-1:0]           probe193_out,
      output  [C_PROBE194_WIDTH-1:0]           probe194_out,
      output  [C_PROBE195_WIDTH-1:0]           probe195_out,
      output  [C_PROBE196_WIDTH-1:0]           probe196_out,
      output  [C_PROBE197_WIDTH-1:0]           probe197_out,
      output  [C_PROBE198_WIDTH-1:0]           probe198_out,
      output  [C_PROBE199_WIDTH-1:0]           probe199_out,
      output  [C_PROBE200_WIDTH-1:0]           probe200_out,
      output  [C_PROBE201_WIDTH-1:0]           probe201_out,
      output  [C_PROBE202_WIDTH-1:0]           probe202_out,
      output  [C_PROBE203_WIDTH-1:0]           probe203_out,
      output  [C_PROBE204_WIDTH-1:0]           probe204_out,
      output  [C_PROBE205_WIDTH-1:0]           probe205_out,
      output  [C_PROBE206_WIDTH-1:0]           probe206_out,
      output  [C_PROBE207_WIDTH-1:0]           probe207_out,
      output  [C_PROBE208_WIDTH-1:0]           probe208_out,
      output  [C_PROBE209_WIDTH-1:0]           probe209_out,
      output  [C_PROBE210_WIDTH-1:0]           probe210_out,
      output  [C_PROBE211_WIDTH-1:0]           probe211_out,
      output  [C_PROBE212_WIDTH-1:0]           probe212_out,
      output  [C_PROBE213_WIDTH-1:0]           probe213_out,
      output  [C_PROBE214_WIDTH-1:0]           probe214_out,
      output  [C_PROBE215_WIDTH-1:0]           probe215_out,
      output  [C_PROBE216_WIDTH-1:0]           probe216_out,
      output  [C_PROBE217_WIDTH-1:0]           probe217_out,
      output  [C_PROBE218_WIDTH-1:0]           probe218_out,
      output  [C_PROBE219_WIDTH-1:0]           probe219_out,
      output  [C_PROBE220_WIDTH-1:0]           probe220_out,
      output  [C_PROBE221_WIDTH-1:0]           probe221_out,
      output  [C_PROBE222_WIDTH-1:0]           probe222_out,
      output  [C_PROBE223_WIDTH-1:0]           probe223_out,
      output  [C_PROBE224_WIDTH-1:0]           probe224_out,
      output  [C_PROBE225_WIDTH-1:0]           probe225_out,
      output  [C_PROBE226_WIDTH-1:0]           probe226_out,
      output  [C_PROBE227_WIDTH-1:0]           probe227_out,
      output  [C_PROBE228_WIDTH-1:0]           probe228_out,
      output  [C_PROBE229_WIDTH-1:0]           probe229_out,
      output  [C_PROBE230_WIDTH-1:0]           probe230_out,
      output  [C_PROBE231_WIDTH-1:0]           probe231_out,
      output  [C_PROBE232_WIDTH-1:0]           probe232_out,
      output  [C_PROBE233_WIDTH-1:0]           probe233_out,
      output  [C_PROBE234_WIDTH-1:0]           probe234_out,
      output  [C_PROBE235_WIDTH-1:0]           probe235_out,
      output  [C_PROBE236_WIDTH-1:0]           probe236_out,
      output  [C_PROBE237_WIDTH-1:0]           probe237_out,
      output  [C_PROBE238_WIDTH-1:0]           probe238_out,
      output  [C_PROBE239_WIDTH-1:0]           probe239_out,
      output  [C_PROBE240_WIDTH-1:0]           probe240_out,
      output  [C_PROBE241_WIDTH-1:0]           probe241_out,
      output  [C_PROBE242_WIDTH-1:0]           probe242_out,
      output  [C_PROBE243_WIDTH-1:0]           probe243_out,
      output  [C_PROBE244_WIDTH-1:0]           probe244_out,
      output  [C_PROBE245_WIDTH-1:0]           probe245_out,
      output  [C_PROBE246_WIDTH-1:0]           probe246_out,
      output  [C_PROBE247_WIDTH-1:0]           probe247_out,
      output  [C_PROBE248_WIDTH-1:0]           probe248_out,
      output  [C_PROBE249_WIDTH-1:0]           probe249_out,
      output  [C_PROBE250_WIDTH-1:0]           probe250_out,
      output  [C_PROBE251_WIDTH-1:0]           probe251_out,
      output  [C_PROBE252_WIDTH-1:0]           probe252_out,
      output  [C_PROBE253_WIDTH-1:0]           probe253_out,
      output  [C_PROBE254_WIDTH-1:0]           probe254_out,
      output  [C_PROBE255_WIDTH-1:0]           probe255_out,
      output  [C_PROBE256_WIDTH-1:0]           probe256_out,
      output  [C_PROBE257_WIDTH-1:0]           probe257_out,
      output  [C_PROBE258_WIDTH-1:0]           probe258_out,
      output  [C_PROBE259_WIDTH-1:0]           probe259_out,
      output  [C_PROBE260_WIDTH-1:0]           probe260_out,
      output  [C_PROBE261_WIDTH-1:0]           probe261_out,
      output  [C_PROBE262_WIDTH-1:0]           probe262_out,
      output  [C_PROBE263_WIDTH-1:0]           probe263_out,
      output  [C_PROBE264_WIDTH-1:0]           probe264_out,
      output  [C_PROBE265_WIDTH-1:0]           probe265_out,
      output  [C_PROBE266_WIDTH-1:0]           probe266_out,
      output  [C_PROBE267_WIDTH-1:0]           probe267_out,
      output  [C_PROBE268_WIDTH-1:0]           probe268_out,
      output  [C_PROBE269_WIDTH-1:0]           probe269_out,
      output  [C_PROBE270_WIDTH-1:0]           probe270_out,
      output  [C_PROBE271_WIDTH-1:0]           probe271_out,
      output  [C_PROBE272_WIDTH-1:0]           probe272_out,
      output  [C_PROBE273_WIDTH-1:0]           probe273_out,
      output  [C_PROBE274_WIDTH-1:0]           probe274_out,
      output  [C_PROBE275_WIDTH-1:0]           probe275_out,
      output  [C_PROBE276_WIDTH-1:0]           probe276_out,
      output  [C_PROBE277_WIDTH-1:0]           probe277_out,
      output  [C_PROBE278_WIDTH-1:0]           probe278_out,
      output  [C_PROBE279_WIDTH-1:0]           probe279_out,
      output  [C_PROBE280_WIDTH-1:0]           probe280_out,
      output  [C_PROBE281_WIDTH-1:0]           probe281_out,
      output  [C_PROBE282_WIDTH-1:0]           probe282_out,
      output  [C_PROBE283_WIDTH-1:0]           probe283_out,
      output  [C_PROBE284_WIDTH-1:0]           probe284_out,
      output  [C_PROBE285_WIDTH-1:0]           probe285_out,
      output  [C_PROBE286_WIDTH-1:0]           probe286_out,
      output  [C_PROBE287_WIDTH-1:0]           probe287_out,
      output  [C_PROBE288_WIDTH-1:0]           probe288_out,
      output  [C_PROBE289_WIDTH-1:0]           probe289_out,
      output  [C_PROBE290_WIDTH-1:0]           probe290_out,
      output  [C_PROBE291_WIDTH-1:0]           probe291_out,
      output  [C_PROBE292_WIDTH-1:0]           probe292_out,
      output  [C_PROBE293_WIDTH-1:0]           probe293_out,
      output  [C_PROBE294_WIDTH-1:0]           probe294_out,
      output  [C_PROBE295_WIDTH-1:0]           probe295_out,
      output  [C_PROBE296_WIDTH-1:0]           probe296_out,
      output  [C_PROBE297_WIDTH-1:0]           probe297_out,
      output  [C_PROBE298_WIDTH-1:0]           probe298_out,
      output  [C_PROBE299_WIDTH-1:0]           probe299_out,
      output  [C_PROBE300_WIDTH-1:0]           probe300_out,
      output  [C_PROBE301_WIDTH-1:0]           probe301_out,
      output  [C_PROBE302_WIDTH-1:0]           probe302_out,
      output  [C_PROBE303_WIDTH-1:0]           probe303_out,
      output  [C_PROBE304_WIDTH-1:0]           probe304_out,
      output  [C_PROBE305_WIDTH-1:0]           probe305_out,
      output  [C_PROBE306_WIDTH-1:0]           probe306_out,
      output  [C_PROBE307_WIDTH-1:0]           probe307_out,
      output  [C_PROBE308_WIDTH-1:0]           probe308_out,
      output  [C_PROBE309_WIDTH-1:0]           probe309_out,
      output  [C_PROBE310_WIDTH-1:0]           probe310_out,
      output  [C_PROBE311_WIDTH-1:0]           probe311_out,
      output  [C_PROBE312_WIDTH-1:0]           probe312_out,
      output  [C_PROBE313_WIDTH-1:0]           probe313_out,
      output  [C_PROBE314_WIDTH-1:0]           probe314_out,
      output  [C_PROBE315_WIDTH-1:0]           probe315_out,
      output  [C_PROBE316_WIDTH-1:0]           probe316_out,
      output  [C_PROBE317_WIDTH-1:0]           probe317_out,
      output  [C_PROBE318_WIDTH-1:0]           probe318_out,
      output  [C_PROBE319_WIDTH-1:0]           probe319_out,
      output  [C_PROBE320_WIDTH-1:0]           probe320_out,
      output  [C_PROBE321_WIDTH-1:0]           probe321_out,
      output  [C_PROBE322_WIDTH-1:0]           probe322_out,
      output  [C_PROBE323_WIDTH-1:0]           probe323_out,
      output  [C_PROBE324_WIDTH-1:0]           probe324_out,
      output  [C_PROBE325_WIDTH-1:0]           probe325_out,
      output  [C_PROBE326_WIDTH-1:0]           probe326_out,
      output  [C_PROBE327_WIDTH-1:0]           probe327_out,
      output  [C_PROBE328_WIDTH-1:0]           probe328_out,
      output  [C_PROBE329_WIDTH-1:0]           probe329_out,
      output  [C_PROBE330_WIDTH-1:0]           probe330_out,
      output  [C_PROBE331_WIDTH-1:0]           probe331_out,
      output  [C_PROBE332_WIDTH-1:0]           probe332_out,
      output  [C_PROBE333_WIDTH-1:0]           probe333_out,
      output  [C_PROBE334_WIDTH-1:0]           probe334_out,
      output  [C_PROBE335_WIDTH-1:0]           probe335_out,
      output  [C_PROBE336_WIDTH-1:0]           probe336_out,
      output  [C_PROBE337_WIDTH-1:0]           probe337_out,
      output  [C_PROBE338_WIDTH-1:0]           probe338_out,
      output  [C_PROBE339_WIDTH-1:0]           probe339_out,
      output  [C_PROBE340_WIDTH-1:0]           probe340_out,
      output  [C_PROBE341_WIDTH-1:0]           probe341_out,
      output  [C_PROBE342_WIDTH-1:0]           probe342_out,
      output  [C_PROBE343_WIDTH-1:0]           probe343_out,
      output  [C_PROBE344_WIDTH-1:0]           probe344_out,
      output  [C_PROBE345_WIDTH-1:0]           probe345_out,
      output  [C_PROBE346_WIDTH-1:0]           probe346_out,
      output  [C_PROBE347_WIDTH-1:0]           probe347_out,
      output  [C_PROBE348_WIDTH-1:0]           probe348_out,
      output  [C_PROBE349_WIDTH-1:0]           probe349_out,
      output  [C_PROBE350_WIDTH-1:0]           probe350_out,
      output  [C_PROBE351_WIDTH-1:0]           probe351_out,
      output  [C_PROBE352_WIDTH-1:0]           probe352_out,
      output  [C_PROBE353_WIDTH-1:0]           probe353_out,
      output  [C_PROBE354_WIDTH-1:0]           probe354_out,
      output  [C_PROBE355_WIDTH-1:0]           probe355_out,
      output  [C_PROBE356_WIDTH-1:0]           probe356_out,
      output  [C_PROBE357_WIDTH-1:0]           probe357_out,
      output  [C_PROBE358_WIDTH-1:0]           probe358_out,
      output  [C_PROBE359_WIDTH-1:0]           probe359_out,
      output  [C_PROBE360_WIDTH-1:0]           probe360_out,
      output  [C_PROBE361_WIDTH-1:0]           probe361_out,
      output  [C_PROBE362_WIDTH-1:0]           probe362_out,
      output  [C_PROBE363_WIDTH-1:0]           probe363_out,
      output  [C_PROBE364_WIDTH-1:0]           probe364_out,
      output  [C_PROBE365_WIDTH-1:0]           probe365_out,
      output  [C_PROBE366_WIDTH-1:0]           probe366_out,
      output  [C_PROBE367_WIDTH-1:0]           probe367_out,
      output  [C_PROBE368_WIDTH-1:0]           probe368_out,
      output  [C_PROBE369_WIDTH-1:0]           probe369_out,
      output  [C_PROBE370_WIDTH-1:0]           probe370_out,
      output  [C_PROBE371_WIDTH-1:0]           probe371_out,
      output  [C_PROBE372_WIDTH-1:0]           probe372_out,
      output  [C_PROBE373_WIDTH-1:0]           probe373_out,
      output  [C_PROBE374_WIDTH-1:0]           probe374_out,
      output  [C_PROBE375_WIDTH-1:0]           probe375_out,
      output  [C_PROBE376_WIDTH-1:0]           probe376_out,
      output  [C_PROBE377_WIDTH-1:0]           probe377_out,
      output  [C_PROBE378_WIDTH-1:0]           probe378_out,
      output  [C_PROBE379_WIDTH-1:0]           probe379_out,
      output  [C_PROBE380_WIDTH-1:0]           probe380_out,
      output  [C_PROBE381_WIDTH-1:0]           probe381_out,
      output  [C_PROBE382_WIDTH-1:0]           probe382_out,
      output  [C_PROBE383_WIDTH-1:0]           probe383_out,
      output  [C_PROBE384_WIDTH-1:0]           probe384_out,
      output  [C_PROBE385_WIDTH-1:0]           probe385_out,
      output  [C_PROBE386_WIDTH-1:0]           probe386_out,
      output  [C_PROBE387_WIDTH-1:0]           probe387_out,
      output  [C_PROBE388_WIDTH-1:0]           probe388_out,
      output  [C_PROBE389_WIDTH-1:0]           probe389_out,
      output  [C_PROBE390_WIDTH-1:0]           probe390_out,
      output  [C_PROBE391_WIDTH-1:0]           probe391_out,
      output  [C_PROBE392_WIDTH-1:0]           probe392_out,
      output  [C_PROBE393_WIDTH-1:0]           probe393_out,
      output  [C_PROBE394_WIDTH-1:0]           probe394_out,
      output  [C_PROBE395_WIDTH-1:0]           probe395_out,
      output  [C_PROBE396_WIDTH-1:0]           probe396_out,
      output  [C_PROBE397_WIDTH-1:0]           probe397_out,
      output  [C_PROBE398_WIDTH-1:0]           probe398_out,
      output  [C_PROBE399_WIDTH-1:0]           probe399_out,
      output  [C_PROBE400_WIDTH-1:0]           probe400_out,
      output  [C_PROBE401_WIDTH-1:0]           probe401_out,
      output  [C_PROBE402_WIDTH-1:0]           probe402_out,
      output  [C_PROBE403_WIDTH-1:0]           probe403_out,
      output  [C_PROBE404_WIDTH-1:0]           probe404_out,
      output  [C_PROBE405_WIDTH-1:0]           probe405_out,
      output  [C_PROBE406_WIDTH-1:0]           probe406_out,
      output  [C_PROBE407_WIDTH-1:0]           probe407_out,
      output  [C_PROBE408_WIDTH-1:0]           probe408_out,
      output  [C_PROBE409_WIDTH-1:0]           probe409_out,
      output  [C_PROBE410_WIDTH-1:0]           probe410_out,
      output  [C_PROBE411_WIDTH-1:0]           probe411_out,
      output  [C_PROBE412_WIDTH-1:0]           probe412_out,
      output  [C_PROBE413_WIDTH-1:0]           probe413_out,
      output  [C_PROBE414_WIDTH-1:0]           probe414_out,
      output  [C_PROBE415_WIDTH-1:0]           probe415_out,
      output  [C_PROBE416_WIDTH-1:0]           probe416_out,
      output  [C_PROBE417_WIDTH-1:0]           probe417_out,
      output  [C_PROBE418_WIDTH-1:0]           probe418_out,
      output  [C_PROBE419_WIDTH-1:0]           probe419_out,
      output  [C_PROBE420_WIDTH-1:0]           probe420_out,
      output  [C_PROBE421_WIDTH-1:0]           probe421_out,
      output  [C_PROBE422_WIDTH-1:0]           probe422_out,
      output  [C_PROBE423_WIDTH-1:0]           probe423_out,
      output  [C_PROBE424_WIDTH-1:0]           probe424_out,
      output  [C_PROBE425_WIDTH-1:0]           probe425_out,
      output  [C_PROBE426_WIDTH-1:0]           probe426_out,
      output  [C_PROBE427_WIDTH-1:0]           probe427_out,
      output  [C_PROBE428_WIDTH-1:0]           probe428_out,
      output  [C_PROBE429_WIDTH-1:0]           probe429_out,
      output  [C_PROBE430_WIDTH-1:0]           probe430_out,
      output  [C_PROBE431_WIDTH-1:0]           probe431_out,
      output  [C_PROBE432_WIDTH-1:0]           probe432_out,
      output  [C_PROBE433_WIDTH-1:0]           probe433_out,
      output  [C_PROBE434_WIDTH-1:0]           probe434_out,
      output  [C_PROBE435_WIDTH-1:0]           probe435_out,
      output  [C_PROBE436_WIDTH-1:0]           probe436_out,
      output  [C_PROBE437_WIDTH-1:0]           probe437_out,
      output  [C_PROBE438_WIDTH-1:0]           probe438_out,
      output  [C_PROBE439_WIDTH-1:0]           probe439_out,
      output  [C_PROBE440_WIDTH-1:0]           probe440_out,
      output  [C_PROBE441_WIDTH-1:0]           probe441_out,
      output  [C_PROBE442_WIDTH-1:0]           probe442_out,
      output  [C_PROBE443_WIDTH-1:0]           probe443_out,
      output  [C_PROBE444_WIDTH-1:0]           probe444_out,
      output  [C_PROBE445_WIDTH-1:0]           probe445_out,
      output  [C_PROBE446_WIDTH-1:0]           probe446_out,
      output  [C_PROBE447_WIDTH-1:0]           probe447_out,
      output  [C_PROBE448_WIDTH-1:0]           probe448_out,
      output  [C_PROBE449_WIDTH-1:0]           probe449_out,
      output  [C_PROBE450_WIDTH-1:0]           probe450_out,
      output  [C_PROBE451_WIDTH-1:0]           probe451_out,
      output  [C_PROBE452_WIDTH-1:0]           probe452_out,
      output  [C_PROBE453_WIDTH-1:0]           probe453_out,
      output  [C_PROBE454_WIDTH-1:0]           probe454_out,
      output  [C_PROBE455_WIDTH-1:0]           probe455_out,
      output  [C_PROBE456_WIDTH-1:0]           probe456_out,
      output  [C_PROBE457_WIDTH-1:0]           probe457_out,
      output  [C_PROBE458_WIDTH-1:0]           probe458_out,
      output  [C_PROBE459_WIDTH-1:0]           probe459_out,
      output  [C_PROBE460_WIDTH-1:0]           probe460_out,
      output  [C_PROBE461_WIDTH-1:0]           probe461_out,
      output  [C_PROBE462_WIDTH-1:0]           probe462_out,
      output  [C_PROBE463_WIDTH-1:0]           probe463_out,
      output  [C_PROBE464_WIDTH-1:0]           probe464_out,
      output  [C_PROBE465_WIDTH-1:0]           probe465_out,
      output  [C_PROBE466_WIDTH-1:0]           probe466_out,
      output  [C_PROBE467_WIDTH-1:0]           probe467_out,
      output  [C_PROBE468_WIDTH-1:0]           probe468_out,
      output  [C_PROBE469_WIDTH-1:0]           probe469_out,
      output  [C_PROBE470_WIDTH-1:0]           probe470_out,
      output  [C_PROBE471_WIDTH-1:0]           probe471_out,
      output  [C_PROBE472_WIDTH-1:0]           probe472_out,
      output  [C_PROBE473_WIDTH-1:0]           probe473_out,
      output  [C_PROBE474_WIDTH-1:0]           probe474_out,
      output  [C_PROBE475_WIDTH-1:0]           probe475_out,
      output  [C_PROBE476_WIDTH-1:0]           probe476_out,
      output  [C_PROBE477_WIDTH-1:0]           probe477_out,
      output  [C_PROBE478_WIDTH-1:0]           probe478_out,
      output  [C_PROBE479_WIDTH-1:0]           probe479_out,
      output  [C_PROBE480_WIDTH-1:0]           probe480_out,
      output  [C_PROBE481_WIDTH-1:0]           probe481_out,
      output  [C_PROBE482_WIDTH-1:0]           probe482_out,
      output  [C_PROBE483_WIDTH-1:0]           probe483_out,
      output  [C_PROBE484_WIDTH-1:0]           probe484_out,
      output  [C_PROBE485_WIDTH-1:0]           probe485_out,
      output  [C_PROBE486_WIDTH-1:0]           probe486_out,
      output  [C_PROBE487_WIDTH-1:0]           probe487_out,
      output  [C_PROBE488_WIDTH-1:0]           probe488_out,
      output  [C_PROBE489_WIDTH-1:0]           probe489_out,
      output  [C_PROBE490_WIDTH-1:0]           probe490_out,
      output  [C_PROBE491_WIDTH-1:0]           probe491_out,
      output  [C_PROBE492_WIDTH-1:0]           probe492_out,
      output  [C_PROBE493_WIDTH-1:0]           probe493_out,
      output  [C_PROBE494_WIDTH-1:0]           probe494_out,
      output  [C_PROBE495_WIDTH-1:0]           probe495_out,
      output  [C_PROBE496_WIDTH-1:0]           probe496_out,
      output  [C_PROBE497_WIDTH-1:0]           probe497_out,
      output  [C_PROBE498_WIDTH-1:0]           probe498_out,
      output  [C_PROBE499_WIDTH-1:0]           probe499_out,
      output  [C_PROBE500_WIDTH-1:0]           probe500_out,
      output  [C_PROBE501_WIDTH-1:0]           probe501_out,
      output  [C_PROBE502_WIDTH-1:0]           probe502_out,
      output  [C_PROBE503_WIDTH-1:0]           probe503_out,
      output  [C_PROBE504_WIDTH-1:0]           probe504_out,
      output  [C_PROBE505_WIDTH-1:0]           probe505_out,
      output  [C_PROBE506_WIDTH-1:0]           probe506_out,
      output  [C_PROBE507_WIDTH-1:0]           probe507_out,
      output  [C_PROBE508_WIDTH-1:0]           probe508_out,
      output  [C_PROBE509_WIDTH-1:0]           probe509_out,
      output  [C_PROBE510_WIDTH-1:0]           probe510_out,
      output  [C_PROBE511_WIDTH-1:0]           probe511_out,
