`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7216)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5IQJj49NipZ8M+awYasSTowTJrB6A8rap+B7QTb8RJkWl5DfThoyJO26
ObQv6/qXG9aE6JUc50CoYD9HN/OD8vHbTe7nQp1teAdlUzooi29P05rEd+oaoecfMIHz36B7ZfYS
46Ei1bhdJNfoLMugMgmrnnt4bNWzER2TfJ7DD+wML79blnAV5IPP/+U282PO1btCnOnUhgKHu3nl
GLpLWaqRxLCb6h1cdDgJYqpv3fsJCoXxIPs28c2wFg2Br6Ia9AGgcrywZGCYDvgry+/NfmIZOWLc
vXKVpA5D9jAOlCDZuQiKOdBearVZxTsxqH+knRr40x1WpB7TbciC/X0gRWFTxAYnmU+NhDqQXcTH
CaHVVwznGujbNjKG9+BwIDTGEcyGM1LNC7PtZOG+kujQQY4+oUA59trzQ76MeS9dpk+J6MEN9BOE
IUSXDaDxEwHomYjVt/S0kUYoLNqQelsKk7d26Z58hpLA1Z8C8JzMVH0YHElBQuPoa63TKy20bJIb
2wW5htlQQS+yCzts/upHBVpWMbvMLx7lj2LzhpwWvGgtwNWU2R4QLkMfm+whA4TyTYlO6tRvRiba
95tsqF7iGluKzooaRPP2nKtceVDI08+upV8bKQ3OvMnFczg93tqV7Tf6ubFa5f8sgHKUHe/SDAxY
e2WWsSThh0Klw9pEpD6vhb19TIly5z4gBFS5c9efoMs2j0yWdkOgaNQnquu3uoiQIHNZ2xCR6en2
iwISSkKOL2BAfguchLRq89Hv076XnmOC6TL5Mpg/QNFHlLC+wwE0VDMFBUI5aJH2QFEG0Oe/IZEC
pfh8p3PXNJDKniRNyere1rRgRwB9/AqiGtZqSpb9Me+6Rj9GXTMRPIKCmGv1VIkBHtmTjjvKdlAf
LsImLCcUNq1L5NmMLlUhKOMfDbz7CQIBfGxa0oVzpckniZkhHgiWAJHveLCb/GRO/Fw2FAVnUfjA
w5mJ5xPx8Q2uub0SlfD18oCPGnmgfs04ZwI6HnE+OFP9SBJbE99MChS+FLEAQnETsG+0rc8ObOL4
vmU4NlOQY+Wt9xT8oCc7GMlFmbWWviCV8FTgUu0h+AkNkcLkYmW2YBXE7duI6Nn3QjbY1duXc7+3
z1oAsDED0zXkfUQH94RXCRaAB8ZNMDYVkMSAGtRwfJcr0cuGcy0GUuVJzEv3Y9dW74q4Oal0+2Ih
gsYgIJOizfTQmRrqzy2255clEHPDlAWqv/7Nwe7eB6SvAwrNar5Hs/ChWKlofhwomllWa3zvF429
o3kncKJZ2hOimt+7JqmNjiq6gOlELFwDxljszqT4+7vlUszgqqpHjssSwzcnOf0cY4QPqHeUXDrz
UsCEriE9rhO1bBkZaO1X852taHlAqwtzMJINw+ilszMDl062pv/YU1/ecX58GlNopgKHQLrkwz1p
bCgnPH75gptXB4g/B/9lPKnRShqXZCVG7SMqBTqfJ3tU6kxULBxWPirYNgXwW0VrlDPqqDLJJFh1
/ThaseOQzSdHMBPzBAQhh1Tp6iiU60SAg4jFxq82Ptiv1AEof8aASLMBymXLAHJLEyMXaxotTFcf
WRpQ9mXGa8a10oQVbCGVEAGXIU8qnDBf7OJhlJIBXKbci7IAKrF+JT77x1bSOp2yNnxQbuJ1CgCo
VLkkmHPyGeTY00RZnZ8Nk/QZzDL5vXkU1JyE9/zPHwmm1+EHnZ52tmzehto2PhOMvEcRQ7dsqYXZ
2a9SxEGMPw/T6ZSMIIayb6P1YHPxchKciyj+4qzlSP42Qr4Xf/bEPtF+bHdbp25gx0NXGNtZ9kkf
GnZutapwAjlQu19EmYOSHS6OXAHBW5KLuHlCUw6cXBD/Amx4h17dWtvOnuVhsCTK1ipaU+r8nmcr
ToC31kJ+R8ELXNh+FeSuxsQxHYG99HlgcUhxfVTi4XFj557rWhWObFS2BusEDXvs8XypHGMmBeAm
C4j+vbkpsnzMQPf7Gxd/bcBKURUNBQytCW/ABZh2kJBjQwa4WIOBVnwfgd7O4Up6op3XnPrl+aRQ
26kzDHIIJbKDn5+B3V0FlRJYCiy6wNtD1J/uTHy5tuVRNQR4yId4qFYpsIiWSVCdEgbQ8gw52qZM
sLzCpkrwgZ7+ZmcdPmprqiy7Ba4haeRPTKpoL57V8ny5FPIW2wo8coycu4Nr8rI6a57ECC7ifMou
U8IN/g5u9d3pHbwhetKCKjs/3CsqWw4LCzTJXOK5HQky4m3SMQGrYugPjNzU0/q16m7MOyCseMj1
Uykj0o5xA2PE6fq3XVZob0uZwCh5JwkYCp/r44CUxFXWiD/M3iZFu6VDFdTUsUURRlnk615cEX8l
PXU5eOJksgtqbmLD+Gnh0kcCWdGux11SNJ5aK/C1ersKMia40p9oG6LbcPLExcIbhCqm2jrCEE70
R+vMTWGdANWMzyNgkfhVx48StWtaJFIvNC3sJ17BUxngtaK2kweU+R0sNDA4ORu/6XJDcX/F++t/
LfnygN8flVMNF/LrZv2TDaInaZzy8PzBqKOrhVbso36PH8/7DzUHN9ULpb/K9rjtZArwXb0ro3oo
XI2Q7XKpZ1+8/kymlD6qfwm/7EbckufRUfklj61G+1TpR6qdUAy4HFDMg9khLplk82isEipRM4TH
btkThJjYnotNNMKpdwIEwHA6716/jzzMgjbiGsZXbjerw18sA0bp7mYrNZqk9CMkm7V1USB7mbgf
vdpG3Qb1mihJYYIlgVDpvHImfegoS116vKLnUGP38XNtxRoYd6nbBgWwcH0kSv+4TMFdx3OJK+Tu
k7w22FTE5IOoMZAzFNF4bR77QptznNPkKDAJrRIwDwLSf3KxXd9dpY4lvvPqQxuUV96Vj4BXNOSn
V9OHlgrAD6FV1QbdG72+DZo0D0x0n6ntjfnK0l5LeUWjdRPscgB8VXYuQvE+b3b32JR7t9x8WpUO
EtsYr1igmCH6tiJ8UyKVHIM6ZPrSKnM+X8zVnb/dEwSdXCD4TpFgM5nNlpzinnJ6UwUkGpdi+2vg
j0QRW8+0eVdU5H/gGBOByiDbja1r/vMJ7nZdh1IVvNFoMfoum934KORkmU/EACzegi38CErdepnt
CC9QEWsErMO5YT6bmmTvdqud4k8MH9mvBU1/vRn/me1AGVdCDXIG3yCi+/FE6U1L6QoI+7ajMd76
PNai0Qp0MArf73DCDJ+KDd1VQH7RbrD5P0GOMeNChRiwtlSDZHgKdYIW3MbR5zZT3DWmYVhUzIIL
oRAGKBWwG60hEBsjYDp0J/laL8ztcvqA7z5Wxc0hDB361cIm0N8GAujFWWEs+TU+QlBDZ/N/KS+O
hnN7ETH0k/mjSikRLPXYtSVZc0fGbGOfMWIbvkzLKZyEuLn2YOIk7NcKFomokUu/YX7vA9a4Atu4
JlTRBglweZpJU7yPpv0dvVATIHO6vIUOxGIpHPzbzHlCu5fIYQ8STN/YsHkxPF+CMEz60BkBwZlX
+ONZcYm61YHRD6D3xVU+HHbhL+V3Tu3FKB+M/VngWKakjOIUtUEgwz2E3pZHlTuO51imb6XRZ1aj
g//B1gE01BGJlDccS7pawajP2XnI59noyYLZKMkpejdDqkyDW6u94Ql4ArKnCZEaMTiI3bCyQi9t
iGx/YdTpNH5rXlkIbikMwQdME0lU2yzsS9wNBFioG1u6WudpHyx5PNWBF2u0fSE89LfENpbLXhzX
uwHd4Hy6pHZjQhsxIdreUcaQZQjDrj20VThlath54u/+L1gZ2/QpJSYavSoSlw+eRWa+58BBUBQt
VEGIpDa/H1X+1TGAuunzxTSUzBKYwx3T4dXL95YH2uh1r+IDBt4jRPMvCoLwoXTKlxMCE8qVXqM2
pqnoOeWys/EnXcghyO5iYQKvxuHzXB04pXhu74lVcTAD+ktdJKvV8jIj5W6jvuHrc9Xy7l0X9d51
TweAv0LfHb8cKg2k8U/xh1/eHpddTG+2G36VCJBhBYpQqutDAYW6+39O/uQzIW3PfeHSfcfjJmG1
0oTgCPArP9xx8YMfxu77ZA5MfSEF8rquiE6vqD1Kg7//09O3XNnoj2pXAhlMCKHRY9e/pwbgVWhK
spz2fqjJqYZ32S+aN9HJ7Bur4Z8JO+a29eqMLW/UsldWkX61QmzI9JQ1DSGCINEsYeg3sEyR0XNT
JwxVaZ6WVD1toJ0A9Q9ITlbjqKxd8/LTytLWcM7KqZPevZv6WDYd+WH/ICbJKrX64lmYcEjGbGx8
Zv6hSUvuQNBbO6JTvTNEG2xWJMSdCMBumMhGiI2nBwKzU2lXwWv7ZPuxiqcQ/CEhLWt8M7iapSpT
nLkWjWBTicjGeTWvcCCf8PS9ZAj+KvKxObofuo+zxK3zliEFabcYpPg+aIpnRmABPtcmAxXPUHYq
W8lD/IAv4OXyZT5lp4B+GWYXg2dE9bLOJshZkPgIr0i3sIOegE8QqMS6QxwUgq8mdi7IZljPl39N
P17Wjp7jc2q8hpW1NWkFzM7VHsJLv0Nb+cZ2lGhrLRS0oNxOlU/kW2aaGlxZRFd8o4/kc1R54Cnm
sJ8yNph4xx0fdyyVXWzAQF746PQxT/8ET+McQ04NRDafvwnM5wBVOYHcsZK9RJDN9OGpevv55yW7
2tvpDzk5sax/m0FKHsBsXGWWJxugSzNZNi4YocVSQTm9K7u9nbW25Mla/jmM/2oRnwLbBXUhAuFy
pUQiahVTnhDxOLbFdU+zlZSe9ZD/0dOiAmJCAX2Jd5/WXjwcca+xEDyTCfG7nQGcV2MKqMoS6EFl
mO+KlHhHLByuDrNRjtWnUGPXzkREOMemKsR+DqaI0AjXOT8DkxBwnOuWLEM2GFcq1Jj+lA+LidnU
f+0kArucWsuUIoRFaB6hH8LbN3YTRRRxbElKubHCJ3NbgIE3LUHI9pXELEO2yTAmoHAVt6Ldw6XS
i3SNHYHC/2c0gRageQL7F3Hm6wpdUtxsgrOmB86W6q2EnMQfZZsPTRbZvkXaKmGjbaJBq86TCpLg
y4IjiLSp7pvzdLtEjPpUSgyO3DEQ9I8Jmk/4cgdSIogvhnVmbWbav46kCVZKnDguzcmnJMUsH7KW
kFXmNv+lZS+CCFeH72u+XM/S12PqNNJ99hWu7GB58GAr7edpiI1jiJ5JH8pQBrMZTXJXYQ7gaqho
roZ4bvW2VPDnWfsGtkcHT9tMRD4+8UMszl6JT+4YsuIz4Xe6X4x95Yc1fczMgUXGV0CqkoNEYyBW
vhw3N8jU54p/YL9QMJuWHlhEgKzoXsV14VDy7bFNmfcxFjoQIhqystUdy0Gar7WqQ0GyLsFdCF3/
RGMNz6pRQQwyAk1M/oo/mOVQ0fPMy3FyIEANx/E0tkPb1uP8sY2xUVRokuS4YUORoZm1gRR1XDwk
ZcbLY5rnOLcxXnP1t5ENRqg5NwZQj9qdOGZMQd6R4HkcRbRTA08MksI7FqWd4FI2frhR71rkmkPt
caXGT/+FB2FghpCX57ylbaWDbetgjLr5VT8gqqZPlBWn/rzfDyqxl7N2Qa8h1+9MlOQ26PGfrepa
EKPraW9ZTA4PKyUdizkNYXYH6WDg6gdTQUkx/Gmblw3kPN/iR0bX1uO3AEaaezHK0HJ26mYJ3dn0
B3iQvB5AcwB/++8UEEMyB6AYkA0QIqhf2qQZv+Dx29DWIDZY1l1P1DQbEAKI1Poyh5CWgMgEihr1
Khk3CamIJK24dMUp6tFPncWf1CeH+C3jnxIpqym1sX4fyaKIpyZAaioXMTLHFBDC1ePMnixv27e4
xk4SpV4medTqWPYYoMVim3CymgAM1I7YkhmBz36i0K0bCkhJ+GgVlhk+FJl1qtqOkQunxGRiGMlA
UgfOYnXnIm48VZXyLmUbAVKDM+91Q3ZY3uJCq6lFTwxVZ94/NHPVvEA+izHKzxdHrxh/CoeNW25i
/gO67ylaKygg0x4CLJcp2XvT+tE9YMocw68RtCjNF3duMi6tR5s6Vf07IFxV1vLfQpeADTIg3p6n
vtvqvAQpjmqc+fDH43xDyLMV2Eyuxb7Efw4Zh0rNKSm4h++Cy/w2bE8LCnPBuv8N3EqEVsR9hANp
A1q0myqnPKSHs5ERDtWjcp5CxbLjsr+EGB6/euVAJ9/lTVMfOAnZO0iLW6aR4VRWblRiKIj/5QRL
4Y//U5ein0Sadk/H/3FgdHSClWFVVKknH/c5Y0m8QhrVrYCvsgSWN+Lc+Tg4E67BCa3vG3nvZXaV
mLJl95YbfN9A//6MWRMQ5M+Tq4Kl9+YxmmoQHZxaPsWgsp4LM8KYDyHpLZ3BYysnBytgHq0QUABT
aDsRFPBlVuIGmxG/c5TdW32WL5umTt2c1OSbDPuA2xNVFj5vMFl3tKyFBRqmXYVylIVQfzsrCGL2
UP/XzL+harHHYZYUm+hh+WVnFZDrQ/BBSjaPYAqCOxgOG2+xadz59tEBTcVAUobhkT2CyexgFdqm
iKsChX3pGBtLS1fTAvhux7dV0WuGViBiwP9KtV+wKhTb3EbFwZCQH1I6x3dN8rDpr+SakPg1aSMt
4PbpkwWIy1sXeRLjR3P9QOmyWLo1yi4oBrBHcmxHNzJcxG0ZUfUNYySsLQgUVvQK0+e7caLmlYs4
qZclZUS/SfKWsYKtD1jOIMHnhQGIQT0g59ZuVOasf/ItCLqSGHUqU2X8+Pc+roa1OkZX+mtb3GqK
y2mKxpE6IVw5gb3g7rlMahpazmMDr7uesZL6Is7zeYPPdlpcE+/o03bf3ibR6pNuOLGAjL5TrUpW
xGJIcgnK5M0K/iwtN4TlsEBIBOgE/RdYw8NaccMwBt0vmii4bZroTmy4b4IBsOM81WpOGtxMtsB9
P1UknAilAjLddauUr1i5VPF8zn669ByhXRrD0xVcutJue4Ihsu7oovqjIWBzXGjSvo5cl1h4DnBT
vGAeTZIyRTu7MKi/z+f96Qp5Fk8tAAcoKtMIyV4Ide8UFf5/jGRQptPaMM2pXwNUpT4NmRUo4U++
+S30rRJWpbsZTXccmn9TIkW4hSts1Kgs2R3nYBmTp+ElOGOAQD3N9jHierTS13SAWTHAnL0XXgn0
CzuVrC30TQk24SZafBFZyEfGmAbIH4P8e1NB6aBNXQm+w+P4QVtqnnTJ+rwAZG7vyoU0Aa8sPEEa
TUV06STJQujehWaRsZKL1m2XPnerHGSmoIfa9l/iDDOlnZv+MXo+6MRpWJsJLcLU1M4GX5gArNXg
W3y64qlsvJ+C9jUcjUby3kgnVf6mnt6tLbkcAwow2HthST8kIHYALva7e571VCXvvRs7gIr25vcP
CQdZBfo1k8vutR3U7CtGUYfhuX9/O2+cHs7g4VjoLRjw4o/SZNiy+VkSoK8SO+ZKlhjHJ1R1+QKW
EbSrAIyG84eEy1B8nFfPvDLXyKnL9/RCUKOEY0QTluvd/2tZ29QN8rZJZ4xoSvronNUngJVAVB7s
PV7HQCs9VG5PCJnz1V5CDskC4752Ko5aWqqg4Qofdmas2uvQaqfP/zLzQtE05wQmqMg7ZH9qpkgc
wSQ5Df/wDid51Sq1HATYor8I7W9K5iUAFWaTYeLlPnNfcNKVsuszr8ycIEaQGisTA5tT+WFFJtQe
eeHe4nCVn1hd+1HT3bhtAjgrZOMMPQyNS8mWu59+uwX8g+Q5GjvvspmAv4/VoC2MwSouVgv15SjK
tmIMHMTrB/idnhBLPwoZAtr3CGErwIrCRjcXVbEHNwbgCgl48BfBpVApXM3srhgAUjb5W1B5YT4T
6khIdvcPy0skrOilmKUzTPG14z+acMwKwZ7+az1M3HkPO44KFm1A15HCQJ+oxWjYhiVjE3ZUqXZ2
pM0wsWQxRTit6AYpn1Ko8gzz1w2mEUxuE4jz1w6cbd1tAqXu/HLXennOqoJfYqXPWnhhXtZch2TA
U2R8e97GOcG5EDwsqpqeo0ZKXbwvyzw0d7y1WXi+EmyMBnNo6KG/xSVDqMhNCVj00jlz7xQRWjNW
1aqTUa7tkGUqvB2U+iPp7QvHK5r4JvIUfZ1PJYi9m+Tggz2IQq7RA1AZxFtpLWEHphkKHTyJ5tNs
u+8JxKH4fR8BzpwoGXoxomYBtxmWPbzaB2zkU7gKvqvCJfAEWxcwam9dBxw/ywvrA48j8GpmLWoV
AnWf7iSp+kZHwfHsA777qp/t0LtTd05zqIjcTJsOT4sfAM4996wMNz+iL9KZm0R9qAiJLVNoxEBk
qLfLUQ5zJSNvfoml1DDacdkMLdKRKEShBzhiv5CnV/4+acWtLq7AS77zPGHv6cU40kvwWGsSwY66
XodonlowO7NAp3vFdyQvF8a/jJNwQ54WIMvam3KC6xOi0VeVF7c741zAmJtDu/WxoAjcy5g9PDeX
ylxriAeMlu+Ww3n8XaDpomWz1jn1KK+K2Y9JdRSvs2g47cO8E40LNUHBmz1B4FnB6zRhForT6I7g
t92TQewmawfuVVHU+94foxt31mTAp53Hu6SEm2SDZ4pEUIA+8bwrIEzhSdyMM77IhxLrcJJypm+k
PCBzME5nu0cxHeiCiCeP8CSCvzOtaEl7N6q8SJx7/ZrpJcnhzPfGWa7XwQWeHNNo9Uu8GWBppdRB
LluX48XqFNHVvqhN/7AMjLT2XQz474183b2Ki99VRh53paAzdi5kxna665aBVdy0I5uENLa6LG6W
rrfKtrBLcr2uqxFuUixuwcW/Em8xgCpxVQhfIqPBXk9QNlxvepQJmGqo5do4K/RIRoWN2Og3j9t0
GMTym0kOH+9dmbplQ+38BkgpyGc1VdyVovvx3HT5eTiedtpNcM8/JHBr8Gt2rHxaevKVlbvQZd9f
dnSDgxjfyzTP6YtYeL3WQ0dWLOgQT0GY81v26tsF7YxnLKrb9mBczfHtFULH6s/ewhqr0IZ4aQnr
eYiml5PgITlf1/vcSncK8F31bw0D/GITEDjIv1SbOyuJkHCgxqPv5piYSA4+pFxbsJW5iod3iMhw
nx7aKBpqHR6weNRR5C2nmgeJNYxa9SucNF4klCVjMhn74Nd7X2o3hb4ce5LwWKX1agtk4ylw7Ltg
7LSuJep21ROQUXiBmz6jnKcMrVY+QwseR4qZmFM+20NrEHb585P4Kf6qNds2dLxo7w8ioLEdAJfs
kacGYmlvdNmGwtIiLjF6P3yLcQOGPrPPhkVNjov2AnzNR+TmYOgQn6KqhFoEdWDKVSEDe8DZBnZe
TzhldqAtdObpEfNnv3o1cZK9Cfkl3apTTJKzdcgoMBDrBZPOTnaDDyTJ8hUSdFDqoUxJ5ztkWZ5M
EX88TOTmPtGuV16uyVqKMRK0fGCDC7B6WkEl0WHbbKVO6ahtRDnTOVntODGwfVLVV2pGkQ8sWY+S
vdhPH2Jr3ZGX4+nGpnfAPStqbiUwhZbhGhV2zh6GS0gVQ8Z5SUTBW9Bm7OV71tyQyAeteVlS8cSE
NIfjrR4G99KGv+P/yvd+vba0BMi03oXXFAur0uoylM4F+rGWrmjY9demGD89zBhOoc1axqgs8epD
WL3NIXsgcpnxwT2VpASjUXcvHEe/d6VwKvHdsVsA3RmjXh3M+oA613BLuIvw5vTJp9HpYVN5BRK2
Z/FyqXyhaK3mRKDZa45e+NU+ufcYu80LTg/1ZnGhBG+scA==
`pragma protect end_protected
