`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14960)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5IQJj49NipZ8M+awYasSTowuZocoHyREJavBHjlmjUV15riyMACdDBM4
9FnBKwYblJXXfItaP1UYfC790iu9J97/877G8BJPLKtKAvL62tFnSf2QpVPUMDvD9LBqnf+Us6Rb
MJ3ix789DQkR+m/O2pBQw15fLV0LRUO+Jt9cYnH9Zpu/HDXirQfGDrAjBGVc3wCnhhcVwR7DQ69F
ZvcZySsaciDljO7aYmKH+TEDPF8MITP8nsOlhwo1TIKrQeeKxS6ZuTw6ShlBsCeMovJM7NKlV1K/
iIxKaiSFUnOPpI2Pan7u4wHcB0sw7EprrFcHpRTNjh/L6YtWzAZlvt0D9/m+QFK4cQuTuLLYIMNn
ZUIx2DsuuBtJ9P07P6uCrMtw1mN/6Ff+9vGWItrFMxzRPGxyZgvq58Jv2ARG5j2FIcJ8Q6BVS9gy
X3YhvtJplPFiDv7Lm7QRQExc06jsh1OxxTv6jLHI8b94LIAfGzrvC+EbxFj22LDdiclr4kqx1a59
Yc+JrDPVRe0nkceBdY50Q8JijjFm/WvC2EMc67ud0XR/RcADk+hV4uAG9lOKlPoYniCTUVxnNitB
HLSXqMyHl1CWpa61ENNr4T2h0zQ2wijBZrW9uIvsxrT0R/ngfWgz1qrQ71RImO1/HKNwZItdLB3x
GfZJ3t4k4TDGTsOH//c09m5W7GI4Vu8sd3un39LQgX0A3xqgkrvlTprdL9BcPa5UMnEZ3yIz3VNE
iUFW7+SwvPxfAPG9yMPHuh8jdkSUU29BJzHQfJ37WUP/epWQ9VKLiwsvFEqEIDVisG3swCghNKwE
yrrk7jMcqo/OqIe5OJ5Bv31PRBBjoy2JuHyg8jIaAI4+oQprLoYb/XudrG80OS9OModSZ7EzAhYs
4NjZbwsxIUJNKPJ9QoYFG+Uq30s9dNIUofSnZPT30TwuhuAORID+1iT7tI1bZ7GQCof2K6d2hk2w
w/xu3NRbftT/f0MTV2uJjqH7ItIz0IJWro7UJGe42skYPeg4qDRZ49hDtTde9qYkWQrw2pX2qLRG
NIDEhkQcDImbJarbUzaAUxDrUPyEvdKtEgvX0RbnNJ8HqKpsbkppaUEg9SB30xYHQXVCzcikBdDN
/bFsk60f97yxsZeixtagFwtV2K2kza+RETLT7Jd+k05nLaC3lfy5WyccoO+KEVC+IVUanmjpEFPs
cLGRW6UP6fV8et+WSmoR0Cn4w1uUYt+3akcbd4jqN3L4qLm7yhwlR2rv9ez7L5uHB3fi21tYD6aj
iQdtTXLED9VvkbV3L3XuoqNQejCbtdxK1H5KlL8MYB9LVHphKJp48ffN/bnzexOrVBPpnZ0FZU8g
8El0ETH9yzlcg6rdMdObWKtaf15tJfBWUXqH2mF6HKQ6h0S1Yd5Mn5cy7IJWU/+OFqouv8m3l5BG
Jonl+uVrFhD/QoRhSRmK0wDG13KwHgb5YXBVXO2f1vnBmr4nW4BqbgCg/uvQBEbjgdK0JvQj47xK
26PzKccimffDgX/aUk8o29Kte3o8a9cOLUrUMktou5EzoUb1CiAxc+ZOGM385AuJnMVMZWmq1+py
OBUgCoFht1UcV3vQTK7OvhMFYS1/t+AWN6y9+Urbq/nVbslD3fdRzAQ/eFp8+paCwiQypeGu3Tx+
hAgUN4dYUg1RSptUElxDSzZABrVprZBQCoUMSwVdLJMQX9Uq4JdMAtwlDLgVWiXCuu5jwJ4Yr0tJ
YkfuU+ILnfVSc6N/hmEJY0ilcHRW8aUmVnUkS0i9BF1wxqhw5SPoTubGWrifG/CQYzvMyXJOIMNv
uIzPUjKbfjj4JOqARqHMKlv2ZswuoSL6kHoRLseJZx/IJZMoypTTJvx8dow5r1rIksxFDDKmZdSg
g2zCvrxj/5DxUZAUYPnU1eJn7QhMPpPNa2LGHwJxMuDQYthZJfHBqWjENKhwzE49rznvUc4sgRJf
CBdVYJjdb4ZRbuNiQ8E5xZIYWiqH4WLREYQQzVXfLeWgXB4rf/2plY0TREjtxlETrg/TIGNd7va5
tvKAcCyr6vpBg9TSKQYwDfpuS/eHabgnOr4eg4H6wm5SqFOZhZpeDxVf634/jPhYX8LTAPtqGZOl
uOb7DYRLgIpTBLVTNR/sy2UQvdXWkhW9a4rxXCOHG+ZqP/O5bXz/iUiqSoRrcxsCehixL0yvU3xk
HG2TqW87nTgRagzkmdr38oEzqivssNrGUgQIyJDcwBtS51OiEADn4P/runLOfaFPE/smHBw+GO54
xLntacVL8eNG8VBo5vMtwOAheJu02W6IqqBQHihGFYiF9OFVCM4NcKMzbtTOsc+owdFy/lFLbuQ4
q/tcJCIWhAneWgxIQSVpSUS2oLLJpTs2OG5zoFflpUcdBTgdoBKb/PtwNEOK7pqXOrcfZdj4bcRz
tObge0e8KRMQRCG8xQfwkpfJRDNyLkT9FCZTweHkxGflGuu4oCfvZ5dITqlrNAP/h8cNcH43GwFJ
QveRMadYrLtaFX2c0SdcjbKWwEB7UD7aLFvNEvfglBSIU1ZD/+I4tZAC++hqYX2fE79+SNFOEX7D
Zme2jMreoWrLdd7hcUqJwzvMrxzpA+ahg1yy9Fu6J8BGDNnLxi489SO9Lqk0bxF/GOcunQ++KNg3
2ORcquTil33ODM1Rjy7m1ZhC0ZxdewwIxihDEfPQmgHsOG4x+rQbortmsUT+jYc3IEfw4ah/APRy
8g8bxjhmRsBgIxCW1Mu8u6r/KwItj2/HrLE/S3rqADfdWMoYxcBnfb/Rhh7HuxqgDCeeA8DlkBwS
EQza4AFanjiJAzreVmvPcABE2tjMxoqy2JaCGhE2dXyOV4idpTweSelzjJotNM9jF9EDueloeldP
66JKhPsU5eRk4UDYzEFZ0+YSw+z9pGNEgzs9yEdGq6QphA29IVH6jLvP7vXH4cS7W+PEmqP3eZzL
qFKNDugEAEFJu5H6u+ZS1OKQOf6RFBFBrMpVmlBX2SKQxNIsRUsLRfn91IprdOKRZWyYR3KvZ6in
fQPXBXod1/TqRu5kSoZs2L6s6zrxT2IEN+GzIkLZ98Cdj1AQLgfUWTvKm/QFxwU7TwQhK1OPMElv
EqV1TiJA21CFPe+DEwokAojMhbSnCQRjXnw9ZxfWQfm0ouMwyhQ6aH2AzzG79riRwyKwXWwcyxBQ
Ddl8taU/vZSzW0dtlLCqcuTSjTuFiPcRVJ0TyF15j3TPWWO6WKFERyf++fco4YUC9JGCCwkUm4NY
1C/Uq7NdLnvXmQASo7a6bOcwTrQIyUYZM9LwDEea30/M6ElZ2kU10Mxw0PNzVRImfM1idLrKeNgT
pZ1iGZAtE7DAw+fvXDphoaGla8BN9oxX0D8nK1Ka4y29xGr9opXUdCA7SXP8baJK6Nfqf2DlOyr+
ROv/YtRpHO16jD1j3NtxHSOZW7/DNJ95oRyfkcJiKU0eIkE6kRNfSKRffyIybPpXexTL8VTMYUJ1
21j1X1T1uVAXYMTnmNAUGXLOfQzDBnWEr9TmXpxzEmUTPSSOP7BCT3hSAWlyL6Pc78Gf13pkDkSo
m3pIfSAekvBnhafJc/8sSlEDnQPUmMI9/l8xBeW7Gab0JBVRAcJNrILPfO7rInczStHCkwHGZ4LP
h4O7an5K0BdGha83Wgt8q1pDYyCzGpcz6tUMXPzvSgsiya5tUv9BMNb38m4/bYSyaQyAru2HVLgN
HCEHmPGgM0Euew7HVWhQF8kHdUzXPUpW84YYDaQB+RDchyh65jPzMHsS39W6FcywHm8fAiRM7HX7
7i5ZyXdsh+ZvfkgQ78HafE7AR7/VqyD9qz3wvYbvZKYdbXD9oqoj0XLxi5I647LnsZv3vybNu40W
z3Im+xZCI1jv6GXQT85mmqGuexAzUmroApIYpB4KIQqwzE94iJH3RNRgvlV0tUG3t9eahFmb5gd9
L36vBk6ptA6YvP/dprBcdAKQkZZhZJ7OJM5OGJrbi7d8+CTKXfzvT6VcTD1mAjSCx1xAnKNa+MSN
rMvAVEtKgaIRUXcxbWSntlJT0gl+3SJsJfe8uTefWXsDYM3L/cwA9CJX7Esj+ay1f6bCbJ1c6DmA
jwqiBImNNdKL94jNsjDmbmamEE7F0Qkq8t7Gc2b7e/A0hwSuEcZA68UrNDfko401Bje0Y013oYLi
ibpjMVlvY8xkujBbgn0VsuzsG5t3ZUzqi96XKF2tXxfcISxneRA7wdmlzoYOyQ0oxiA4KrMThdGJ
jmvGPEptWSt/sreXaz6mpVrfaR8F22ZtzwLHZSWGs6wHwGkYV04V067YzCg77wqFpp3POGKomThn
cD7lxNSRQziv1XjwjOk2haJFOu6Zmy+BtnG7ILT113lW2ARtlwxrbMnQArkB6fSAQ6Ob5UPe80mj
K2wH6sOPHMJIPGwOvQpsOLoSbfeMxkqdehy76GjlJs+iiHX3WgBEnm9oBTz7pVREGQF5UosdhdRr
n9MJYZ6U1eckmgrF9/z+VVt1QiW/gbIVXXtMaUlA902UTxEHJHk53BJuYklDUmBNOLNAEktrLaer
8fHsOPymtZfJhkhs8Q4WtsqCI1EVYMHPisu0oZiStxO7OeLnGJX5iVp9bQrZcFdGkay5JHI2Lwop
+AbjXl43OlBQBEs0AkHm+3Rw0Xxwj2GnsB2e9nSKVnp5SLfcxYJX3Ru1PlU10RZNwx0U2DiBuR8z
iq8nDnPLbdqKyzoVQnRJOEX46YyrFoKB0X7+s+0MouIS9NlqOLn4HIGhPodSQLXBrl8zD3JHliV+
hsjbXDapE7eMmizrVOSQUSac1GL8S4KMC4sxzsYXDDZHnJINWuWZGqqyT3ymbOTBdEOpd6kkgNEU
eMkmlfWg8cMw8WHNoIcB/PqeCdAxSZXBNbHNSz6HlH22KkDcRSh7k5gQyrSy3LQmJVxM1BYywhpH
nfgxOvUL8wC0D8mbwFQvyZBT/QXuUCmE1PfigdoM0vfZTlmpRQngN2l9/VE3MijCgqW3AOIAUrN7
4VIuK7GxDApQfEUgUW+S+oeE6iTAXg+BWn8C0o9covJ3ihZPviYk5MLZz3sBcsQ355D9AM+3QbDL
JT3I9dJIXNJXEsC9tKxEl4L9FkL0Xb2PC5KfM/3tx6l6mKhsTCkirtGJnGlerIXaw62OcfVFQoEJ
MDas8nP3Yd2F8vyMTbEs7Tsyq+Md0YkIyRero0LqL0fQggcTNL169gdrOGjos8BcTvyCaOXNuZM+
ixGHDw2sa8HoARdFJD18ECp1tMqaHmbPCZ+W2sOcL4X2lpvuHbDSKUSf6aKxou0vFdxy20ECEF89
xVIFPq24Xo5NwrmQxVBTmZqJXqxn3FGhKS3Bd2gx+zTdH62rKpqjI/WfudhvbMteiCDMoDtS+q2p
1238CmXwaxfLxYcGcQ4RFbX0Do3JsgLq7cANGx0c+qpngkocrIfTAOvfIBhbPSB4+DddPM0ObbiZ
zARDO48uOF+AIbGqC+n5QjZLKSiq+QNWTXFK7HYsY4PT/vnd/tIkI7CP4AinwhHJL6NOAGimBU3/
DYKXSJxlxu69Rxatvet84TM9uDlCWlcf5uxlLVadhQTukBUh7EpNC02ipMHnrwdjsnhwk36E01tx
nDr6AdJ89RopR5ZLrdkoICSuXDdg9RsoYN2EsehorPpjvEJ3stj2QtjBE7Y9cU0G+1G9kWuM5U6b
bMbnWXrD9IzX4pdXbhAvB3ydSwfOjcbHHfy3rFgyDuXd8OhacF0aXXtONpeN895LpC9udNhDQE50
UDq8bkc6wpw2pKvNipo7mxZ5psC4NrIDHoTQ0BUZbQNiRCyUkqYwStaSJ81RluQMOSWtuHaNqka3
cLMAKu9SHE34jFjbBp3ZA9WEc1MSD9luQCCLEJugkIAX2rfFNINt2Wv0kgaDU7oaXgc9XxYSzL2y
2vHzc0Ley9lxSwzOayNJMelmVImkqcxg/dEehL0uoDCwYbKrHDL/V0H4PqN7iMJhYlNbqblO0sv7
31su5LXU0zWmmw6S9+/atZVbbL55CJwNNOsXkNRxSl/FDIsCm9i/XZskKp/r0MIluYQO5MZr7G/Z
8BtSuy34MNndqp1sLhqs5/Sv7yQjJrG2r+NAjrsBJaaraDHicZYGictifj65XC3+E6Z3sTc8vtnF
o6N1Bb7z4tz8e50vrpklQJyJBrXUrGLKyoLJoQ/tfjp/RkjlBOlc7+hsAR8qn5bjT0FKGgKaQBzV
0MARUHUc7RIGiOAmuLoTyBH6nACIua9g/swlBCqQ7QSgCpo0qnQB7/pjXIvkxLzJ4okBPtHdBf0d
4jZQj2pg7rnKwb+jH2rhET/Q2sWqeP83oe2IZMVtD7dbtSM5a2PbStkNDrrBi9fZqGF9aJadrQi9
fpxx8YvjBVBGv1rL8j1I8Y8/8I0HpeCHq9B3vADlAoIJ22xpkBLY2SiQ/N+wFjqzd4bnXZRBD7aL
dDrBb71seAnEMn6UBpX8IEn3duwomHsTJ2JnbZbUc+TbPkVCoAO7nxbA1IkhpX+egWbKxE/Tajgv
EsawgWxO467n6ILQOndzLdlWI1B17sEYI4SDQk03ys6TO5ZcGRgC4UUd7n3GF23n0JPGyMaFwZpe
ms0KpBL/5kPFRLKjm2xGgd5ZCOUT6lSx8z39q28VPBpUv4Xp24Vxt/z/fM5sLOat2256sKbYSrUT
vDohk2u98pseJwTBE73pMacEqtlT/yPGj5a2ZoSo012dd0HU6kxWpdx35MLDIPEzQ5cWxFYYffzQ
uXYvlWAev5X7zL4aIQKHkEUzqnUg8o6Cs7/uqEMXRwvZW5YAjQWaiO2pJAajTDQSwGBNIQRyJbph
L8LHQ5Y81f7J9USfcDHaYIAfKJi+L+SWpSpjDel5dD0MqyUJ+XnOIG0neKH+4FixP7OsA7u7ih40
vWRP/+EL/2UmXb6xXGCJzpTw7vhRroao5hVz16ahbLzF98DfaKuaCHF0I+F7PvTg481Ebbebet6T
085Sez83YJloGTWLKGSeS418FbSB8lCPPAn+JcV0r1X5fgK8Qki5ObnpmZv1MFJzH5xKd8BwAex8
nykEu+0rD+/gUpMD8hlmB6+r3aZzejD3D2zXMSmLiEHNjzfzgu3TSMFeF0VLRP1ZWsV9R4g2Y8i0
D5DTCYiSaLtdjNGbX3KDqn+IVMyNKOqX5qKkFinZN60zl/XUTSNsOHPFlHJY9xeIn+QDnFrip9h1
g2Mr4mAhT5kcJ4D8CS3YsymoeRfgx65brsGN8kFseDc3sClnKtM5Wq+q1wIL6ihXigH6DUnOy02F
Xonb0PEb5thrNaKrG3w0dDRuJkd1VjaE7t8aP+cfatjlbKmkj+VGV+llXYucQf2mDsTORva7+HQR
pFiOn8lNGLnSdj47LWmz0fOe69zPbWzdmWY+hAcHUPYNNxdGXLATVFs2aV9Q9JsMeFAf/G5D21Gh
ePD1oMqN/MNxkKwx9IvMDrNtu8RE7V2KgzZ7giUdlnMuxAkLAS5prHzZtSl0xDoy0u5GRQ5QIxd3
i1pKdqzwFyPFuLmKI8Q66N17V/UB9tp9SR0ENNLZEX3HfaoHQxkpIdJhrusV6/L9sp2lyzshm+1b
F30GGnerzhIyQkjc//ii1LVFcw8TGbbC96T026kFsoAY/YCVz506WBkKa436npm/vLwoyVLy5ETL
5LmZYvPFRHmkm5M1ivcMVeyH/2vWcERYU8hkHoT9X3m5+/DHfJXeXsxY8RLK7wFa5Xl5ZmFGO/sj
agJoszm6kBC8AaKAhUCl8pLGVoPqFeYhI8xgOA9Nt7KnPjuelgfhsrkd6Vzno7Anb8Zsj5BImVgh
DXHTsl+YueR9hBiqvgBZgvkthvM4v5qRqmrO1GqzAsnbLszCYXNfCvwLvq24sa2JbNct9glo8SEM
js9LJXyH0seC7sLzzxusTDaE7bLCRS6szNGW/HGtW9Nw/TtKyuZ90kEeYkg8Djrj3pPI6xKrQX67
qFkQD6zfEWqdcL3MgIinEcFCLmsPd9BTVwpw4s28pnX4pqFsvcpLaBAoqjIbSKTCA732GjgkIF26
R+iPN+vY1Xxrw3CemeOHYn8zb3e2lQIJCplsyFRhMZBSmsv/dNVbaw9UxGVX0gAqknid1/b4pOIw
Ktl/w/VZ/s+ynXIqr1OPIhCSwaKEfxFG/gOukaepptsB4rYT1H9uC6ysOjCaiwqOQ7FaI4Uz1tk6
cvage4vXWoyvGG7FZEyOK9YKtbYakIcdMPQm5nIFcDm6ml9MzY/+SEH0AnkEp9nKdqaCAyIMkZgp
imG2X7iIILWSDOUvBS0+AaLxMvi/1lqAbltwqHuLqKAEmDcRNsTUL+SxSIvkUf1xpTKE/Ee0+CfT
bmJbhKK1AnKXxXTcPucvT2Un46iKbcT7nF+WDB2XDMYJmYS2/YV75lpY45ZCaAzEU0SYnyeSPi5y
vuRo4BNXnRLpP7DMH/HoaaJtgEusoDMEqpujTCRX1qfgXYQgypl4I7BcBiYQy3z2089jQ+Nf7b1s
iqGyT6HEbdmOYEnN3xQnyJg0t27Jx6Cc/Dv6VeiJ8sSSrey8nmDVyVyWU7p92mJMHEDqQKn+bdD5
i7yj49e7T7/6+0ewPojn5tLR0PPaTWZ0m1FvWDwogYYg/57t7OHGj0HLcvZWyK6nLe+V8RK1jtzK
Ta8Ca39TsFmaTyL/CVN0vC+41VenQKHmzSM53HqZ4jgKek6t4GChd0DnGy5CRGUdOXSsROSdKE57
y8aVcrGTG7qsoor9zcSzNkISBnFzFQmmMnwSW3GNzcfltiFRO9UZP6U28QM7GkOh8s5AWcWT6Rpt
4IiZoYXdggb5aKGVoe96h3mn5suYfYss6n7fjv8c19oxh/QKa6xTWWKhcdVRsaau9xqPl7hFcJtr
DZlikTnP/WzqpNz75zl1AsPD7ONgrsVz2oyL5JbKvGIYeTKUl++dUN5Nmro0zRhOwV271yEGhGRu
tOvD2kVtM+FYfwMlHPlPvY8MfkHCRbExV9XPBI5swyWg14OMOwAcWaOHUl7ePySjMz0Q8Hv6hIkA
rUlwIc7qcnr4KKPaRNntKC2xiavIGGlLc97ddPTLpXbRlAoOijbbNV2O8H6UGKCMvLogXbwol4cu
rvpBukYJthMXkUX0PjwiYZlISSR/zHEaElzNYCHu6lDHYxVnru+HKaBDu+mQT5qD7X3Zy2frjscs
x6Jay1vcjxoH7/nhK4CwgAP+XpPgDpGDxPaJkIWEHefDpM8PXySElfJ2XwhYIKvRxdh0+0Oirlxu
J8l6X4r6emiQL9yOZdmX8LZ5vLdp+EcQTYgN/bjso4HXFpSUA44DusxDkWYr71TIypALrS4gYeJA
03eLJ9/Gfg/gQPu1Bjoxij3pSSXv1v07uI5ZliWMtxUT9++EiXLbZNX6zk51vJSrKycMnVklRVRj
xk/uUbgxXsW4Znpsu2MBkoLsU8MwCct60/68T0CZkYH0t55b70XSB4XOfPc18vmlA4QMWGty32IV
Xp7Rhge4Py6tmhxXGcQzDkOtt/mSqw6MJ6U3J6uZTY419RFwAt14lbqDQVLn79b7fu+sIJ9DC5aq
g+B1/TcSvpbi9SCCi+tmTQg/ar9WdIwb1aLMRoqWI3z2zsU2HITlisZOvz9ZUhV3OyU12jRuKqzZ
wNBPP9lt/ixP1gkmTIa5FkVoTXNVT3zb2fuG2kiuFfillNFL/Q27ci5hdkFTZURZoBFghI0GRaky
sGUes5NjF7mCpVER2XrFvhpDRZ0vO0ztF7+YmONW73t690yNFFlL3aYegF+hQPfdI+w7mryF0wvm
pk9Mc3F0eTl3gITfiWWytnZSzr5tAuDLRvHwxBKIzOXYVA+NUWV9DUtPG4HLH3pUsWViLabkLGZG
M1Y8HIn7YqOLJbaU1p7js2ORF2SozyMl/lPwemjvv1nIIu8w8BnqPEtr1VzRbVt6kR11/kzGeL3G
twuhtzPFV2ehO41tLEK5m/LWxmRp+/BzICnKm5V3uAj2bIPeK05dcOdrOxKMJ/tnD+SZRR/w+xWj
WFJQRv985DdBTgkMKOl705UzbInPuZVVIJyfWNMFHvqxftOTUWGeQWsEMKl7r5cA/O0nCENRi/og
axkfKgeQyVZl+G3t+fonlVdB8GRggJkDCH39ysxtW8ajCRQmdc4vvLy9iZlJJ9Ex48W8OJKWGTWm
CiD7R3AQf7JFuV1Zy8ms9O1MIUHQOd9EYmIIEt7lOgMKD6PqYQMk9HQEzVYPZf2kLA25FsH7jrxv
ddlMe9AWMam6v23ImS4Yd8Vb8AyKQv40PoyXcuTnFTnKnsYynprfnmNQlb49tt4cXPQPLF9x9PqB
aBP4Sj5HOOalvXxdoo9FOjq5AnyyxJh57KDi9Zog1l+WfD0RYxOMo8dY2+jK2cJzfNYi+8lVwP/X
g+qVsA2lusd+dd1L+kAX2SMqyx4ZLDU1jnCPhVTjkchhkLjO7M+jJB8s5L+vdbQoP+GIUPiDGg5t
8rPXH2DaFlAMwIHi2WgSHWmL3jNAZzbHtl+mdy0BTv7F4jEM8CvJNk8f/AqmETNrV4EXcuGa5eJK
hWuW05byFzoRNibcZFYInqB88DidbbEjBSyEXcTpowDirXrc2I4polieIpPxqX1QkwnL8QcOPfRh
veOBHKVzVmyuKdBYeDATEOPQN5fgono6HhEYWIBDCjO35MSJNRogjnzJH8cqdms11fGBgcLTC6Sb
KSzKX8Ijy1LN7jqbUWOIXjsU8b+1ueBNt9Bqn8zzmprx0J5kLvFWKydwGr1fjpHolk9NUwrGIJaw
I/5oE+qt7OAWIxk/F3QT8Sm20HFwa/mX6IPBxhFLDNWSqcWqNZx9Nkn3k1nZVK+jWWIOQ3xU2vdT
jp3H2wHPuEVnJWoOG1a7s8b5jE+wIt591p417i9LXYG4RYYt4VYwdSDKsrX6WIJsS0vMrsqvIie1
nv0mMSZCWqVeia2RCsiv1PdjSqsH7pUO4FlPCdgSKNrm47okdm6nKeV12HEeIW+b0lm1OzxVHVsx
fAM4nhNKTkHE84UaH0AEPmJxRuPV/iSTrJd8arMhY598jk7d/rO2sWEqq4KU/AFqI/2RIBJy38Cg
Wy+UPVmkWBQl73Uvd1bd83drzsWSLVPDewUln4kITNtgmdPxs/g8KNz64WczSVDlvX5V+J9JbMfh
gxrNuTuRO3djDSMwrZ4uMY+D+XvzHr4CLyismqOHaqBQq5OLLfr+XN9tIu/gDUJ/ASfuYCHKvNr4
jMimavIFUnFzZzYi9hzLy/ohvz/mdWFZvkNzqIBJSEU1ZOmRheDB4QIjrAr91A+o1/RTNUy6XVtq
hYnOl2k7XNGcgqQvsRMks+EuP6344+F397mxzZVG0v7zK86vjLGo50aXy9NbbbjG59KEzubWBMW2
+xQGTZ+fb11t1oSsITex6wzD2/Y5kaVEkviOoN/+HgxX/041AU63zNfxwNxt87K6rYAyktjH316Z
tfj/grNKeR+uIzvzoB1F7lcm8O4r5y8k5YaCOeLCcApC8Fxt9MYu4eSW0q3FXvqCwtc8Kl36kWl4
9EUBGDoXKR5a6sCbzKzPy8iB6BDtWObYN7M511wXT9VBn/Zm1Y2UKIAVpFK6UzFSYAD8fHPccIcN
kMDrd1vw0p5h66SiJhqc2YecAfTqm6IjjPIqw6WgTBaN9L7QOzBJmcw4YucCGxbE+buTzfMOWlVD
lElPc4ZWzJNLk4WHKGKazw3AiJ2/AHkHCcBQd5lBZhj3XZrrl1UOp/yZWPfWWvF8Nt8sqa3mi+96
w1bwPmQRaypd1k1f/OygLbcteDPdUagLdZYZE/vb/y4n2khgGn6YgoVWRiLGdqlCr37+DFViOLPT
o6v+w7ngo5MikUsrekITTCRKZ1/a0/+RPmo1DV8Oc03mH/YmfujBHxeEsk2aBJItQAuxzrfGA4nA
/5lpnz14D0tt8D1Sf+OYyYqRvln3zMcfsWeFQT/B6Rb2CxeEhc/dt06SowuaNGawRjodiPll2pe+
M/uFG5bkbIcn/x+FtTfuzvcqoaUg8p3WOcXNsB7RzbUI/AhuF5sd7FTZQnV8vv+O7Zw1YToolBfS
JXJNR2l4gotGtphJ5rNB4L1E235fKPtvLlf10qnS72MdFK7NgzVrC96uo92j1+MVAhe+vWd0tVY7
959CxsXHE8qG1SJRiqRmuRGn13xY/626nw/KjhaeTD7T9KCGt/6OjA8PeTWYE2CGaYrEK2XuZQv0
/9iy/3gWdinQolfqS1MO83IF3rBZnuDc4LxHc+sDnfXKQFm2bNGoHi0BhrBUJAJd6NGfPgshTnUi
CpR7DcQoPL6LSSNpOn9JhkJ9KJ/coNEP7A/K0YgHeyDg+UZ9DcXUi7hUj8T1eGck5AD9yOTrLIqd
j6LJwB24a9l6+Ep1Q1yvxeot1EksooEl/qcU1jVgrGOaWnlnRft50scoPb+e7NOAUl0uxPxlzVPZ
IBNfLdbwJzfZi78QJWeWncO6bPLUvhLFoSRCBn1wFrTeVF++o6uMeNO/hawL8vZ3GEyGL6b5c1IZ
urPeGoI0gn6eXXQ682lUC7CpQQK3CUiXC2Ss2QDJp4Dljm0jF71OgBlCQ22qWJFUY6qqt0l9kGcQ
iCgoZ3avdunj7Vy8+fjabJqpOaQfDC12u+4Gz6ofiwMUuNz4BQw7+eo2glO3LlzJZfRqeyhbfU9H
lPjo2H+2mfZOO+f5FmmvTHA7uHAylnsPogdBsN8nZeVXnyQLlP9i8XflcnDqks5cf81PqVmGirMn
utZAos1rZ+7ARvz8PqtEVEDkZ+hMtJRQeDw5GufIf7oMH5jXW3NQ7OJwKpiPWZBgmMnBovAndyhc
WJzNDWPJbdKcvP1xKvIZWl9i3JHsAC7Lh7BBXtKONfqbEEbDAQBNuiPOFne/J3emwbRG7ZiHa0ZS
NvSuWnlo2e1MGT+mpcp9txEYGxGu3pfvKtAPLEdb5vq00jxqs276Soi1z89O9dpz8O9Hi6J185SX
OSLxUZ0Nw1VeLjWgb5fskJPtsefQXVEHwfoCvcwK8Q82nE2sBHk5AzAHpnO8pSik5TBP2xW7L1Lx
P6y+2ERURTSD7VNjWx5+pdxCqgm6rP0duTGOCh0cdwUUNC/oENur1XWS10Fsneo5HDCjhi06kT0V
2CVkaSaG0pHHSzXr/JORabIqBGpFzj6+zPqGzjRN3/3bD5J+f1KbaRIs02HAPkznTSMPJHmCnkln
J8uXr7smPo5Wc5RKOOU6PIQoGdg31/iLdFVGRRHHK4nDgCh/DO+iiXLIHFwHqYn3vP20U9N+mM/H
aiV6VUYAtLI9Ph4qZhJ3ZKPTql3pIYnRKnetFAYXBkDLSippamwXaEziaoxWcwBjkW9fd9hJVEGe
zfrfLIqoDTBkxSLdV66A5qBWKp4uOjt1fBKpM4d4H7WkQ/uE5gWUXcaZVOPSjNsBviOHz6hC82Nb
Jf1uwRSJst5UbvFjd7gJD0IE6Br6iSCAQDnx1QlrCN1OxPqlcWftRbXOFYJS/FtBmvUVB/tm9pWO
ICXjPMYSmQTGuPUjEi9c+eXfBehBR46Df1WW8Ehm0C0Wfdccta05euUKCYsKUR3jxPzD8/OGiRFK
mLDq7YXfZmXrhsaD9ufbvfB05QvSWA5iYGo5HYgvBCg0hG4JnOC/D92bSo8hG2JqVNceyD5WB5rW
yfmqaC14DNkjlnkH/Tr+xjdj8arSkQVbDR/NLU9IAkPnrmoaHqn5VkpHBSZkwR7+2t2U8Hi9rSWW
okgewuq6tjSP3fTfXzLomdnTNNzggYb0owGpPyKoWYztj9AHer91tbLTsH+EZHHbwUElvk5/mMJz
zVkIWu21ra4hqmPxqKcLvf2rWPevQXaxMCUOxc9Dg6vSRzk1AfysRRtT57QhNhg3mcbe0JIzs+Co
kuUP3Q1Fgt1ENlJbqK/KcOF+3/4CvQ61h+DBCYyB02nCPMkgyG7Bta4N01B6/Ob4O3/W9zA2F0Bj
qfsALR65RK5yt5O361FjjYoCmWr912L3hFxqGZ3bsaL3TiJfrls/LCFbFwZxJLWVmsrCHqaUzK0U
S//Acz/cP37Zr7FCHqfWW37hId+T033ZyWFxkk/VKbpS4+zowZUeJp8RLy8CIymuLNUupmPoB47/
Q6Hv96ZwqONrGRSHYuD6DaXfTgwB/PaS+o6W/VZzgAb70zAOg9Uw70b2qzjzb1463CZ/XgwSrxnA
UzPtfHTAfQMWRuC2ph4vncD4ksT/5IJzkdnA6/qWtaZ3DqJm4egkUMVH+6okj1Eil+3iiPJ2FVC3
VHfN6jzttXiWvLRk0moavNYujIzt5MG4LOYwXNX9hBFSQ+1C5sqNFbwdisGBRjwnXN7NV9VaWJ6S
h30fJOYOWDkKpKbXN72Qe2Nay4lUMDCSi7coBa4W7bKmw4NZftd0suiSb84X7zBkj3/MbTUQR7Rt
qhtV5YHxziqZfLtRUh4daRQwM6rojcEdzJ2iZgjK3PVhRJ231CaDXrAJGyEbCjXVeeWKOZrnkkgw
BVPsv4BgH3N03tZMPbQ5Xg9x00ilxvqX7NVzwnMYiUSgWUFeKw4Ru9cPue1CF7bGZaG+Kv2jAbGz
i1AzqhuQ1SxdC8zhpIDvUR9BcjJw+9UDVJ3lzebmnk8iz4mkMwLqjpsEaVlZIRtN2cH8qm2GBUgj
WUzRS0Jx/aRZOgT/OhJTtxQUSI2V27JPFByyjSYtAET/wlYJGYvQYhRIz5JK4VkdpmgYeeEEt/cr
MdB6bJhesIP8wR0JGvtjmYN7XTzS/6OnZcW13ePaA4anpIyyQGbRtSUO+8pVmFis0ZTamB0GF4sy
CqdP6JqClRCsZy57YB3I2YGZSfbA1VGZfOrk1CFSvt+jYsUVi1iMRCzNoE/u9z59mHKLADfc8hMu
CGIcvMCGQ6JJdbhyPJEsJiiesWZoc97WTXe+7NoqM/HUXE2xa1jYdJHBOTWNqV0L/WeoRyRf7W/q
xM6iZICnDwkQ1CctSR9xbzkwMXCrxY1Ol2quMaDaRNXPj5crK/5ayTePbtrGOvDcdCNwVOF8AadV
DHfHwYuAIEQtPlaY0sEd/8WtspZEXRWCX0ixFrpmDklAHxBl8/6q9aE2dHDVUaaX99NUjfeNGzSe
/mo0khTK7i+Ulljvzp0QErgiU6eWtQsNi2D8AW9Fxz+iNIzFSg0bYkprYptR5gUlthi0Nuhw1cRe
N8id2Ct9qhc6yMjk/d07+PfDgrSq1MXtJvyRjC8mlFMe//je/ftF7O7EweEG/fwZGmMw4Ls/iGEu
CDCcuZrpel7U7YwLN6MiT37Rgdn9tqh9zaIid7NTRtxE7QhVHX8NlnIWkcyfJMTZJ4U+KXhpJkkT
vz1ckLEhFVzr8EXI+FYNBMdYtbICeamqX+metF0557unXMiT3oeQl+qCLff9fZ6O49BF2KgMgDyY
JDqP9ik8J2BjniBqaFIZ0u+B40Vu0cphSgWrPihErgqmZZ0lcJIYoGY4NEUCaVn5G3DL87QiUsxw
XM3ZNfxXBIseQiIv+oLdrf1VDG0mCJVcBr/7t+R5cCW/wwpkQ4Z7lv711uS56jIDG663h6PkHfHq
oB1glhcXtfb3mXnLjuec2W/ggdLaQ6Y1wlHBEmQKD01+wZw0oHOjhrKrHHxAdU9qizcXhGsOmYIX
0wEDg+MK6BQiSzwWaJmOEjktZIPdnzkPfOted7KVgeFFqGzNtihJImJjogaHpfppIgFk1ayIteKO
2NeqT9KPyoKmeF7NuEhorBGg/QvMyxBjip8a6hNim5kVUZvnkVbkqL4KFwrC422E/yyLxS8buomo
qz99/Jto/ODuHGznx+NyAAMcgwEuYAAjt7QJ8sDbFj08zZ8FxfBqHzEi4ISD16LSOgaJEVxASe95
WHPokuYKrSx/n48hFTiHQk2nzYsB+CEUu/VDizLS37FgvCtwa1Pta5n9t7rkY6dFpSoQdBjaWlA5
+AVv2gaOzFrzKvqbzIXB8pdZRkXJu8Nb+EM7NzIaoJz2C0CG1W8vm/Ooz5+sECP6Hvy0CdLrFbpH
WAcyTUVkp+3rsrQfu3b8h3mjYlyHJeU6pUCzCsLrSSNCV7UUCdDXypxPjq//SRj8l82xZ1W/2deh
bBf1yNhiviDBrdOOmzYdBRYrrAusE8Usf1YcKg6G4fYIWCkwqtHAfupMej3/lruoykmxKKQJ5syy
Tyc+E6sZOGdPOB5QIw2Xd4Owb8YvIqYn9Q/21oY2/0aPx6RlaFUY2sdGwQ2fLZe/iMMy1ng++elu
SvdanmlURCIvtJD40q09gxjDKhZYWoRukqYQ41CMNSEVKWVAU5cW5ObRjCzgfBWXsx1cwOgOx1ii
FiF3eyQRVbQQVeB7m8lI6hHwmKyPeNFFiQ+ri3kKxSeTy3hOpIaPxxO5u6Z+u1M17iV8ROiSVafJ
UwWTCNlms4nO8bI4n8AeAQIST1sUIMY099WVKXwqwK9pxpNwS0V05WWTAp/ltqYgev7MDHpAyUMG
/+b0p3IJaTZXAZkDtXdXqSvcjnEIL4Xk6nWZK3IiRdUlPRADeIG/pgoPvTc6/OiatwpdOutIQldn
dUZx1ArEoJar/T0OexH0DiRi6tZycGoMhqjb1Ycj/cmyTx1GjL1E9Sny+yuqRcO+nDzxWLb6BUTX
Svuq1xksVp2PZMtnLfde5GDSzhB+IBbQPH1vvRpJBFZkegfrVhiyZ+HqpkCB34pVv1Vkbyhg6wLr
kx8nIF5ZbrIcFMcHt9ep8ZohpPmBoUhUWHHnxlmcnIKAS39M9/XR0AzD0To6t3But3KmNhJLDpAz
TNUWRjUPOLO0s5JiEV5Tr1/zDmXhHadq2hgdShs48yAx7h/m4FB/0YIktc5iZlD8KgVQ21aNd0Li
kaNNz2xZCEiczRm0bESbv+SdNFvsy9lsARSB8SbjmdDk/UtXF4cgpdgFz4J4eY66lrrWGtgNB+qd
XtT8gyYonU0b8SRhh52mCyaq7cVBNylppue4AtNCoBKj75cqgdIV3ZZ0wExRFUlWZ1j7cQaqANKF
K+HReAmTrdOKNS4z/vnO3agtwT0v/w4H9jtGlufVMyMGMBq5Q46L6KSDBbUTjEvF8PJHCuTlXXSP
k9/ijFDET2i0KEiuI6JjXdtG6xC7NmJMDpw43J+OlUcjYP0Tz0BT/oSRUlIn9kc0MtXs0s1GPK0l
D08k7vdIWzvtFrqaOch449jXQPR94pLGMNvyGmDqe4zeMFkRFMPYI3mATWQMautaGYz2CSZck0pL
iujX6Y1gsn+LfAZooRECzJGbCVPYzUi4bvIukX/XEGT7AkkpeQnHNOXZMec22wqWts3Eh06RdbRR
IFDTLWeyTcA01SAmNJvVYZywbirAFsQXuuP5dY6ljVJhPHMaNBqdGA4Dz34tiQz8oQKjhrdK769R
oeOCD4vVOBDFcDutGiNNQwzm7IXG8DWvMITIJJF5wOy3+Lc03LDnAR9F9HM0kyo9AERtQFT+0ODi
YekxQyup8j7nIUbW/qyJd/mm5+m3aOd1+lfnd1BJoJxq87OW5NewkhDRGl8JhQhIRCA7YI5AoeeG
BtR7ddp++11nx9PMeg73NHaUFGIsyn6uo97hVQGvdolQ6hVLRINCQVwirVMOt0vWtSvVGUP/BSAD
ilh8nDk6KBGPw+olV47Nzn+zOXSjhghjU/A+ztE3EtrAjuGpIJJlcGaohp8IbcXOPU9wZ0kgtQxQ
gVHGe2DtTnh6wDiQRYXPHFfzq8bOap/oqxDsLB69a9SscrRyxSLQmK7J2bOMNglDMLr/mXIyTGr9
9biAxC+97S/qIZALmzWOA6hkzAaJQmY7ACR9PswsmX4u3/1gjO7NxIuK/R5anMXXwAlxGBWTXLVU
vKmf2rUlxkbHLTgUJBa995DieFNYyNY/YjCwMm5Ws+abIil25kZSHgGwaPPOPl3Pt/7iH0WhpzpA
nwXGCoxC1jM5/sdpy9hVY4nIGmAQbFoVj7YyI3RNT+iDc2HmDhAPShoUrsi4nL13VeM1AbtEfu2n
Cwak1HOWFvZ8XSd3jKK/08trIgF8BhpOrbbtvsad3MazMoPjiQntawXFihR7g6Rn6mgjp4mgB+Jj
01v9ek1BsmWDruPIRkL8r6ooWZH/jEebC/q4VCP5Pj/cyIiDJ6+wR1bkGdT7A652l4WWWR77tc2+
o+QUODX5gPqB/erk81ds/6s5ZJHFLAJxkXaiWkLkhByCqjYEmux8BdqNb6UQx48dys2qoOLJwHhZ
X9zEzH5EgM60/G+CfYeX7yAY9gII5fqu4BEcC6K7Gt1wE9p6ZUTgFZ12zsHlVBXFF/6hHHNk3888
H0q1/ai31So8WctXNbThbjFVhm+51AvJ0DgYmN2sZjfCgYgd97SAot+1brmnorQaJnFqkAOGHqpU
608LiRLvd66Lg3ZGXYSvPvyNx6SA4QP9KD9fKEhqsu+sFvOBXea6lLjAIE374rn/CGZCzbapu+03
cy2UUsRid7R8E/HVzFR3zTzMQwZYaF3Xoa/rCpnAz5q54xgFMxUI+m4Gzq3E789PzUcC5zT21Y39
w6HAKCsIFpe6ngzfm4o08i0EZb0SqtjxST9svrWEKDSLKt7MzF9CFqhUp2ouY6C3SKG4wS9t1S97
gfwVGQqf9oMkgCRdKGKiA6kpNQ5P99fyuWVM8+pyfHa8XGOBNFaQtVR3hDRW351hFoNsjUdAwKYP
ctMDTe3bzYO2ohMhSTJxr+UkxiP5WJV2Ee/A4LPJXxrybCdyBwEQffrt9yE0q1Ay36JNg7Bi6ffU
3FvgwtUZVxReIQNkcsjfT6z6WCOQ/CHNJdF/67JKe4+dVN5APWeGyfdVfN2CQVqhJeciKsjnMueJ
L95Me/WB+3bZTJdGn5QHhDWDUUSSI3n5udpG+doZfdmP23wdLuEBs6yhbzjTgq+6ZFb1UuGKs7Wx
lRmt73/vtMeS/Jt7pQrUlS5YG8lRMkuI7UPqjLkIcIOHdsmwVm3p0waB1DjsDpuWsTHxaWi6lpkO
KQ8nKpN5prJYBCGPEMoZ2mYgM2LUzHmd2gAaCI7BQz3KuRRbPtP4h3uUD6VVwPaxEHTEhw0elmos
oVIPg+5J3RP83qEJdJi9METJ8verGOJVt0c+Qel/Uo/55Y92vtwBeaJLmdQlgWnM7sYbDDYnviNi
MJ2eEydAbrpLufVutUQ+tYMMCEMrvEGpp3HQQLgFIoQjsYkK6cRtVKvqz7kM/7Bko3usa0864Sgv
J3l6PedWtC7n3pMAe2atwscto6cu8nnrC4n22fkWgmXeyUbC8kLnZmUjHfBxA/h8kM5+RR1MUUac
tfDFgLBT2yQiKJ9IK5/HDAADMyHPIP36dH62Be2aLukzqwtSzU24JQuX4woPaq5TE3UJpcasrj9/
l6Uic1qhekeZBiOZrdXeWKevJvJSXQaRZWk8bQYDjuU3bhS/XnuenLjp0PqI9syjq4fNGmDJiygj
ZT4jA0n4LO60GwHfydiOPOUPd2AUpG9TdexiCO6Sfa4mPMcKWPrqQpJVibgVFUo7ZfB+Z/AUNDfk
baXEpM2tRv/n2azCb4Iv2oFxVTL63KF3e3wrlO9PyuNO303frZokACx6UOZuzvjhlgE2eRP7i+ub
mJERCEWynamcpBkOYOIZdogZjnSiNr7lPTXHjZSCNIivyh9WGJuuEAAKuVmJETIIvO9OfetIX8MS
6GCJvXgphzI7UEn1uCDWHIsKI49nx8D29qq2gv4RZSGplGUa1DePCp7VCVYauwKvFQkTUj8ECmeG
wtKn8z/Ya570Igj+e5/r0hnkVFGV9m1nT1S+bCyprfZ5gq/Ofic3kaqCJ0depWoBdmmCb3JZUvYz
vT9VbEB3oaTIHnRAPYBCbvzZS1/Y8mU1dkU6xRpiaYye1AY0RF0wMV5uzex9TVEB7WdtrxN4CCir
9BWdbEtxctr3PWN7FVGkwKdpVtHR3eBJLKM=
`pragma protect end_protected
