`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
aaWX+RXW+JYYxLcaJSDmeQbrMJiIG8RVLefhQMpF7ok8yt3AUm9zAB3YsxEY7DVnt+0Qi7cyP0i/
Fz/wr2+STQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Sag9X0VTvdmkzilN20OH58Du9EMZQ5gTXlFiJHAHASj3LslWwaG5zS/uF5eD9jFT1EQPrIuITcaw
KB+c6/DgdzskXejqpcM4FNY6AdDA6baFoWYxzZUeAUKnwIiwdOP8h63ejS0WyLm/AkvO1nYAUuiB
xZiFpWTO7SkEN8sorqw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
jx8iaN93qft5c/Hgh17wVfud/KVXPDiEoE/gCMCyy3LV7jURoNrSWyx2OLUdD8ukOlS1hn0kBPu7
bYWC8mw/azUcnmap3LEwhRmSInMgDcFKeS1Lq8O19x1lpRvsewqkgouJzcVIB2obNMQ7DnlFlC02
jgzC/fa5GNMpraEH5SyRDR5N4rTjh7HJRTe+/oiiPyx39H6797vFWIf2SVQYcjDLM4UhfB9yPGNF
aTRVeVEtfzDrBQUjUBsrsKzirwdGNFwIf0mkP10DMtO5lj384IWKEzJI1MrV8Dj5n4FjKNzpjy5l
08Q0IvDYJJAXeNZnRgRbB1VWikDoIPcJAiknmg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
DvGBQ8pckqaDVW4OigHVkkf6EgQ9MIQSm/7Rix2F81Za0lTs0bgtaHXv6/nR9MM51hW1f5FYuY2V
ypNlhxpCXEKLBEkF9pCWhZMYheSldu4qRY2OJC+mFSTDrfaYEgD3OLGHO/rHCnvo3V0iYCH8SvWX
CIUPQadkro8JnetXqTwuAH6RNujz1KFkvdXvxQr9j5zEMP8HlSuf6h/+L1ODRCiIDsvaZnr7nE7I
Y8H6AQedqsGwa2rRPlHQpdL1NU2IbY4SuQ5LV0Fv/00yFwTbepe7j7t5sx01vhSPnyaNK1Ysives
oVkWncMiIL7BmCfs2YNArxhrImECBuDd4w+TGQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MGHIdF8GGfDSJK4lEmSE/nyCK1MX6mLVlTuBEcpJVf8NyQjT3Ti8+eJ5UOE1O4xk+r7vzOASf1af
VXfR0sXtqPVjk74QuiZgtFmYuU5PLfPrL53k2kpKTDDxLZn2lFTlWyWqMTD+csmj3kRbRT6hFAIy
C6+23tsLFw+bWE/hBcppE2XlV8VhnTDVVM08bBmCpWmIluZrnH4kms1KSmfWZhHVzVWTrgIkSwMz
ScYdW6ecYu2T3PwHjlrJrpCSKRuTPOhbz82d5g/2wWsF3lkCTDN2RC+CF2rLiSoCkWAUJ4m5CGQ9
bWGMsW1OJGvotzPkVSKNKZe0X1JM0XqQMN/AtQ==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
GWgzgUVU1lVfSOUuslwLB+vAEv3+rZLg19FjytWV/KKdSO79OvGYuOu+FfbB3Ha/J/HS0Dw7VoWi
eOeMRXxZCU9Z4fN5mvv8iqET2JZrsoesPM2pJyFRvHEtt/cZ7vAWdrWdJxcFMG91HOYfLy5SMeLx
+aOXNcavImdd/MowK5I=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
q8Bd0tZIiyd9JcH9UY3+hAw6aT3ce22Nj0E60qDMBWsL1MiNmKwcJP16YB8IlMiawH8O0WrED2Yl
kHLIV4jNwRUlRlpw03IPy3EKIJ/2eXWHfVEhAsClVL6JLS97Ubf+Kp33wdrMhheuIUvI5wil5LXL
YnXWiETbzSDVGvg85l/Rg2cDHKJ4oyztKH/oXw2qLARogZRajVqJvnVBAUP+M0JfzUWw+PnH9mGB
dYZgqhMOPExtIWTxork6D3lQ6VjThwJpHby22N0fnLSFFAQNyg8u3eKEpVcM2YlkLJGVQX4Rd6xo
49eBj+86JemxoZJVqGluCaE+BR61Cws8RrWlOw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AX/loxH9jMcRZyAdg3lMjqgfvRpTRm0dSidHbgXZc7q2sp1oyE0CrcCkpw3blvX4/EC/I2riH+9l
+1FqxWKE/4MvU790ATrGbnIK/qmKBHpL7EJtHvwnzSOMalYr73o2TUH646NjjlbIiteaYPbaeJ+z
K80PgZ5nvxBKeZeLpRLnTdgQZKMBMoNIu4BeUPfWE3UYgmI+c54aQ1lgTkNefYtchiHKStAhJdKR
NEKNJ2bMR/F40w/mWIAVh3k2Tv6d6deXS+e7aJ1PCXTp9u2niOMIUqgKyNj95sK2TAw1u5g0D3wo
v8SXvSkY2QTPNkaNSDgVWSpeCT5f2pPPt9I57g==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 432)
`pragma protect data_block
vqBPi/8C/p3AstUOgdZK1QiJRLUIctOwgw9aqOtyVQxupVvg9+OfRv7Gf5z6RsU4sX4IK7sC7Cv/
7aiy/o411DfcEPI0j5bKMZCeVzxSLPTMyJSyf5BZq6LmJ2cA7IJA+8naShesRdKc1j6Iw3FtIOch
Vyae1yPNggixyIT13qLXiNKHJH2uL6ev09QVW+4c+X5UUj4br8Qz625k+y2SlQi3Z8kmXzxYiFID
up5hxfAzsF9mXKAM5Z77xM0kFyGgpK1evMaP9Ui5A0QYsq8UBfOV+UworKEPlRaBmmvPls8XrzVv
fvKWJnG75U/eD/2irzHHvxlvFMe4AR8qdDjRKzyMW0JQJOu75G76pNeyh0YgD8NIj+I37evHMHVF
jeCi5wkcFslsm5nHTD/h0ZcHkfZY+yf0ydRbgpDwzf54MhWDpFZbd/PzcQ981eboJefNXirfBhaU
4CRCbsJfo4Kt1taQXsL6R5LnXgYKZiT15peqHaWXVi8pQZUjyfTRAi0vwlOEripZdITsuYdWaJ1u
BZ49jfGqTJ0UOywRvP1Q4mZqgG5PAsPbHY16so0BR0qh
`pragma protect end_protected
