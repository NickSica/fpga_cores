`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5IlQqxgcm6JvJjWDD6TdiVcpoUm9UV2fn8fKu4zaQrqxt0knSu+3dFwO
nJNhXa5YddLGKTFIwIvB+olpChL3bS4BA7zG4aUgZtiT+I455tRkBYmGJq5nYb8CqXKmdo2xwb9X
VxadQZqIY59v+gFv9e7d4FwIBPTbzEdcRwW+bS6QerrynDvrU7lUV6RxEsHuk1ePzbXIshyeSeKa
bBb8GhOlkkPrs8k9p8UHPE5sW4ANpGH71ZkpWy1gP9fUyze1c4Db9cr7w9owmO2Lvc5WKvuVzPDZ
bKfg/hfE2FwW6PdtVJ4m9EzjAKiIhWAgbsYgJr1sn+wiOjntp0W8OH/bSZk4RFezzNFsTGjLbBoI
LCYQTE7SsnioYbWR3MAJG59cZ/BmSJGdO93mdAzmCaH38Gd8ei/4HkWeuHxyI+Wp53hK2B2qQ7Qo
X8a1R7aDuVpTzGhLITIoZERwWRQM1iBlLMCLZtk9b+Ws8qd5LxuKFreWTiIEaI5dnz6oKvwPsDMP
q43DuAbfnZk1/VSyeGJ4o+CMxZ6HlbyhwnyKERchJ8VOQtZn/i5L8ydN4bDJ7ekvDsgJQNsdps/V
j0YeTK60W1Dh37sYkwQFo+OXODDnw2zkw9UyEQ2wV3sQ2XNecRveWP79vHhaH2kbig7ekC0Wq+t5
SzUgHZMlNqg8mfVVs9ro7vi9DzEqNG9gvNMuku/iRUbSnMODpGscgHaJ2FD1hK1tKM1Px+Y2Dy8L
2wahSkk3/0agGQ/Fl74fzPqCsa8/eh5FJVo4M9hleM34cFFxtxiILiQu6bGHn7T386PgpZXP2Uzi
SbqV5ybtIO3BIJ4Tz1i+NMl88M8yGPw9BnOR9cK7RXSzf/IgE4ITW0bpQJTHjX3aOViP/48Lz3Dz
1poR8FxgkhJGyz6jl43zM9V+gj3ZdsZaRYDZyDVNA0fWkkhEsudgAfeqS03N3k01kwfBLOT7E7SB
btn+/DI4tUyQT+EJo90jch3LF5Oi1DRnnsv/VkK6d84oNXAkH1libnY2FP0V93IZm26LUySDVBmt
Od/u5B+tdOhKGLMkArIr2FHS0Wg0iNzywPydKi6chWaHgvVTcnuaCXPUb2YN4m5ufws19SLi5UHH
79NnaSrS26o1MWzFnXDMQSzfIwaPS/XC9IwzDs6dc2tqQdWdNNkRYShj1sF0B8dIz+QcOOzk0obm
zaRtS4UUFmpT1n6QjLcqEKaKzhO7K5qFX2L8gSTiCUanoZORAM0QVEJ40hwi4nprLnU7eIFoECFo
XfYVg/H8gHbqfJHrr8zl5C9lKgXy0LQhlV3tHVQB6yTJI8XUM2MiSKHwjmE06n8egJyX1T59V6BW
/+kyZPmkhfWztdQ5n3iMwCQkO4XI7h2TuXrfHHhGskqMPiPSgyLTm3aGUw5i/OiY3LwmgHxY6d/0
De/fbK+yRvlnIclpKwZLWI/pKlmjLZqzETMj6RMQKN1wtR/9aSCF2OK5jeg6YIvElMcHL+3j4nrB
ZdzlM/qHvOZBjARDB9Fr8As/iRYgV5fDelQHcHvIf+eiQYsA0zTPFQyFYzb2A+JXeK1uhAuTh9lX
KVo8iQ0yNFS6ceOQTRk4eCvWtYvnZSVWMos+CLC/aXefCtnlAWvX5fpDfcwWsLoXAOtnALSovvTN
0EaZcrdijZCKOnX+UZscCfB4j+bTMJ1JjVN+QV/+7hfLvtKqQGmstr6IvdiySGhwEyN38NBOR4Jb
VXeWBP4D4Rm2Lx7/GaVP0JAOpts44fLLguoo4ddU+MtDT3mwpzT2a6CeHTank2khwEtNqlxkz6BA
64jrMx5erro6UYD4olShDbOh0npcBvj+lRQIx1ZYtgEn1Nt+0zuPUE1+dfTfJ6N0hbErzlIWmlIq
fT+tNopSFFZK7leNKFIaV5xicwmIZUOzvsSIM/HSlBovZzk79qcrVmvqRdCPfhX8Okpeejn8qBy6
vnVQb9jhdfVVmKx/HpGSvKyGAhGk51EsKSHJWTJuSy8Hlyn+RhYbsKQI+70ME2Bf8bM4XYxdJz9X
N9+zNqdQ3f0a4wQMFIjaUyp9dDyJS1dPsQiUVZK3KHQf4ZYZit4WwVEWYIh3+YWMRgYz4T3M4Gjz
fiX9b4dLvrKFh7F2/1V+ELezxOKfs+GSdpxrUhzBVkb+1e2GBnzBzyUIUE9dlKU17Q0ZEpfL4q3S
e6A3GQN1pE8tM8R8g7/sZwWOFbWnsVe+dBtfHlJ6JRfKpPAXMUNI3/c5BroXARQkK7mXlkiFzs6Q
h0n/0GUDB8pz3jPpGaKx0qlPfK60GpPYukDMq+yLQMbCIablAE1J14/MCZ/XZKFIt8bAXh4EaP5v
MSpGjbqXJOtgS33N8EqmgDWBIfRP2bfBEXnJM4OJtC+fn8+zzj00c0cmR/qWzxZ7BrP1uYE7VUiC
yjwfhTdPxtm82oUmtwHLl2pN2HMPOxO2lxYY4QkKqKArXNxNCNeYPRjTpQm2z0pyau7DqCDPUW6F
OXzkZbmOI8SeE45XqtJrBxDR6Dej4KXQSgYUZZC4zX5w4qu8Ak3wvTLQFRUAKHIaacWIwaSbUmp9
OprGTinkGr9oA95WEEX0eS5LGKFSnQ0/BSwWCj6T6+04GoParw8rgszRn1+gmK3h++BQsFxRjCDn
FM42prWV5/eLSabtn0+IIahXiQCbo0A14wkWppc/CuXvCv7dxUWz1HcLIocogDz4vcRRt6ivixQM
VWRBbKRwHM2CxtUE+Koea0GmNpzx6ZL/lzONYLu5yeDW9A31R0Mk2lIe0zLNf9riaV/vkyWjkxMy
5/r4KalFASrsjAWpwya/4Y+QmSxi4pWQVn/smkgOkfZHubLewWa36cRHNao8uGhafWTDh/6f3A7D
ApMFPrjCB7MY3H67tuE2kZvV5MzfvSgRGV3B9jRmsYe4xD45N1IIK7hf1eorK96tYzPBQHJt9N/T
fcbqfxfj4EKUMlRUm10u19C3oc8XbtuV6cloysfWHx3yI8bxk+99ZSGr5tlLycKebjXwEHRcgf+Q
oMmkyRVkEIBk5x+8kTVSFVqJTzq8Uc7mPpe2tPdPP73wSW7vcM4xPoBieSW+98T7hGWu4U6pGOJD
BzcEppEMY3cJBBDwf4yV67Q/JXumjRn3tskAiTZqlOuKht+KPMxygFScow5ttlrRpGZGjBDvzj4W
b1OuIvljE8R8S4DVL1iYpbbuF5tbseFoHJT1vCyIwiKcWyEqpnAW56ypmVfUHx0iO7tvyPPp5yso
nOB+cmtr8/eTWW9FcQoeU8oIcwv+WqXyP3whJCmqvAjSA08ftWWpW4MTIk272PMnefFDZINhVP++
WyFJJ2MWYj7keuc03cBb412qy0/vTuWaFkIcJL4YUdGRDNAMm9xfnw8NcpZUHM5J1k/3Nh4y3x+K
bT6k5kzPmVBu1y5i/Gz641GoOrchBHk2Rb6WMaVt9lpr4SP+Lh4nbI75CzkWUgid+wjWRFOoW8hM
Aae/X21r5lbpJaxXDxJNweBXjCCo42IVPlnmanvRvj//tjFupQYf1kTzhpaqCZ4VNUkpswsHx3HG
BfLhjlZTUlZS396uh7TAbRAnYVcDINeZtJUvcJp0oSLO4rTGWeDyGMxo+8fsVJmytwQfmyK9fev0
W1/YIR50YBR9puMDIX7hIukrh1dkiXRQwD9xoOd+oa7ZsQs6vwrWiziuAIymQYWMJgVhL4UN1S4F
1vDv5v+eIGeZzW2ZwLBEhEaz0ZXmaDIsGbc8ouO/WXUbtrmhIg9Aai55VIRxS2LB7j9JgyBAOp48
kp3I+rp3Sm6PRvVG92WgK2hiKguZzmnZ+8mMsaaCYTMmpKULqvbbT5JVcFcwNqowLJU7TyU3aSJ2
UJQcsLIqWswSJYGsOH5mEvih4yOLXnZx9+OkoPebAaB+sJWW/fY6jvv9VVSBswq/CMcN4izdjFqW
ytWtaw1YSCnFb/9Ftx6+b+2wVC20iPtfQ42Z/tlIvAd3tVTya3aMOtQ6JZeey9fjCGlEa0q8KTTL
8HSutPD7bVDvkUsXYQEFvwdCx128uTN/GqG4zmAQsbtP96rKqx8YeimWTIv9bCghiLhEAOAKyAcN
wuuB6xyylRW8rUmzZe++K/HTKPyyWaHeCzntUAFFz/Jh5B6L3NRo5u9JhJ/niAs7RC8THe19RVfB
zLj1kozR2+uGRKE/vC69gL4zjLNqZ5WlZCJZYR5tkl8ZOAUDRwvTwjrGJdgw9XqoXx/ty1Mpyyf2
mG/ZiHU5m2aZ097BCdO7eInQ++Z4Ul0r+4es36stORs4T00p2Opcnk0DPo0t1Ll8Hi8/HfJMAq9V
tl8M1jXy+OTg3m6Uze8g/QhqYiswrE7c2psBqr8z5mpX4V5oM6VUzf6s3z35xjBUfICZO0REAUJN
mas7PYLEXME3jjblC0WjISG4ZETOr7TgVs+dUtLFHBUYzAoXkGd+8SD3X7ueEqxZgUtyWvGBxV3n
RD/BHCEuLS0geXha44uXFPSYG5aCClM7nF86YeuOtn5jNu4Q8MRxMNGBNWzsnj7+c7HzhIGgfN4Q
Dlts0lJCcrdls38QRyY6iqv0GW7zHLn0HhpKvPXWy17B2BtZRcZa3IFtOTX718OvLX+WWc5+BIhR
X3Ct7y6+4cSWh5qDZA1XtefAHq4BCKdqPe2A
`pragma protect end_protected
