`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
R1WqgqFekyFBf+R1EmSjRCQxUuOx6MT9aQyodTNNebOe0CK13nDxh2Wir1luIC2E+1RiIa720P7G
30ynEHVRjA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KNMY+1Jln0fE2Hw6EJV59uwRAjQ2BHIWVdMuSpeAltv11pWP/JZCrd4z/uZcVTngSRY8jZzhCZTQ
WJ4MxCfVaXUWBZm7mY0qLw6qcMnyzincQFakqwRdOx84IckfsGjNGJ3OEjUVkf7dW/J0o6KJvGRq
A/P9gVOYmGcnWb2CkLI=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
sL7gG3oizEXkzDHancu7/45cwKfdv4EnXAdeK54QMEX/eoc5P95Q2IxqcI+tnVljSH1drXWj0Eb6
Of0W/iXPKZ8OP77HA72GpMs5rDnQtlgP3rECZlxuTJ9RMJVfJzzO19m/vMWeqMysX1t8PW29rrsf
0Tqwcs84OG2uxBTuyDEWCBSCU7Yk0aBYU4VmF2rkELqh6jo2Q/udlKIUXrwoYSdX0O9uon++5ahv
mjzu8SGK6zkA4uqzG9ghLIe8qBE6KYXQuzvdlMdTVdy8eHbCbzVTNoB6j51Qlq+S5oMMSQvxBaRz
DIAN76FuevwCbX/XKHESsvee5Sen235LJDeW6Q==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NTwqMfOwske0aroynepwGO4Lz00SLylJkTISN8LAcq5uE8ZoeT6aFHS3yIuZsI6EEE3s5mQQ8Cob
RXh00Ler2BvOA4K7lNGJUpMzGqJI7MZao2GijCVpdWL1r0vSvaacAIY9nlusgQmU63NqWs7cQx1t
7NMmVlpgPTHr3KxO5lMNWR2EuXJ0I0zOxQbbrTneEEip68PBGwJFyFdSjQNe3iwSj7O0u1NlI0nF
01F/RGHelGngznubnZikT85LEu94GTbx+WNlMlaxWaxuIaRvhH8UG7MPhsxH6x7sS5ZS9GHBkFDK
gyo/ARDW7a6331M9HUgGOcgw3trs1/Klf0nskg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
F0eZzxJQxbI/Xk9S9oAxZw5Tpi91CrcqL3BrQB2lyqn9Vl25Garq+8JIOwcSUfEju0nEdI9Cvd5l
ooe0NMs4K3iY8tnE+FiNZhFGnmyV5djhXaAeRPiaySzeXAc0nSnoahW36RgdEHyPbHBrMfq1pT3d
S/0aa8cloJNV0EZcGFq/QrhQOhscPpDi8uk4IV75ihx4K3Y6D/SPBsIijokh2lVOyPsWt72NbpFl
R1J6iXczzSEND79HNenePfXgQ1Sr+h8Z2ujGHirxn/++xFCAHxWZmhGcFFwVO7AI15b3pfNiyQF1
2SACCg7/b/5q/JpHGBLoFY5e10UGMoGkaXNq2g==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eShHfvBzKaZ/Wp/QUxGlK7/6Td59dAgzaJsrKOgtjc73r+sFOocLpKUK8YR7XmM0pkfLOBkjrXYq
jGiy10qSwBo8l2eE17VZo8T9nQ0IB2FFGgVl0zNGiZaKSzE4a7K5so8c5gtUyyVlyHWXKqYAj6Ro
NzUEnqMqJPppbTPQbvI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
VtDvfrNdg+YlmytFZV1nO9Ch/hNzGllGY3c+wOLUGxBvYhloxzDDcAB/7/ljwrwghZilvxZm/DJg
2fzdltt6rugwiyCDZPTj9bYqZhAAM0bSdp5YpZP0gTz8EvbCxUo8+Op+ufZee7A2QX4lG973f4tu
FbV42AkOjECD3RCU/zC8zhB5kCMonmYQSEe1sGWBe2+Ga49sur53s1VC1GSUOY3PQLHNqtwSq2Ra
owo+cSlmwu7mHpq7nDvHG8vWLm58VKt4pglBRfC9BYdbhmSQeWT4IcMsVz3wzwUMY4HmFkj+0Htu
JAA3fKLFH4/svF3ilwX+klAmiEhOn+ftw2QOyw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HHgo2A7au8S1PE/PLf9TgssZhqFUk1LyRHoBPoQd7KZOhYH8iTwJV9W8hjvxzC2Na0peqSJ5zF18
7DRfKJ++XfNw8OtnyxfjOhMGRjIzpk9/xlZOxoCpZPFsl6WTW8CoN0RLlh22HuIAeiFQu4jBiY8s
f/eG3F7z8aDUIS222+2y8Lc0ifWDx1YbNoJritsavlDA9L9WOwq+EXi3pvUCyXszhqfkMn1JVCVR
qUhUx37i3M4UJEKXpk5rfAol3dwNa+jlOtqwiBj8/VnhZxY2i53S+bX3OP8N1Zx5wRoa1UkpaXLd
9XQOggc4VKKTgU9CJZPlRk8FrwN41qv2G8xfRQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3152)
`pragma protect data_block
eeCl3Hcc/V4mGRBHBrnlVHJbOUqReYew57PSt4XNTtv/cVnC95TSQLlFiNAG7mVJNYxV42w7+NAq
hnUTIUlB2M+iwMZtijptu565NHr68aJ3P1otL10ii1sbqM71LWvRHazEDLbYrdurQ5e4W6Yd2z/4
AAUXElRery2ITm2MmgTEU6gRv1sBZCxFua1aCrxWTz/IVHfzcA/gU0TdmG4D45wn3S4WLixmevSS
uUoBj7qS/o2aqaLJTFU7AlK75EEP7JA9/H7sdMUWIziMycex/E4lOViQmyry0OwkRBEYTfvAhBCV
SEGmj2D4vEyfHj2MNM3ifcupJ71O/gkmv45gvSEuNurkfu5jqSpq7f9TxpiqBRNGk7XX1yM8ryYX
b2/GdxZU3X5wBg8JCtR40UQOv0DIc7udxOuLvk8VUb/Nfcavp+3mph7sOxGJrLkaw3Lj+9yS/9PM
TBpCw5d26qlAhEV4/s3kyPVmocO8M+Cmih1uF0lzHqwl+9mfdHp8bh71Mi9khH4qw5IMmoJv68hi
h2+vBnElCJK1Ishb9iMJgoxmvh/DN/jlkvO4EP6ZcXk8zqfyjvUeG1ot4mQlAB2LMw4LLs5WrQyj
t6JIakPAsRUFkoMk/LXAHgVq4BW9a0ctKpkyhqVhWoixGT83VIx9THW/YABtyvSCFk3Ty0ddb6Oq
ffHZi0+JlpzhfJ4v8vcG1B5HSjdhSMQokG6bNETo6FQ3VvpMfOGi4BVif4SWf/XYOqOyBuB3sbdu
RajCsQbHm3T1fVfq7uB/OAibMw7lOLx9orGa8jLvL9Jcvu65Qxw1gG113HlFchctrdFrEi2xS1A7
3Lx7+0tmq4tjjxEKFHISM2WQQDFcHtWvKNX7S059ZnxEVaGlSzpDpsvNt4sRqCSRdqrDIMMt61D3
OycJUIMC4jiNrzn0I5LjzzVAS5NF90NkMdsfmqU88xfrMqZxQ7t+2VYbWQqI62MNVy7gnb0clI7t
Wg1h+pzOSfC66U0DS2czqc4+ks2bHvyCHxnWgY1OyNQGyeyFosl9BlpksW6Tmf4Ectxb+7nGzzKn
ovAEeiTNWMLG4BUM/q/mTSFEwbja0OybENAzAOkL/gd9ckzIZSLL7Ymxv+5qaJk2rs6k5iZsjoIJ
7rB8A61C9RdASpgfp1aePAx6JMX+6xSBY14E8kiyQKFwYCOe0vqE722HYNDAH3WmDiWbvVwCehV6
BpNTr7whON1+9V0fP39kDcX6M6KbxknRDpY6mEpKX2dXuoFzCvlCe8MrWI8/Q070HdIQ5BWUH6D9
eoAxXsEtzGc7o9hYsffBL2l/JnKXqz/WXJqfFIHHIBsCcaEVGH98gJGz1QsGXNr4PP+NiGwdijA/
YqixG4EOzVeXZ2oDlx4Iab35xp4akSueka7FiMy/qQkYNqOaDYxF3SF0sIeIB2d5rYkSvthFmFY0
nKqiuMs/Y7GLsciKjMYm29zDQBlrHg5IsTOXeeMKeI7aAdof4Lcy5xP1MWC8s6iuMdaUQnBpkZLQ
De4Qr3jqzn/FjZTYa+k6FYweimioJKhu884XOZJ1tzntb+AFzBoksiUCVTjnR9M+DpBOFW49WoDA
a5bcSV4Vx1MVjTxmtc/sbnkI72G3kvDZFz3okyj/Pmpr+jVBtsLfZDGTm8v723kRrHv9mJovItIS
hKDmrgqlFVvKmVaR+9bXrs5HMqYTYWSC6LDymMzB/dsWIw+G9KSHAG4+9Xkz06fItwlxWBz251c0
81qhJe80vKjfp3NX4nbmSsqliQDx6G50Ic8v/33hoogW9gotE7i9yRIyRPE6scG6IGW1BpCT9Qfc
mhA8qfwJpWw0njI06vnMyx0+TgX/UVNBAW/qMo4Z0Y8Q0lWORfb9ZA/Mfw5mEma6mOtFEbey3Wcb
GA/DMkBygBtKWVJUTLV1WV0nJPUisGLBdqwGpqPQye4IcSE79//0zLAGbKF78nmazUD8sGbFwyhy
xO6dj8z626AeAVOrwFZikFPqNy0sdHBJ8R2xRCiR1489sjiX9q1YTmO8bKPgHG+y4vQPpw5GEYTL
TTsfBfqClBw4a9Lf2s5+7LaMfzJieRXSFyMjkmTfRonBuW3zL2Hmwcz+oYVeOkQGcozjEzmcXSI0
Ps/WWhOJWAPuYNHyulaeFMoHwB9nfnMRwOadIUO68+KsSYk1lEg9b6bBDI2OdUsSCtySThCbQOXS
65bDYfC2FWcOfsZMJ+Gddv8y5kGkBYDHMzljAL+3QrFwPqO3Va1ZKXsApCM93ZV+xfb72QrnzPMa
klonwdmIyKOI8VKKVuUsAOgxEtf2Y0AH7RXngF39V6GY0CGoDNX/xjkw2rU8Ate29dDmuSsavZGk
VWrsXXSS4QsmLwUaTb/uU32JCY5B9ZxYvP49lmQUOp7+DRucWgQOPRq37ze7NzyNzCRW8ulWmLlP
dbnG4shgmc+W6ud0jO4IcTqhNI9coPVXQCfbrDFOKhUtMK+Tikb4Lu++9ByKmxfwXbGlwF2CTyn7
3+Laj67WLH8501brxz9ymUW89JfyuNL6beeN4hY1dtR0qD56c/eqWH065n27qsR8aF2LV5Lz9Z5s
k0QThk1s18/OoSv8ilzgNrVR6rZDregEHpJjNBzKpdf7wDy55Z3P2bvWHyqwBwqFuoxU62R1A3vH
/C7Wqo8d2L309R+E1KaW4KWKC0hcyDDjhVfVV6Bm968h47EKyNOKwHBZtcK6AUEOSbpuA57LATaW
xu3rOV2Ts9jYYtyAujGGWyRQBia8Cuclyya33uau7qXm9NmZDccluIPN7IcsKNnWsE0UHEyJvkou
TVIbMRi8ghOkSfkpjCbAEENmXt9GqL3vRmJvtmdCubWAm4VVKjb2jAxfeIOubLac9sU/ikFWlvB4
3M78800nEi0dxlokQVDW24yCTq/cVEyu86r22hCmiRJ4SI0ZSsPV8IgB0DSXcm1FVkyzfY4wSC9X
GhMoBGqNsR+FH5qjrLZbrmpipfKmmwnFHLGex49IWIz1mJozOGjx66TkVGCSS6Ne52D/nG3tR313
zxmgPT2yLZKBeHJexmZgfG9mxifL6WSIgQTL5hfgT4WLl6Ulri0Z0P6wFfhCZo2GNb9dfmT7UPaf
qqP5ZgwOVqZdedryy5wSm+XyMv4mIm9Jb6sUBjePdazr3q4YSH1cI1DuD6AF0hMK3aUvOMnBd1LO
P/x9ecYmR9H2itE9g1ODyxw2wPEnKe8pItROZM4dkQlo1F0CWJCBrj747qjWNqa8KUT2/w0EBEjf
vlPN+UkbDTwVrrHuNK9r1oaRJCP8oo+nzqQuY8e3YSIK8MWM4DTVksEhszlFyHhobd1Xjpk155m9
40/GMk3MRpVdK/zZO6lDuT6pr8NhVQZhjnBgnf3MbT5zjWnfXzrhyIuMaVDUP0rNcC+40XhHia8H
PpN9YipatHeYom/KpSUxR5/a1ITVfcfv5pQet3yfKT3Hk4pdW5tHD4s3fOyz5OX4vcbh30rR4LLE
Pr7lQbCPotXqM9dVZ1n6DcRAouKQIf2layE6PYy4+wzvOCPzbPesH0PDpqiHTkIOt31ty4FJQzQs
s77l5/EVfDMohCcUPPHKwE932CyNb/a3e0qN+RnyCToix2feaQQJdxGVRRHJQzRWpo3tBKLW/EX7
q+4reFQXov3oMuYKxwixF/LekFjHi1HNnQAasRXDxom0V5g0kh+J43i1MHcm312IjIsDxwSre15R
nzAQg01DKli7UiaDedTa/eQDvlgqN5XV/4WGC2N/M2jDcRRMbgVX8N8bT442Mlthruk3HCCMacry
TQUYKl22vhJZYxHJ2tL4o+jAlkvdIaqUz9aEIapXYE/zMbqT9Sa8qyxxd8UDWh16GvGwvwgvnKGH
j7Kzo3lol9aZk2fSczHjqQ3ik9d1cJ0X59g+R3tX9EtVleNjocDmDFmTCeG5sqV1c+CGSgDy0mlP
bT2m6F1kkfOTo2NL6rv6BNy0fx6shWGF9e3WYXgaya3sFFmR3xNX1L/zflG7BeOAlKUTAPbKlXsm
m6lxoxJUd2gdXFiHZvWGcKkyVhBdBuz3mWz71ljBhf2pyP0oxTgsH67US5Co3dmCAmVrOoSqOS3M
f2937aIwulHVnZelZ8vgosmKywIX6or2cOXmh6IH1vLIP6ImQY4AssQBRDF7B0r3P8sHvT6ad44h
6PrKzAIl1/f29ddIDmhAnmo=
`pragma protect end_protected
