`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
V82h/mp8FbHcv3//3zVZ5VW10Mue/LSt5dvjsUkiSGtG5WaH8H9Fv7j37k+xy+3/pQvfXcpqBF/k
iaz4/vETUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n4WSOWV3uUjyMD/l4IGcKD1bHONRRplCKgax9lu4YRYlORLHEpckVBvOD9geZHtnlLIjTLNUcuHS
rc4oO2K5x66eEf5+m+hNzaPYWCrVKWQI7/tyX0imMAsD4JQXzU2CP3ATsQoldRyYOQZmggmbIMiB
stLQ3uoRuVc4t0kXI7U=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zgo3FUzRcS1G0FRTCr4C/JBs44dp3dv5CUvkYU2vM2fDyGtu9ekJcjDXnFGi3Qx2X0BV1gEyWxsJ
xqQkFlu/f/1mutspkUjOMtKZNCgPGDHkGfwBEPN/xT22fOBwQJUR+Oj5KSeDWe2U4t5UJ4XXcGMb
ZV9syPFreDWYOTWkkl85cAKcf/WXC6oz+tOUowqV4nSLA1PaSrK4ohf8oaOGNVX+4Ji/w6ViTIJJ
OqmPJQ151npm7Kbt4RW80tp1OmABkNI+o6h4rwtTS1IHzM6bJ1Krrp0V+2aEmmqoZkuKINjX5Pw3
P4Vi6iUmJI0uMpdsCPr3MEC8HH4v95WCnjh0Qg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A45QQ9IEoKpoNXpmniz3AuFZmGAAZIhtA2hP4/pi+Iwurx8nPI4ZkKpYXPnn4DfH42bSsec35aiS
Ve+A8f1Q00bmFgtclspinRe4YgFesk40ftn1mzy6g6sLCNXhUm/IIjCSNk+ie6jVQS7STfOdio+z
cvSm8QQePoJjzlJz/jkNhsD110PhDAevJWb+C5fforY6kT0k7ZmJmE7btahod6wU3o7t2HM6+XGU
DDNZ5E+RLS+IiJYVCOwsdqQFDuRaWwS0k8Mk4UuDiVWtU0+QLFZ/8UGJhy2ZDSYlL/8TrrsWcD/1
Vku2N+fkWCj38RSMWEEe5TmUHSSzP7uBI6QwVQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b+wEsHDGMmVXUM545W/2toIjDItLsHFsIOyFDid8Fv6KhzBePVZlc9t2c1LfdAa6UEpdqcx5kgIr
+oVEglJG3R/fb6dRp2mvlu6+x0AYh7FK0My5t84q7uKZ6EPBxHnDds9FLGQdMDUFv8E10WtGrG31
lkto5q+L5WLAzYgiD3//MgdbP+aqLc/75XWIRhw/PfRn4OqyBU7xSBeoK9TDxBwOscUv0cQ+dauJ
dUQ0W2ZCXwF6cP5c47k76Ikfu69J0/IO+FTLKMkjAB7Wzsyqbpl6RMVdJ/iYscNROh1xxo2k+52w
4l9VnVKN7wTWZdW75B3V/MsNTrKb2I6dBdveDg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyn/owx08GdB/M0CwlYM5XwpK1DLRGgNdNGvCa53fvz5ftb1LM2R7yhWTTXlm8iqXlg1S70wvPmw
WVO2ZNZ0csmDdQcX4HNMiokrI2gpR08Dk8n3nzdOhqyFyh79/eVJzQItyKMQmJZNCvFfww0mtX5K
FbNe2x6ria5jEBEBp3U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J8WwILioFJtk4e6vNsFHYZhWTjvAMbsqHcnvhYKYzsY6fpaoYuWnjTNNNxS6JYZj7bKOFgPjdnBA
rKaGPLghV6UU9fx6UcBVLjNOj95AU3CZPEjWGC/GqjGRPxOkhGtDka91PZuOBRTBqJT8F+5qIgQR
vO7WJHaKezpaUm2zbeC7+ShM5p4Wm9L4dzJ1OuUGZNm39p9FbORAZNzAWa35wpfJ6PPOgATFMi7Z
sN0Hg00oxMFCKSg1bxvN3p4iC3rVT+wV6yuzOecq97B7Fu+tfvP+shqnUhodTpF0WYfGWHeK9ocM
Mg7nt62XJybi4Tm5rgYGMIIM0i67934etK5Aig==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AF8EDKLpUnsf5U27caIfzjHsL1dKCT4FvrlOxjBwD3ZJ9vsXwbWO+EJTOJOFymKnoSSFnuslr7C8
ZCAbkJJLJrLXJwfvC9hiPRksxuYzuxWrtwsjJd+5KWtue3gL5kHClD8Tbo/V+Dnr3gvKzMRNdFRz
i+4p8dC6/32xR0/NITJMYT1uOYu0oBFDHGLR02Wn4PqghcTR3gQMVeL0RsDhJibeNnf4Q0NsKqCF
7OscDpis6r9ZAFao+mdpLGI93rreTlZvJBUPh2RcpqOjL/8IUv0iM922KOCZ6j1LtvD0igXehvHa
5hOx0DDcMjOoejqJiwIqLij0FB13lDBsu+fjWw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16080)
`pragma protect data_block
BMP9G5RAk03qFRu5UmzfhEwWXVNssrcytF3IPfT2D1YwzbCCxP6+7+htF0MH/npmUrtgaolQ07up
AJvgfINSrtl4pXRFfkf8RTrA0VMQEie3q2THB5/DTuYICjNZeRiqDRdH+ddgVX3UdUwta5XHYfkp
SX0X0aeFTGVB2HJdYqh/2qbmZiVY9OjcL1flz89mmkIccHpy5Wv6JWn61wSduCtlM7V8wtsTf8/7
p+yzDkFWvmPwXFC4VDRYeomCGPFO0c4Ds5IQkTgSC1BF4MF8U1GN0t8E9x508I63TlP9gR3ysac/
ZoWxlrqPYK6JQ9JovbCQm5UiNShV2je5n3VfOK7JmlIOrYFuuJ7E2UYxP2nyOdn7sLnNDtTVD15B
5EaioTmw8w2R5QMjgSIgE1hRAXhE/NjCszb8JDOaIIznDzpELDaeNd9dW5lxlrbg9KONzKhqSLSc
vBIYT7qLPz2A4WOI/zHgh4cVnqoMG5wB3QHJMcasItPxVVUESnye5Rqg7TSARZusGa6+9x31jpH4
PGD8cHv704D8XLsTUcq5VjmVt5xLuOlbB1pyzIi0mHgSPGTQNczuiZFMTatkrqj49zvOYazPp5xO
FMcExg3Uk1jrlSPQ8qpSLDHAedDHFD5Q5oaliasgmgREOOmsshzPMJqaHuxFAeL9tDvzCt+FzqdF
peF3TEKOgDz1jsy2z7ys4YByyUCRjaQ6485C1K1HE02R9wzXIKFX0NpSuuoWvnywOxjA6thQmnp8
zExGOsetnTdlCl6xzGJX+ff8ob3jUsdFuh5iEejHWYi3wIhA2KZhhHWBYcdwlOiJ6eOY8qxpe1gL
KSQkWgNVz/2y7uqop0Ban3dlc9JjlWvNQumg6WGa/4xSE6ftLcDIrhCFVKq1xLcd5sE7AzxfN+mB
1Deo05scC8N+dwStXRUe+0OiZkxyiwXitTynD6hmulutKx9VerrQ3b/yrqqZZNO3zOua2aFftBW3
WKd1p/KMt/x0xIJrkab+9Aodk0iJyxo9j1OKvOhl9MPGZ6sQgm3K38YZd0x9QlUm6XD+kF0YcHZj
LLqwO/dzWH3KwUaR2/N4DiwNL06q9AHud3+73DJ8Z+V/dz54mXFr00HTUCE/rt1FIw8Olg2IVe4P
NZPkjjfAtrikOzm95LDjRWYCewK+CGnAGK5+9mKl7etuoOhNWz1L6YW3G02StkYVaX0fdIiNlwqj
E26j2Dn831B7nWKo94dZDNmW/ZY6hfhF0uPgdFi4VP3IP12CtWW4EK1Lt4eTY9Ps+LMrL5P977kP
p9y+avx5upPqdV2s4J5bJWmSF19kiHrTaIHRpfzyWe9ApgUeaFt6JFGYL+tFwQlL55OZgrqGxI9X
anNiF62eVLBnAs6EP6BZU81sBkwq973n+xIsbUseasXmYuLGZxgrBy91DGMwh5stbLkS7xDqa+HQ
bdUosbNipQvqbgsLzXsFtXVHBULglHZIPwB3W/wKaJYPbqwkxJeZ57oBKGDlkUim9U9/nOpd4+Gh
IH4bABLbQh3WyVBxYCciOrjuO0QBWFqxIVFfbn+X+/vkk2QKAHny+L5+Lp4tBJ8Djoe0bGwZpZ05
lyz/vUGnmKekhlfYZllvGLafshgqUymBp+gZjzvCjExFt0PtPlcf+SQ79QnnMxDenI1b1hsWfUqw
rah7ACYxQSj1Dc5ZfUYsPy7uZRyAWM2jbyZBmdvM/qw0AuZODxKfytlnADI5DbNG+ztXZqrEHADi
lxxHGujAGmJIrm32ntZSy3nY4LQCcZUR6AjVPMBWTxdq1Hkia0Qf5jQDK/jqu5qFz8DgRpPj/p6B
/see49Ws1HbpNmOWhY7J1gFGW1L2FIRVWqW37tcWBbr24NvPj5YumjlQF/uhgBeag73Lfc2nGr7f
D+MP6zgE8pmMqpNra9Ise+h3g/zxNrmIyQXmyNucsU0wysWsGtwG9pc9bX/qzZtLGUhOGdKN6M/f
pD8uzcLBi2EwLfYZ9u/vbwrfE96PjxdY1VHADNdd5jfZXhMsUQ+bstwo2U4tK4tgn/eV+KSLVb30
2RI3TwlUKv9W1m0H0c2uEXSj5roxUHtdBOCnN3KRNKDMsaTrZ3m6S44zz3c5a1Mo+FmaYpanKU9e
DEoXWfoOKsUnjIf6Il6/eqsllCGBH+LdlIcIVnyd8xLuQBvcdFKJ+taDi/l7A6Zcl/kVrJ573I8f
rxygsGNiMGI9Fn4leDQnkfPB7/x7542dmHHdCuXDlGV7F1rTpGkKicsSH9YKPzivBwBNV+V7S9zW
PE/dXlK/vwijUafHVeNl2be6e80GoiYrrY9avhEwPGry/5Q8TA9qaVn2zXT6IjdF2ctVAg4v9DTq
WxGp2kJH+ki6vZ81UNvxhdLkbYTZQUdO0IkaJDNJa1hEPnTusCDiqcou/KHsyXUTWoATJ6La6bg6
YiLYsM5yato2bVuF94Ee42CsK1lmuq4JQmw9wkfk//TlnuKJWR6bFyeBbaml49f6zfb6Dr8yNRVs
u+O1mn0yZ7LEfznLF9P5HlFwKETeCFv8KkYBGOmu6lcWDTXsAkeRfGdzjuf03jG1BlqjNgfKKrJi
ceyIiH/JXSaSNsJURIdq3ctBxaOfzjsr/gbUL87yE4/wPjAXj4T80aO7f6IWHpjqhjVawHQoZNM4
k/v3+FyPvRZfK5ntE61TOxKgjoPZ5LRMV+eAutaDvEPZLLwx0RYanHd5lxHJkY2EXaZPWD0Pz4qr
bDOkZvbAfD0VQJj/7Es/oirb/lPkLT8p+W0XgVlJcHEtSQVpDlidB0h4nOjYXDIH2Ozv863w3DFE
coxSenY+C5bJH0ulZv8EJ+xLyh82i3EcY+qr80kwH2TPVdwgJepKDT/Y7M/m7xbRZJH4XtjUmYJ4
ppp6Lg55KcEB4ImWBgyYGPBwlx60oa4txCq+6O2KyMJbAJ8dHZvTD7w++IvdTmFSTsqGp8iCcEsO
SDiTx0ZCMY+G05l1nX1e9ey/UB06bLutbLsiaTI+2KuOTX6eupbLGpMWI2R5Pf/Gk+2QtNGDPyr+
DpicPMLrtl7D6fvPSgDggBrQmfZArAVRSFFFgcq1+XBrS9SWC6K37dD3MVLGNJ7kgTpwXtxqcNkB
M18Dy0A3YSZZunJXrkKbnsNKIo3Yy27sunpDYg90OebzihcfIjwv9RmnmkYoKubUVhhVlQLrWaN1
0H91ckIixkvC5oIZ/3j91Ev5uyUIXZGSweXQM/KCQb9INn2wOznx98yB7mX98w5uZzEvjxAg1wOk
xKxr/t0nsOT6JP2zPx85HCUxg9fwfP9mfRaSSAo3kSGwujGCEdVFnxOPnk27I/i1I5/5FiWKtBrB
YMjd8uJKE+nC67cDOfW5BBHNidvbStyfxD+ogwfW2y4ykyYsnSIjUCLSQS5aPIpkgAzslaNFHyj6
oxN6jMrM3ZBKKGDikA9JsO09b3jtcRnlDPZIvHdAwrgAYop17SVYIKERHjowdGk7fw7TA58qb6wK
6dEF5AW8UuQlk0RcMYdXSOor8jZaWk82aiUeQ/s/v20tirc+XTjo86z1UZ8ynZhmfgHgjWmYNoPv
+8vY79rxOpfWisyU1OuGrpfx5z27i313l3IeqBpZ+hioY8A56JRIf5frCCtwiTgVBONnMu1cowrs
f8dfWIzFFsg/FHwDzbM5WO9nH8maMo/IXzU51xZH4kYskczaLZzJmHbsoPTxNzMxIScGbkhTEuEx
kNP1DEw8PAHhckJp8Sf1moIG6EqKVu/iqvgCwB+/ynxDp9I7w9lM5xB819a1AYasOTbidj+KYbQm
967mygxX0F1NCkrBIZxNaCXsWX48XKKMCbOaY8xYvT5+N/E26ijiPnX1HNJ4x0togI+6IXNxwRWo
Kcg5+AeF4ejIFiT2kSWT0E3rSXJ/NMhdZT/CkdnfHGkL1ekXwgcleR5psepIE2+1evWwOVDrW+Pl
Zi3FKy7dIoWVHOsnzTc0RDKiftSQV0Z+b3AYOl5dRmRQkDd7z30jFzv7+KV+OaQagZgjSX/CqUta
NJk/wUjNwvd1VBhqoAgu7QStNVJfJNE71A2m02cNcir6yoo+IvLrmh+CI7F9ir7U7C7UsvhBjRjD
RELE8wECuC81yPzDiwGnh+d4TaiWjVtN27zsIe7+N/VNY+VMIydgMXZ/xZehWCfQI8pb88AUpmMY
YvYZGlxaWV60CMI0detTKF/V8Ml/XYlupbfTR3a5MLCrvT8yfbuLeo/Y7qBrhDZ1q1PNZPAqaU5v
coKibsXCX0hQKKJBUyAvCvFM126Gn6uiKY0NdMDsCnYrfF7XXUT82WxVYcYIPHilYUsvor9hcQS4
qOZ4YPTvXvykEIoTd9grd+wNXaWLBph+9IAuObOmG58EkCecNhckXcH7KWkHmvLQkuWAbQjID/9G
hSHgbVrQazdJjiNVxwuo2zOR/fVlbxajwrOgaoCwXOKTsNIGcSS/TtO6jpZD4iv2DDN1a9rb75Gw
shx9BFrF/MT/KHI4uBg8jbfFxvRB5sjH6uOJ0gk+aUHQJloJqdX+3HtBTV12BiYLWOt6bx+27kwR
UFtMtOSsIU0Oiu8ym4DwUjcE1nRBGSvBNRT/sRVOdsun5mEpzXfM7Lkn3ScXBdlUKatOQoLrOJ9B
h7/G4rBdDI2/6Jjvt22Nzb4tVLU2n4b4vTXCKnJAm8OgQjSDxFCT8LgWv3l7o7arnOK0Uou9vQX+
5zaet/TJgSVdl/pbYk+IjdtoD2N2jwZMOd+k0C09GA3aCoeSzdWKNmjsbXX2FTU6P8eRfgvrpNfO
AYubMb1Tn5StmXnh1L+WqVMeT8xNeXly5p6I+gcF9FYbG1JKS0IUHrZQCxz9WXC9GfodvUEE5TW9
CMGUjpdzNOCkyYrEuKYJJ/BWjUoLAY7vpVbMFfv2D1XXcXm4vc8KJYHJrMaUwJnQkwJRfvmgVd/Y
WngJYorGcwMf36Fhf424m7sJA0LbqkIZFPFdR6KCna/DyofvoAobGVb8r0ICFCkS6JL8+sBdbHBN
KBEl0arWchNEHUHIp2DGk+0yagshBw0N9ETbsAgSpN8dfjHtMEEnVfkWqPB95rI/NprWz+iLIOga
V1yxzrOUbCYh+m3mvAPYV/t9lTGqanaNyPWOZIGD+eYVVgazUf3RvRSCqBR96Den4qGHvx9/Whfe
nYjpbCNvUW0yRH6e6qosWPScjTv3P06RXQC5YjiL7M8frFWnU5Ghw/q0hGDvlMnDvAAct6KMcyqd
GAXb8Y0VzgRR9ee1Sz4aoW5BWRHA52O69BULgJlbqOwUmf6oDCExvcNe9VHSAEGyGLjrBR9Gf02o
knpSj/sOE1+CAe8D4vQRx2QalHNGYqlSKsdgrXatqhTSV++j/dlCwlhVEKQC5Vh8cy4AJZiJE1eq
IoBPRWtJWxRxeKG0WJZdfci0x1XIZYKTK7q7k9c2WZnCwSZv9XXBWf6EjUxkSSwWzGwbN1QjRp1n
V2kHl9tF0XaeNZOVEcDTCaOJ5z8po0fdwLRr8FtIxC1rup4lgyrV34c+HdEaVEQl1Hk2WXnZeOt1
SGAXLwvu33y/w1Up6zzpiiqpFYnIbvyso5dKhrUtXMCyOOJhZgdaCKKWNM3Yz7upz1FzNB75EnPm
H/D1469OgwgBmFdjh5BRU42TLJvaMY/2I74jwc6TLIJ0DDMKkk/fgTSYfODsCkGu69VR4YGcU/VZ
05CNEnXO/dG/vfAJVk8qsAfCMVTd+4qN2KmaCFxxuIIma2/nwbSFdj0PYkiUrXJ2m+zwnPQomow8
SBLQtI4UXyDaZKZ02QguluUoPNX/kgkxUKomaRy1ZP+GTa+x5KGyo9B7dmgYh6kGBIhXGBHU+mnT
zkZtrZy8OxnYPz9xMvr25T7gEXpkC31deCdJ7PL4VFX9NEreNKRQtTaaWj4wmTODL1Aq9asOpFN+
fqYtnkp99zovATUTwHlUKyJfSCl/3BQy+qpAa6123bTqHgLGeN7Adcn0r5WIoiMSny6O3PfXUhOr
FaShYiTzkMoo7eP3lrXcb72mZgytPa2ru0V4LcThRtt8HqG3KxA6MIDcXxhQB3lNzw2Qk9814kxM
ml5MZDAv/lIETaphEDhs26rum6WSkzV5dBFruwIa1a1QHcQaAXRordKudaNckMPgsYN0IVtE/VXX
5PlffDxU/CnYddjGY87UlrXtYkqKSA6aBcfiPHrUT2B3WNuQhyC2+H4VB0lxX6/9y8CwEZylDePy
hK04ibcX0ppEs2wAuf6jvyQkUKBhhhiXaYwZygf27aFdBWItjo9ZYdsCLxN/CSygBw6nh17L/S9r
1bQ4mPuLs/tt714KevEjLl1w1/EEfEAfbKYsCU0GewR1Rt0SIQla3VW+qPeV1kI8YqALCyY6X2p8
r8z+oXVTyCjukvFfHK7ID8lRUrm1e+Q0MCWBZ5ixPqROpywXzh563A8TZKMhkkdgrf8UZI+R5517
gnhExOWTvM6e2ckvpKrzvVSsbZQvcdeok6W1OKA920Gkqbk3tqWOuC/TrL1yPjx4OiADE8ppNhA9
2FmZ7FKYej4AsP7utn+7ZudnB9IhBuepV+4NriwpvZdypm2rpo9dIE4W3u3MMaxrVrRP3ZWpQR0c
k3KFTIQFJxzU4xpu6oqdZNnD2/PTNGHXuL+W7mjLAKQOCqzU+b3mAlcL1xxJTPnCVl2a0DRHWy1S
XaWI98JIpIKk9ZYZz/udszwzuOnB70IHOV9qQ9eMoo24EENhzcDfTHL9zFUGziXErjBp+bkcig9D
uIF/gG2CW0rvB7LNKu9+MuSuDHdMaeqzF7khko053TIjQaTctTTNCnEiqtxH0QRuTW6ez3MBsPNj
uTkU9g6T5xMRD+NvuMSYWheY2qzP06Rk1Lv32Gn9sG+PXP36/L2NTA3eKdhAbvE8Zl3mdbhtk3ol
hmglPgNvPso1rqB8LAYKHglr+IlOAJMmh/R2EreAlYm2UmwvsWWlFSDeClEV0HPHkOLECYkCVhyB
iZbUQf3Fjlas3MgYGQRFv6i6LLLu3/HphVRlvI5O/0gRs7XsZOdXqI7/QSneVFKQZsQyZFW/g3zD
ugShbjkiNCFNY/gmBGgRcn0jy9KoG8vfKFeisnbJlwDwt5dCe1Ot0JdOFaySOWlsdBWpcAtvusDA
KuUI4VjF25Ky/noSfNLQ6PIcawj3H483aSsLP6MyFQQJMu5xH/dW/TpsTKawr7payahE2zcUiAnF
tx2E8kehGWILNdCmR+XSYHiDWT73qLMJCrt6QIyagy1NSWyeoD+qhdftHTOc9zqRt2vfOLAI0iuP
z/Tqi+5j9fqFi7eYvC1QVOIQ+ioyf+xClqo5CLty9Vp2n8Ja/NaZUascDrJ8bn98gEI+v6buCooE
EoeO9qcPBKDKn5moXJfXyr/TWN9S8MjhrVnPRO529f7xRnArFqa/0oYGvSkeGSBiWji6ekKn+7cJ
4XAPtvqaFZDCFHpFX4kvwYa5zN8p4uHihOcNpHWU2Fm+6jK0a5DGFhu1x7KsHXhMYAW2UPgNzCL6
zh9+g9W5qS6hxUCNWU98BxnDglsXL5gYhtcXVQWc/T2kfznDog4ip1hD78qYHQ9O1WV+xg/g2ORu
F/oJyGnPo85yOPvAWbmIXE8NNr+UdPtpAGkQ5W1kLuskrAo66NfVCQ9lx+D9yb0IR5VFnO0ekRFV
RtPcvEQSp7e48J0eA9f0r1L3xh49O80M6G8KW1SPdtgQTlHEQ21sZBC7xnikTF74UiJTXfKiJwZo
Bs+2c9tDzEk8f3WJNdZvOP/faTkWgA/P7CVN5xgWca8lYBAQNWTvQYIlF2yBseK3Rw+FWtBvhsO0
qZPiqZ0rnbQHRmJBDGDIavT8s9Bwe7f4+iEAqZddixOJqIqmKrVrhtjA6NX/vhsaDzbvh46Nyz1L
N8yUW3CBR1yWPLh7Zz8PLs9CEFvunVKDA90n6SjOjmBxewB9BBa3tGvSJz8k5blgt0WxXuCBYAVu
wNo/GWvI2g1jSfYHAqNrRAqIaN3DlvnBSoVd/8eWM7xMwIgciVQXdOXZNRxxvDd8TbdVF3FBfCOq
/Symec7JKHgPycQgrZT4lcTLeAPdkLzi9aC7ybJsDTdI53Sc+C8h34mqwEEzzdeX4OYGOr1SIAx2
dgbE4/IzUsNGgCOukLk3XJSSUrHzkTBna1YxQJk8nFHZOpx6/8UrmhhbJhfNjfp6BRyDYp5YVqWf
kzqvqgfpE+YpQ6QCTDsxOnt40fSFm2s7CUWziOyQb5iWa9QACOo6o7dl5sk+dptzHYsdKtmxXIVZ
aMJfwMJ51K3r8RhvvoELbTDpnFrpeBqGai+yeLFjf02Z0rY7FnYIx8RbkFCra/kbEE9+eI9+E+Fy
o0DmRRD9246GMQOqO7WNdYyP1+YxnQ5XYPXF+hOhJNkXDI10CLE2fn/cXQTBBpNjIgv0GVGkXAwC
RAXKe7wyt4WDa8rzKFqlSAz6IU+NG/EDL+sM30VigpzbP3NfGow7JsYMr0stN581Gib9UDdo5It7
HH7+1t6EHw5lE4iqPz4Uwfub/HNXHPzEp7juZf9bly9KMVaVX/ULjmBTMRFXoF+KNN82iaA+i37W
G2VEifk7CPbCaBzJg6ILCqpwfhN9uE/EEHJ1uyvY2n3SEMkzIUC8tnCqtJwcbYRLfw+WAbKG9Lui
hfJo9bpolH2gOsvEXbzAN6fhkeXeq2tsdnlmg+Uju1Hzda+2GFt/sSEDF56YHWRqFMqQo9Mv26k4
VxPZ9K7dCANCM+CdGpcoT0w88CCdf62k0ExfrpU38ARVWOYKBEVyVUjVNgkbsEsk8nvizGp37CLQ
oMmIyUQG6iWNkl7gATeJOcoTB4LXGSaxk9qvXbOxOUY/Rk8cmbObhW6EPTHWF6BnGR+5+HJY2os1
7uiZ8ddMNVoJRBfad0CqE2v83tQeHsOjQrDBOhWaQ8KwQXejU+XsQ0ZzhWZKVk+p/PB1HiIshbWu
3mzey+eQbVEkPz1RFZJVMaSzg/L6RMXEOdW9HQR9lqtr5ord5JMnLyir7McMmKP52jAAndhzItBn
lUabTy+lLHxEyrWY4gOfGWDgIJ+mh7mIrXzsUvTW0nRIRvLdJcW11EVLWnpXRE6vw4MyAJOYwGJo
0izunA7rqKQjRNbzZJBg6FpcbqU/29379SG34LmcS2K2h70+VyXwLGSboV0P6+wUAVoWYeklpsAY
u+fWjlRA7LaxjFTo2l5p47dgGxtEYTtyAPEbeSf2Gqfpj3msHIhgkk5MucHx/JyIbp8usOm1Y8Oz
k5Ax0A+wObwE7KZ4EDo/ziQuDRwg6WV43rjP5Kkwh+K88aN2+3RcV6VonG48nuNtR7VmIMEp+DyK
n5oUwvf0zNcAbgMQTY4pRAAGXsVV7kTflPKqQ9gulEBbIqWDZFH3Bhh2dQDOUJxeYT0Qj4ySYi8h
hwnIAP3yboGqGC6Km1XhpdKhK8whUibUym0PGEIQ5hzY1kOd41KJRs/W5f2bE8jfFXaPRRCYHfPD
m/BkccIBzjGPPFA0MzRgsaq6zcgn4UYPDnnSVM5Nhewn3FU73W2rD6DCx2IpIhqPxZib2GzG9DD5
OSQYCUIt8LphazISHXIFmaCXVyhepqpBS7HDG8JHdXQJA/j/Hcr3JvR+iktggZLGev6U28bzo1hV
aabi+JkEYgXTbocn4RulkPYVbgJu2ZH6jNfpTCGcr86psym/x9+9XxKOfm+U+30of9Ny1zLZzstd
Bw8ttiJEXWDbyau0qD1F/D23rW/NezZJeOdKzLm4WnbaifVIt53iXduKV6Eul6mtWQTgduFr4biX
3M45DqIGyRLJuILagQP7T40bjpWifKao4OrgtIPHcyjXgGOi2msCNsih9qMqT6wZGfg2zt3fcjVU
1JOTvm+5J1hgPqh09DQITsUUs7HV+o0cH9tm6hPNh849c02Sitzelp9VjLgEZJhbFxBInJ/+AYuO
VSzxbsc00apYs6pqEHgnvOFXUlwq15m92ec10sIUy5+ycDMmTCxbkzSKibJPsbN16T+tFcM6f8MG
Ay0uWTcNwKEvz7UalPfbOI34reGU9AhVLFDQexi0pTbhiLF3puOzgIhpKgt/U5BpD4aiFTFobHXG
KxXGxdlKrfzNHvLB4tqIRZHTkBPGqncgbs4NG6gLOb9k5K1vOsJE4/B/1ZOhc0HJnH0Rt8cSpm1s
IidRxolM6hK0DFAJaYyw5uf7j1o7PNODLY53iblstRJ/2P1GUNCEGcIqFkgoR2MjqW1Pj8WRXbrd
/vcjortvGpIW6VGPXkv6OkEQ7TTdey1AGvHmNYFH0bipaUcgMcrJuh25yJtp6XEWnJ71klM7/GoB
s2+a4efeZtMAX5y+4YJcHAYxqacJWETgeTtiorzkSleIdiyFT8+83C5LYkRdiqxvyC8bGKkzc/+Q
Ow1tJChPDGXeIxguHLi0lKEg7e8H1Uv9OAuew9hF3VvbJ7AwfhxoqrILi7Ut3kzL81QUPcu5JGJR
t6p49hWlW11WWzDOqskjKtNkaTPCuhzL6z0uPpqpugZOza1JT6uptjCtlgfoHmk9/i9/yUa6vpp5
qh8YrZPt2gkE6W2lnGxtVOoAwjjuMXpk+sEt7evxyuKKtTxCY6TnXTbgzEm3rWvpReZYZQoGgmn1
Nhule6/EGm+UE/pX6BqIAWE0F22iQNhg9LLhGNp9aVR3iKlj5ny2r2xKvYLjio/QPuii7Z0yO1o4
TgLbZhJM1bC8RSKV8GPy/J166lfddNy9m9zwE/7XlrFqjP8wZ2yl7+EESqKtEUmy9OW3OFkYSnRF
gs8/DgfMtMEVPryTXuOXfKF5TA4IzsymZ8LvskBxREZKeQ3Elfi8aBlPI6pE6ThF5d8I2jfhE+F8
ZJWVToMxoHzFngwF22xwuweRH3Hyf396cRDv7oSqsL/Kv7nubTkIpGqWCpVlvMlUATcJlLXoGbqJ
dp/HUGqienntPsw0aMZIuMDcj87qCbCsKr+ulHqrXd+tPTo4Cfa4M5S8QcO2UPkZ17lRcifFzbWR
D2gnj82pXS0G3c9AGUG+GwWFx67h8XfV5snQFcXAxbhQBWYJAqEBi3fedCjKmlXlxCpIqTgTgUgc
QGVGwm7MKIfkZQ/5jfuEaLPrc/GoCPsG+fd3QhAx1aKkGX0Sdt5Bf15YKlKLimdQdLIlh0R6sLp3
yZUls5A9uaBDZYZBveYUv54kmqR4WFx03lnPh99cg18E2mxAd1ZXD6DaFymVvWHxtl+JVoMBno+o
qmIfEYjrrY7RMezMB9mnbr1zAcrNgchb62jXdgvrTgIwUMyp8q93+WS4k3DVdr16GQ/SMLoucDvV
LzQQNP2eGraCsYCjR4sgqdCF1F898FV2sIB7RAl2qLstZbqgkZLW8n/4W+MpaZFTXwvx5G9NdJAR
ZjyKZhTeKI07fLQ6NOdPO3o2LthfXXRQcDBOB9n557tdF2MqQNqCNkr3U6WgPgtdJFdAscOFCdfl
MA6aV0wa+7hmhA7WhxhZ1BVKTLSLVl+30d0rixylfeTW24IwxzSQPNHXBK2bsoglvHyR3HzfxiCp
TjrdSEsiLcG8waEVL16NsUHhJh4ZF0/97EkB+SvLhbpfjl2gvm7SJbf6sBrgeaW9t4/FGprwzpE1
FgAKY2GZlPZi5mR+EKbCA/FWtyUCRLYYgIrtwKK2AMQEuoj9SN1/ckmBIvpAzXtUWNEs5ppiXC3l
RhMAVde3Mdw+Sey+nPKrOvJuE1T4Urf+fpzbgefuScZGmZMNvPlWV2SjbnJ2DhDf/QTiL4qxgarT
hTpg8CFBETcPV+jthNWMUJVTV45FpNVmvkIT/3G3RtxDuPD//UbcHWPJJ213r+HCqQovQKbGEnvU
bndkqkuKgAUGprkc4lE2phsjTOBX2ZRPwmqmmqGquGhP/vaENeVjJn7wGzDCbM4k/HZKTPZOjqvo
iVrEVIGkVFI2WoeOYuFwlDiGEFI+dkqje/Q2GXPgJnCs/9b1814183l6/j64xCF2jYlRib6t1sqA
eVXV7DcE38dItSN8WCdA0adjKeQ1g0SUQwUi1vI/7dB6vcz36HIpP/9wC5A8qEbU3NK/h025JIYr
TYuIy3lbR/XAO/d2UdBl4KVqzZsTPSeVwczObEuGdfWlKEpH2/ROOijkISS2ShPFOm+RA6sMSWlB
fMiEN0sUFkeVG/+7dwCUP6VEOOCy8uWQ5oJk8q+dpq5hyvHFDtnKDRaJ5S0ERXDxCtJGWVhUsv//
ZEbFMj0JnK7RIgK5xZ0FN2rt8n5oQa91qjcMvK7HbfYuLpc5HUSOLx+mn6VV0t8Wn1f1XoJHwJ1y
AgB9BenEUtr+S/UhhSFOzKZAJXmEubOVuiKFwCmnL/h6tiTdC1BOZpyzak9+WowR6qWYpDL3PduM
9RnIt1lYIC9pHu2nFJ8OIO2iq7apDIYmDXJuuLx/Ho44PYKWiteYfjZ8VtxK1rxGAgc++xPLytBd
N7qZ+3MGD55EV2DLu/WdjVssM/RN85rpwdbuw9C+sjrPeKTgtGL5Ccp5GrlbpmdwPWHNqbsEmBnr
+cDsSPv5vm6KUJUXVgaPL0SluM/UWuxch6Nkq/lxi/XdkpTvYG25XrKn1VhognvvN1lymgjmGwoQ
nn98srv5cBcZo6Cun4T8jbWicl8xwtD7GxzMyAysHvTNcaPNv1L5rEvV/YD/Fzh5ZrHdwOOC+M7g
9uW80+q0wkuGLsF1sGxL5A9A3EM4vGo3RCQN6ewKCJI1d+vDgBfvNZDv2tynz7yVNfcYWfOYPRhq
3Z8flYB8mEn5lMt6nh5RK//hvBHMX7OU+nEQ4qrds1nP53nOR8GEjrJVMHXH/XBvcTrz3cIzuYzB
+kCHYjDrL/Vq1oovpua6rj6Io+qSbJVv6o+kSGwaTv4naKpjU4SVaLRmpRUPp/4GhG3ill0YKPIz
0P6VQN5B/Ax8kMEKkqP3gAS/jM349FDb2JMPIJcJkwuWVrKA0h/zwl8Iz/PWMMNs7fhe+GJqYoCs
3bZ9qcXcS41kQs+2kRj5FsLItONn2TKOc60Bk9L7Qt7QH30n3lXd9Iv88XGEk7ObXCEEvH4UeZfS
/Lqy0GbQ5E+G2AYCTQuQYrhz3PrEam7JzmInIGhWAQzxHNUbwl8Vlz2XQB5ko+MJN8LchuWVQoqK
BngDRG8WIus6vzlB54qCFMiHZC1e4fx8xL/E94bm95D6f53DIpLAC55p9SfcbWH6OTZuVDmpDb6N
7mXUbtzsRtdGl/zTlyiOMmEq9CbckBE0ZvFxmFz7QKtvF5RYc1Q6ny3vP7WGV5pw8igtwE0erdeF
VsFE+OHO1fRFIyAx4XioC6XYqX2bHzy+JH2M2hxrIaD/NC2V5YyHQHgLmnFfVLBY+2/cYWCXtyl9
qyKBi8ckLIf9Ja7RQzqr+oNAqVrSFmm1Fd55h3MpV9dNfhnflxTbkZ9IsRK3+2ixS5Ist7wFP2Bf
2eKRuT12e5sh38QCBJjnU6iBF1ExFjpaqokcU3Bm5B553KVDhkx9wlqx2LffQ/pl544UQ/FzHM0I
p33nrruwSzhiTRNVG1/OWu+mghdSU5ifhmv6TjwEeQ9mrP+GRaEpKRv3HhlD6vgZX5iR3KT/vDMB
Gyn3N/k8yE+P+qF3rtRpAUERh4DUGzJEQJXFPe1DPFuEihCfmuvuzhuUm9aAKn8gw9SB8BUv5ZPU
BVevzvu00Ou2j+Mzj6Bt4PWhy6SsxuLZbBIGUOAaedbG0ZIZncE4/EvOvZq+a88noD0BapiYz1Go
XGPHt950NinvkJs6Q+5QTHdYepUUS7Ni+UVrLVKQqyTLNcZwhjCYh3/jlU1aLm+OCCl6hO05/sZi
EjK2sVp+XRbqaBqJCVrt1yLdEBSqGnL3tepNcRhz8cETSJ9qFqr8TUtob6Ehm9fefrVTRywqmB6i
FVEiC/HLFY6tW66MIcYyX0jurPKAG20pgpU1D2rOb38ATQDQP6WO4UdO+/eJ7AFkyabMZI4/QFdq
NC5/q98W70DZjYPA2zWfZ1C8i3QVFwHMSvWa5QSUlaK8FpFYGIVUIxNohw9URbbR26SCEB/TrNFa
ngT/nCoHkGvR1EncR+CJSFQYV5YSYjv/bZ2q8mlFBH+SLw6MtjKsl7+NkMqkFj4rCeUBoujtRrM4
NREiG2HznKxf0jPbX+OjH2bJ5rihJZFWZNRRjEBnySWWzALAGFV1b3DjwMorB9CBgz11tuXul1/2
BLf72uWPJlCy6UaVeQR6PXLe4kr113xSBO3hLejhEVsYkcK2A0qrTpprdMW0id1GW7JE8thK6S0b
o/M4ZGnOmFF1LzKh/G7ktss/KaduDy7ng4oeyv/N6IuhQtx6S8v02E26WMRcUQ/9JUHRrBAOfqT4
+Sj3B1rp+MoLEc91/jPMyKRymrnc3pRTcsmV9ngU0nylU7+s0AhIR7QNmMuz1bdUQW94VTjXP6YB
TwsHLSOZB8e2abgqWBjOR01clQeWcVFZOVhtkBu64ZXVXSBSPiBDURPvKmRs+2QYRMH+KecAuE92
7LD3lZqMMT5tnQ9EOFOvYxN+SyzCxlbSrIkS7NatMp77y0GFQV5+V7XqPYSnJLTpRI2b6xBPPyB5
Rpx7YeYA06QM5aPz4VKLLl5ptpaDC8X+ZARN30LrmCnemq6dp8+NaEeJcEt8zAEk3M0thCzrw6eR
J674QbH0SxVfUh3k3jNVBHXJoVK1ZNmx81+4qaHEoaR3L3Nqhxsct/ad4Gb55iyycBaTeoce6Rnj
EWDoUSYaMrxBEtcBp4dqACoLF1ASTiv2Q7bremViBDP7WEqVOUyh0rciv/+YnQFX73hTLRI7ssoq
+HY+RDmUhADVopeLbOE4OArgiReLjng49DHEY4LCO+yOIIAu2EVquAF0kcixRSs0AiYTxuKdmiVj
9C5fzRX0na/rw0L1D6B2CFUenq4ZKDh0y8uyeak9908/fQsHRp/ch3PpNLaBFG8yfs7PCQXB6FBO
TgnOn1RVtswet78cZe7noUYzAClA/AqDuPgfgwSlBQ1rQNWzSFF+2Qxjrcp+J8l3k4Xi9n7lH4NK
OexsdMaTv0fqM6jGH2VkoWRvsDBQmsmGJ2+hoHo8Mi1BaAa/pp1QFsl5YM4koQe6tKuoLvMWTuQf
4XqTlx7ZnzfTuIOx2eRM64ejKsCPpWydKTwM4d1mSntueVApF883yahhJA1D18bu34u4Mx2OWTcD
4LCyuE/XnQ5ctOutvtitdMm54aivFIJbXds/8HmBcHpYGtsxB2fxk9uN27050y+ZhQWTakHIBDEU
zboruWW1fv1B69hWqzXovCJkdVaEPSA6j60s6f8ZC06ae4OLBhha+fTDA2XU9D8DzHT90iAr08Rz
fokLOAVVQFu8j/qn35mRlS6Js2ACsZJ0UDDgokhKmL+WpOPh4f+tWX0CWwMb1oUdrx1jGZ+tmhFQ
xygfAv31NlqIWNWIEv+vj9AvWyZIIRSaYUkUwr7CjQDV0SaBjDIVJX1yExoj2OEBWY3JSN0obE7m
1Z0SeFikyYDWLZ2GAd27tJSVQ4Zh48us/DGfKjcDIaozFZ5/7FwDfwBcVCXp123YHhd8SkRzuzSc
JT0V5bF4roJEJtJreAiVddgGifwfddaFNJM0J3u3i+F1P8LLLG046e7WnfyDaUIZR+YKUaAXqsiK
YARii8B9eOqovs57PxFZaJuAOWNt+TBEaKfiUknFW3M3GpZUHDPShNTZZ2QCys7cd8+zZFmCBmgo
FMg28s+a7A7r/j+8qo429XsiRnZKH1r/3jE6FLwh/wrbPkvDlqlsJ32+rdbv0MARTeFSX1QvoFN3
vPpP/VlxDpgTcPjEQ/CNVczx9a5hTiNKQ7fffhTlrdXbXFMBWUy578afqZhKUlwI7JF8anVJRO5D
pOSVtmLueh+WAHIetAM9qf8g5oFIkk4bmWnidMBtXZkr+jTFI7bROWIxicMPJJzPAMWL+/gy/EeF
TK7QlchYYMEykcIIv3CEhoG2L4nszO+I76TMyUgGtXkjwq7pu6ab6MRw1oi7ZJAnqiOf0PNkIwuR
p+slfr/Fuu8j5pOC5LUAUcEL786RbyvRAAMU3hu3jo7dccwWl95AIIEojAqDUfgrEd/7bxU2EcaO
SZ/l4Ty+Xg2EkjqYEK4jH+lv/ShzsBRWeqNB2+LAONDFGZNlLrJY7YjhYit2h7MexjganvpDRp0w
1FF6om4igy9KPlCC8guT4YwCLi1ktcqHvqtWKK6AhW4AoBXz+dkLYc1FJE+45UHdfWZWFSeiWVEW
2qClk5EFLNnH6dAbPy9xTAh0IcE1fySl4BxzhS0wdICRuKYeWyvPpj9URFsQ9dhLXA/py7QHYMC2
SyaWKFPCSTlXi0qHTsY9oYar8E1qExEmTATTmg3fE8Fne+fP/bZ90Q8AhCqV3qX/xu8K7SAy3SVP
hRt/puIpU1tNLWMykRnyE4/+6jSB2/MOtyfUEvOQFBmke/rHPv1JnQpnzAtZ3iS1rHuLXulyViio
bYEzd497q8J1kIlgWqWp4cZWxNZWaJHo6sge5h0FKfHDE56LqySWJnKC7bVu5sXPtc/eOcJkFAxC
qXislbCxs7y4ev+/GrN4LpWbpQ9zB69LwV2p7+3LFW6BRp2MGZ3Iqlf2iVdH/AZviTqIKQciqPOa
Ht7pf6FNZEGMEuyMs+jXDXP1U8WokNUviJ4c+uLVTQO3UpiZVdavHrOm0oDXxhzEtd/reNNZteJ1
/rk61C33uR4bLZ38bfghn3+I9SjquMMBvlUat/NQhewIXnvNJvnvqmshWL//JPlEdZw80mdLGimw
OzkEaSvppvosexqHebJZvFXOC7aopx7PzXPYbMUqIf0hlvQWZ279PPYUlvCjWa4QBQy/Qtaj2ll2
au4ij8iWgpu9MCbRxVLLzXK0xDnP/ptI5DvX7+iv94Lti8r87f+BrZFWcAnzxROpb1V6mIRFPmrI
vdc3L716Vg5cQgFfwGk01ZrTF+ozJrmTkzig9SqoSk+RHjEhiNDvSCYHML/tYy9GtcAjLRERQ8To
FQYdXem1H/rZOCjJ3dAP+HF75OLyDr/NCKWv4Im9mOhubPaSoIIw7l5X115oCXF517f8tBDbUQTm
kztPGZQ0PrrelsLwevusb5K5UlHoBMOXnTZuPlcqgSAjfFdEbTIqglsXDWjPxTEIurszzW3ijuCW
ytqEeCgT7gX+LgWdoW31FtPcdyNYVZoeCvBBnf/AWgyi2FD8AMbYPLTmjYihPdLL7mLTm/F3Teow
1PChSTDYWkm2HQnZ6/f6N+uVZ7o8ENJRKqySUabdx96TXUOm5bC+Xg/TuUi1wnx/kxmSrLShOMqr
mMY9Sg8Ncb9xmoyrXmkKaHFLlWTfZisT51Wgp/Yif2E3D2kO4rbyWn3Bn/n8hd6ETBm5vHhDU7QB
MPUced9TrdHGtvs7lJ7ED2VJTXQ7DJmIV/MAeDM2/znyBiQEd+bx68MIXZqwYBsx5yod+49C2gN+
OKiuYcqgB1lTo5/YCOj7zXWR5T77ek4I68AA71CaBxWmue4VYBLidbFHeVpgJQ+HbFzeJsUpT6B5
DN/diOHcaBSBEFQv8bPLv5maSzKs4aw+AEoAup+mwz2YXyscGvS4uiAmKU2SC5TiT76sMuUo1lpe
DPkytAKC03ZeU8D6kgO6U+Gtn2RQT6t1CnnzD0AweM5CHlwGoNS86rJPgb4ZsEkso4VsG21A6WFp
aFTB/QnvIsJWXniI/pT5cXpHz4A2r/DFZCo39jOGn9EL5W4vkBAipjhpa8b7L0ww50HBnovBeEap
3uCP46Fp1Qa4Ul4NircNSaU46boxnQP8HALmjmGS40lVY0mrNL9pcRc/T7ehQwTXb13F5A+1e9/M
7OD0SOgCeFE2S8SeB9HQE+dBi6/beXjPTna3U4sWeG0D0NJ2XwyORilgpQzjrow9GT1muT+ghPTV
VF5lp9g6f8YhSSAbKWXMyjytXoPr38cxmer75zRB4WibN7q25V2GNzwUDSuXgUr0XTgxDqFjlsLV
3E8ll00R3F2blkgJGz8KaRbX7PKY4469memNChkm6LGnGdEhYy7hEv0fdkUHZFMRkX5hi/KMYZ4O
49LFQSMnivO7MHOHYsIacIncDsUhREwcQEViJXkiVm9ThuEr3vwBt8kG8MXc4WzbspNsBspU8Pql
EDDN73XFcoKJ98zFMp9G1QPFOZ2tmuMkt7Wg5GzLiEVORQ2fOIit0QAk5lIjWjsnLS4DnhLap95m
0wrFfgkDuWNkvYVhKstQlqUBFktrbHmqQTbQlkudBO2sbu+4pUv0fjmfPZzWbtIoa6PzfEkL5Ot/
BF6XMCG8OARtYy5MPHLoldZst/mn8h5LoukqF/a6v4h8HdUDz4u7yVNxV2ZqOwB16fK7ApZOl+us
H8QcqTwb86sfE1gP5/VZoU7ddv2hqoNTTpDmjwFAsb2l/vA0CkFQJ5aRFMkDSVKoUX4HhoclFA/4
9lo69+oe8a2HZlfWYIYxycDgRH1FMQ1JKw4AOPtRQAhzX4BAERRo0b81R56gWqXSOEgART+pKUw+
38ABq1Js+2DqoMQy/Xhe1FGV07vo7PRo+vWye54SypODGMHJX5v81qdKKzVjcgyAt/vF0t42eYYk
vKnop4dUrCyi58AES9V1qb/z07KTFKhD3Q9gWmJSCErwf3j9a0OOkFgDg6gf/rMM2rHPrLf5GO/c
om5xdcvj2r6mvn/EAW4Sb50QfaBgyqaeZOsacd7U4nGHNyDv7i9qrtiEca1ac0AOc8yHWb/0K0S2
z3SOBdEab1ElqU5W0fP+xSoO65ajIYfXy2XgeIpFfiw5lwf1SribImqXMfy0IqMhD1/ePx8Rwi0B
aioFvgX70qGseO5CsNZBCSOsTnyzWnNXh0gF3HE4nLOv9PbdiQk5TZ99xEQ7UNgByW4J9NSCLY7h
1B7qBatwHxp+tDxMJuINBM1MB8R4bbgzpA8SLfc3Qq8i5qR2eeNgGqWa0ziLM2ABWu4jTpp4i2f9
65rmLzDv9oOUmccEQyHjkRn2WfQMsF8vALc9keoLCEEkUhUFZDw26ikP36HKbUwJIXyy9bVCF6EV
tXJpse6JrdNcTd74DLc6XIU1pAMgLNR1hb+nI6zcu9WZY1nwCla2ie7DPdlXqL1a3qQEYyZSAksU
7dkdNyeJ0kdwW2HMSKqhLzETNKp0N5Yptq3/QgqQauGZB3KO5FckAr5Csfs6QERR/q7rzop5xlKf
cOoxczrf1CbH4jZvxfiYpw2mvr++TV9LR2iYzmjRtIYl+65CddR/O/VZuWXP/GoAUrS9tlVgP+3P
z8Jg3zZmoabjZpyh3b3vmP151KhjHe0pA04kcla+c3NqbFCD86yyApDgehCn0/u5bOitygve2dmz
HPq/a5QPEnwUZg3eT8yGNPcbEn3AMzVm8xAxpqoS9DxRr9x8Y5XZrPOet9+D73eFHie0t5E62YrH
XRdm4M/xHpZcwoge6YX+W5ZSHdvFY8hvIJHnpt1GLk6NJe5aTEXF93RHcudduGckHNpTqLbqHu+7
Hz+0l5GxDUEDQHsQ3c8GzskHLAuNqz5RngV/mSSahDKH9jZ+L/gISOGWS85jeQ63on700jsNRnl+
bI+fnTu8h7C/INS9+1HeV48wiMltyjK6gNOB8aqgNIn+Y6cD27uu5P3dbfWxVCerU/VDh9ASeElv
AwTLLDDjgJX7QdSKCm6FlYme7jVLi2eJsd2NH9fR/XbbywoavPBuAwUrNhhkDl62FtK9c8tgyo9o
HdRcKfJSRAoWg/iWe22U/R1UrMFo/6t9NGndvvQHfp65lT2twHk3L3LIRFEPxI5r49G7kAE90yQ8
GugkUq248wc1Alqg2IESWqi9Uno7Em2l9o29APY0+faQvcLQZcZtAeqK6ArQl0J8xMZtTm8vZHaP
FgdlDCK91Z1QHQqCmXBit6rl7rU0rTDn1dOVYHs4aLYPsBlVgXMzs16HgKpydCC/62mD9wFKvasF
GNWoJJY6EOjEfuPNLbg3g9yaG6bfyIUcCZMQZwzP42SAgeWXyWPARgIk9wJoY3bSoaqf8koFbJYU
txtDhMjMRL6M9i9iYku/Ud1LBvUbSiK4mubp+94wTm6Bb3pDZtco0fkqYfYhBrcIZx7bnCOWMXQz
t7OTZy8MD3OCytE7ogxOWEM6wAOr+Ziwl3cO+gm0py9EG+fehUp6X3tOhy5m+OWeiltC/ExXkfMb
MWlEDr+NesUAJ/ZvPHMbNZt8J3/9D4IUYAt1xznuQWc/oTBmGNLOdPJ85ia+EDIrBMeu/0BdoZxU
zqaEB37bQnKmMNQaOK1kXWeCzfTnelpYMN7nBcLOJBDFlmk1zR2OgX/b0WYRdwoSCDCKK1A3/gGE
LDhurFdkuwuX8HhpK/qaGDG55zgJpiC1C0kCwbxuUz/8AB5ZpZN0wBa9G9zOeV90V+3cu1H2IBw8
uPTW1yDVAuTJk72n+WCt1oiR1XtR/pMuKOVroPmj2U+gP7FxnSpZL9zoyLLga49nKcmJ2fwoXDdi
AhuA4My0skgfwkZydETr0UFcMKbwCoRhTJ0edryZDUJV3YUlgthXCn7AHoOMhCpVxHKVb6Q0j1LJ
w5wZKieAEeXrn8TNwiFMf3FmRbeOYrPHRnL2eLphcSZ/kevNSVz7EdkpNzmoAyblsk/JlF/4FVQd
HTVdZlc6HyptLYjA5vEQOE5+IAmRQ2JPUh/wfhJktguDs7R109KqgJk6X3K5YFCZjHtWYcTjZQPp
+1XXhzZ16yTONHrOdtkos180T56OUARhDTc+G4mSpe9yRE4zpjxBC1yiQhW9zvoTHWduWPuJinUW
Bn4DOK5iNKmnsDVV5pQtufT/Zf9Clail1XkUg0Qg9swup76zlIJD0dCS9b//YCztKnve0EzXoRNa
jZRiZbRhWlMCi1dSQtFTz1HSPYiqTQfd8TzeEGi+CKN1Qnn5OS28BPC8O4EU92kwI2qix2wnvolQ
ZTjGIQNfSrd2YLmmjkZSqm30f3cGv27OwOeyvaeNhk4T6b4rkzFE7cFw6U+0SMFG7tfIBrfNqstD
ZgxxieFn72huIflB8RNoUydY4RJpJf5+r+fiIJTO3dQtLZMP6kOkxChaptyBoZWm8jXzJpyjrFQQ
Z0L880a+oAhYNlKjoCtkiI425B9gvUxmBV1ply1/0U2Ggb1TaLVj22glIfS/a8UQYCA+L0MA5zP7
PDJC001Ei9ipa9ljXAwyKGfgqlFph/T7C/8uPvI/1AWFm+vOnj9SSyKaQpht1016oRKwvHdmgYq4
uw/FDFUql3Pr+5ZckOfJNxgcrEruSqq5Z7v3emNgjFehBgwivNkQHtB+bS5mpbASN27DWCM01W85
bq3chbujHy8fOms83Cn9it3o6h5IXWPyC5XYjM0qTSuytFusuZNeEfbxsqvTNeFq80ruYndjJrew
akJcPCmE
`pragma protect end_protected
