`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 14400)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5IQJj49NipZ8M+awYasSTowGOcY2rynDmAB0ACIDngwbKy/y59zVCO6B
H8uZ8OVY4YOx1Z/2Vacp2ZiAQz08sIsIgXoIxDE5XNQ1zewo6CeeYkX/eEyypfbSiPM1GS6MRYsS
b+POFQi6qN2GyDX02Vir2MGqWHlxmxFlCKrtLhDr40prGF+MPGjybwjzg+qP5P0MqbaoANGzr76u
+mCBEup3ycPHW1xfGZEuBcgZN4E4ZYlWPpjNokF+wGqtWN0CR1MPIbAHVdK1F168EUbZax4q3xE4
kdT4z1gTZtqhgrIhPM1Rrn+h760k2P69e8HPXX1jxkmppXBnvjKYEOtkYI7USgMb7SjauVnSKZ7b
Pi8Nk8+e//ruIPeM8bXvNk7gEiVCiv/3FRG+r7666CC3UbmZLqv205v9MGiSBc7kw3dLWPdEBAJG
mtcCV47/mepYapwmEasdc3fgcw4y85DCigkMJICnOaMbnwKSWj0KS6PnuLmzmYRkJw1vZGxDLJzl
96aG73XLB2zJwEaOAJB5N08Vl3KbNuP7VmygomGoMnobn7Yr8ALmORKboNfq3HhV5w1mM77wB6my
3cL/E2HhfcZztNzmofnL7eEz4o6ZEOVI4r+byhvviMUzV9eknaox9hET8xqtWn27XoBalRVSSwNE
1zyeSBpn/GRSrgXLAp7/Beo8cnYyaBpPSZ5XQ4TAvLL8vutxNQenACWCDWAUvogKcLqkmKOJheeJ
F42ojfhQU5D4uDSXoPCkcvSXAW2axGHbJmWKSyF0XecUulfXElhsUSdPBWAzh7hqu1cKVkE5rUOX
AnPDq8K2Gg8yzBazTOll1UmJRi+4yS9xZTS0orRDlEG6YsGiDACaaGMaHhDUj6hzLZdCRw52mgkF
k38AW6n+03VicC76y9YgmTk1GU3IjoFmIiqgr8b0pPxB9ueMZqUalvcSIaL8yJ8NZpy6WPmiPZdh
08cdtVUuDnMGFCMngBKRbNSm2Bv8B8aSUtKvT6RXjnlghmK4ZmXZ8dcFRL6PMLIEJeaHjeP8w0UM
DwMKCSZupkvkCgwM/aEpd7l4S7lWXuZOl/Tsmnx/+sEkb+NI4lksRf1TF89elzi9NewgUR0LTnlY
dFe0gB2GqaQJwM34PNBdhOJDBwVtUh7595IaPEhV5WyDfTHTphgNY2Cb5I/DPEUXKPZ20KcDRh2v
j0Hkb6LeJoE9P3k3X3Ij+rkelkTh6K9x3MlmEJP+6Z4RLFgKCsYIl0wjhCgml4mUAmz3MycbtuJH
F7CaRqLE1MyN7gml3K8hgT4yR/tw9FV1leEJ5IPE7lelrNYA1LGIYKznFzQ9y82N8mcN6STQFN83
+perh7jIzeO+pmt5K7X6jwJMUTtiVRgZ+CF50fuf9pwHxK6dGJMFe5WbkAYGPz5/AascJpkBjVNm
v9EPe0Kpqezcb1EdG33wgxMMzTtO0vDwerqBK49XOQD+kavL00Rz+0c32EzIhFSGHnWF7qZ8BtRQ
bvj+88erkMFgrOWNUtK7KmpfKZMSxMH9+qglBIpdHGOEkgYZd62FnXRwGSY4/U6yLU1KC5Iuy8X9
8sLAWGMPUQZeGQwOjo9HWzmlIcjlIBKYH5yPp2zB0jH6BHBotmGlZP8nGpWRIs7u4z0eOQ2Oh9DF
KKPFLaHpU3dBgYOW9AYd6f4NMKv9fZQhwzZ75YlP885qWdPM8hLAJsJQP77QTiOURo+irJfHXI6C
X3b1Qne09th5HCPU04KtiJ8/T0OIEehyILQjD0Ilp5oj/lW1Opx6/AlZ54b6jxHmyraBkHGxl69z
ndRfpNHiW7Hmk+lmIwa5DI+Cl6WnyEj6/GsX0/eDspeLLLyF3SJGyDYNtAY5+L6Gvi8dUHlZ/FCN
fsRQhORtI7EyDYOxCb4V7WZUQV7rucOVaSy3CpF/7KdnlqiHxYde/VU6Pf3Ny8VppvUGOwhQW1E3
R+eDv2SsNPvpPhDvLq543JGfgNOfs4K/TYEOIFNCXet4bEnU5wd6kScuOh3gLXYxgBaMC8NoENyb
QW2VP6/PAiR9Ru3N9yn2RgvYG3gb0mVcOOwqCg16HLHmO15GXVdXQBZM4Xr94zRbzMMmJWliVFgT
tvDQUxPw/M25ycXDiHYcX3oozadWh3PtFdA3u5agSMbsZUozWe1SkZoioXBJtRWRF5i1fNOOpzqj
5dqzF/BaZdbvAbVxNQ2IiEE1TyAUF5aOfEyJlbI8Zgjf5kTzRtb8e6BgVk210ZPzu7PD97JM3XBO
WYe7JnWZdLy22yqCCzGs7CD+DeohmGalObrik1oQ/BpMz96yXkaWumIjHn4qYUgbGidfBgfWQG1C
78ZXag9LRLiTJqSxTTt4LNmjAVCeSRGnJCsvs2tYqaugcKIbhX2/hbreu7JQ+jO0wbbw7C/KBHdx
CBOtPS5DvZiGFdUz6DgHppQ74NVnTDWGpPxtXEhmbj7DWONi5TQ2eKMYlCnn10JWPeD7bqx+oyrI
FkeamS3BoK7Mg/4+vqySnt8OSdh2vdwMlhRICtsytKsdcgDrhXNQXi1EwHJ8jXxQsDatz+jaQY/V
31VoerYQlGbazeINOlPSz698txtJ1o/hFQfJnvQ/s/sZOh3cbzIdhr8YWB2xOxWFGshoZFvmw4MV
75Xb21fIYIzRBxppyse29hoI1prb1FnDZeDbm6D7K8xRvzW+Ak1Ha6WWf5ztptfIfJ4pyjObtWvC
lHfuPgHr3W2tq662WVZpxe53MP9A2xc1ymBkVYZFKXBPjqR5S9HQejhJ/E6r7TveCzz99MbUBL+L
XOlEGYcl5HaEd/SA0UmVNGVzqPycMq+I20s8/pnpcJLck5pmKyqO28ffDSBSZQBeday32FpdLOEZ
qHoUKkJOUVTXYQsnmL+S7I37orEyUWjx2W0OHJPTX6CPYUIfJRhLNbxJgFbe2usl69AhHFlNLoi0
FRwDoV54phx9da5lNzrZO33puZxrNcg1G5SQTnST533+pVmVtu46H1ncAz2aebvp2lAcQoZsquFe
by+WQMoLjpoEg6B2uGKIZTWBDRvCQMc+FeRPQdeaAVF0NmBUlyuxYKamaGErYph+KYDw71i5Bwzc
OmEQj9s7KwjePhTdPwPilFZVgcfF2jC6HU7x9PpGr7X8AFntr7nAAj0OHlkgSeN7N0bZ5z28ExaT
NQCugXbsRUolEfdfWRjTJnjknuEop3vY4twEy6dJikznbQv8e/3+o4dEVcLn8RgEWAQ4PbHZnK3Z
Kf8VbjmZVrTJ6fbmW9W339UqwBJRhr+QxlR1PHrd1074Fu8dKvo4hate22O8VE7FVxeU41WrzMdU
P769KTxVoN50A7BpJQExjaJr9KxvCYr2zy1672tM5VlH33efy7XHcKTHoE6YArZXlPEvl2D3DZqr
na3MZL/SyOSYDaGNwponoqqqOx+5ZvsdoHy2yQW4Efa+YnrqXbL4ZaOdEseppdGwEHAHbMeVd1Eu
zI8U1arKTaxjnT/I0srVW9oddQg1U3rVG2v3LxxoVw9qxyNAts0Tl1ui6ambKgRzsqLgznEz32JN
xDLnD77a/Amrrd8vxC41TMSenSdvdRr8G6wNQioVZiYevwoQi+ZpwpGue87T+t6NG/Lr/CFd+l8M
iiwS70dPIVnKm56K76tAwb9iODtZ3+fVdT0n4zNy+7DjXT4/gLXdN4jLRresGLOfrK4eM80kOC0d
8tSsnwfs2F2ZJnWeeoJSpwMjEiD7vOTNDuIEpNNdB+uIEq6X81nrRvWnulyCKX/iYOSQXuZxvUER
qoSmVgPOY1TcxBO3q4ikZG6Xqfql88LTDbILg95ceCsp8NW+JN++BAG1tEBnUUdot5EEI9/Qj7cX
3kLRy/J/7kSSdAz4mL0mGnuCMdlxtzQGPJwJdJdusoP6fcpS9gBjWUMwnJmdmbNuwY0MvZLcAEhE
xyX2WTiFhrjCZmMe46gG8YVI4BFMo44GKoQFuYFVuTfTGn3qeisQYbvDkugj0mnXyCNGSFhOaSFi
JZ4E463Iw+es8fyIHzasqmSLTrU/KeEer3uMFINNQ6b3naepVKSSEHsy1v1ELtvlMChWnLy8er8F
SYMe0KB+6+H+tMVcGfG2Rjqv14FJL0CsHpVlhDjAbQ8oyc4Q1ee7czrVN3xC+peJkJu9dk7A9Yhp
u6Bn2mI7XDsfFVLQ9uzStKsaN6N8UWir5jYlEKKtMnwdmTHMybXgtCvgw9iMPsS2CYWXIvUJOGDO
KXj+EZ0Onto65mNO16y5lkVXRrPNrKIsgD2ryovLqqx8PiSoIxZXrOqRvQl8Iz7lEpo7pdCT+0s3
ceqJqqLFv0hTmrYi2/1BWcFKG5rEhekm+j9BjEGX8WSqLiiCpzA+Ft2mhqBETxiqUy+HB9viZ78I
zwTzn9jEIcUqt078QMP05V+ux0zITf1kaBNSU/DaqUVT9e+zLfZwHETXhhzc/bauhuO9JwMfmakp
jQ+ySCe5Rpo1X2maCO2Swj8g4C3EkElIvrPnTrwUVu63aHRKMzRNw9nhcU1KT7jnPNa/PmC+010H
9rvc2UA0LUgE9oXVomMzieeM4DgVDe10bSd7ETDynqPdx7hVcHCZIjWj1S4QemZ7Uv3Ee4ZTinKz
lP4SGC1IsOaYuthJDWem8VFA6YqhXeUOxpMdKiFuXPrN5oYTT6++V/wjD0xFxbbwAwrtgs9r0zOa
eSG4KLgOSYSsnxt3SR33uOgRcKy2a2y+WHFpDNx8CiQq5Dja271BfYnz3BWxalIV+oykGJL9CI1x
TXXoR/VuiAnqXWdheePDc0nH39l0s0ixkUaKcEYscsD0MDeGHbnQ+xFbQ2lzyR2zzIDJIfOPR/vb
OGn0y+YxVvk2TUA1TSMVk/ZmZR4yIeKWAkzu05pe1m/Heh5GYDxyCjRZSIfnfoUzijHVUbsZXLet
nkIJlie5OjMhtk3OpyZIHZ9vunqit6AzRxlOtyZrU4jf/JhPPzI6xnBtcgpDwf5t/9z9jkFQINqw
k6L0AkPf55eOCvyfSLFMxOf6aD7BztDRkMF27Tb9uyVzFRObrVzSXqcMLElmItupztC++CLBcWn/
3o+bFlS+Akce/CRPfeYHoZBpDdl11kWhKToyPc6Oc76OvP26FA506DvdeDaWpB1tSrGIIKBM5N95
4YjGLSfTO7F2S4MPIh6U9ldUMsWi1BI1GUTEUMKVqaVWU3UQgxiuX8xyodmSUBQ/TvN6pjtugr9G
4qWg8qICIMv1bATHcDpxC6kbm8RGUOJqywQA/iVAMCsmfDUhU/Oq+SYzBC+dApa/nwl5Kp9N3deN
jK5X+i12rPHJIeMrX9OWEbslkqDMpey+cN6jV7WbjfZiSvkuPbFaevaV2GKLDLYU9wNhCgtjGpwp
SEl0TDFYV+iJF+5BODF8mCkxMCdYH46AY05900moBM5xw2go2TQGa0N3Kk0OTHK0kexdLA+iN0pe
/MwY1/sA1zbn05fUUSfx/qfMZ66hiFeGmjsayOJRvBINuhb/6ciAP0k9iH/dg2yn/eWIPxJ/3Dgg
y6vw8KH49xBU09uAOrK+ZyBWSFXfqPj6P4pq3cRZtRw1Prnuj/rwmVp8pOvpepv2I5yGTgS0gCcA
mvH0MreSP1gv/If4sHgUqvTQX/ZABUfeACxaUCYmiH7dFXRD5nZkR5wcRZTVThtBSLGIffjGso+c
cXhVe3nvXh+qA45O4htn9ul+2SCghwMalhfg3oQYNcD+MiQC1EEpPVxt9TDimkRYYuvugOq9LxHV
FGIuFTZUIQ2OP6kS43XbPDxTK3eSQ8HtjXbXxT15RHqfDWyFCW+y+ba7lHzcUWE4jCBDcEusejYh
oTWe1XJAB0SHU+2a9TKEO9dTupNVqX48/bW/dRklGM3UNPT9aUwayXq7MK6HLWVmVI1bDC6VoEMx
TZJ1Q5Go0pHGKieD/XrqLZ+zsIuKg2AzPiOkLc/bzNGNxWb43UCCCXa4CJlwdcG03c12DGMNmK7g
vpafh26bjFSazD6+nizmMVr6WEgcD/mAgAekIJvSamXGAD+BF2oIn7/BYzf/GJhAi/Km7V7Cx8Zd
lZWiWUzw9/kKGXlOJDrUQyhfWPYSaSUgtCZqvuW6mcul14h6vyJWIIyvJQiK6Pk6KdLltP3ENNL3
2VuWtY2Lp3JDUa7DQeq6JXLSNFbpF8RK/Y4kMCCvpdkQAamIfuQJcpRFpilzG7uyaOc6n50Xg/u4
7VgUf1BucDhT3uHdox/2x/yvYBhtqh7LKaBVB1uAPfjJhTkl6+xyo/bncpYK0HcJVKo1n/wfia9t
v5K/Xvgu4sPk2EqSnn1IW4mDJGAATdCOZipbawx1f5GT8iWtNxLDpMU8TMTfYj8JlztTvn8pPgnc
240CNCkngZRFUNP6FfzuSHzZfl+MNtIaqGGQVvtBqeXpZj/z3euguGwkX8Ne/t9AGOV/27mV99f9
tVe29CwG21MOOxz/MzI3mselO9vLGOZcc+eQ1d7lASYnuAOHK0FgMtCn8pKAj0MtOv7+V7xAckdu
9t6f4SrB1pCzabRiybACtUmz/hI+DVJRrbYm1adLvJDsuwIcMbldjrfBirBtiz8a4/FfTYvauDL7
2yyJPBiRdfqN4sKTlv4QNXLRMKzk15488gp84eYJO2UAxPZ2WWBaP9qqUkbUk5Otfc4Dbbx/lEde
LPRkUFDHbnZbK/LxQ5Wmzvc4ZmzH+p7cLuvZVQAWg/VK03hVgr3lYyKfNH+qd9VznD85XUht8Okp
GSeCCUaiCFAeaMQJid3U2GJyiG/ulZ6rGDl4Au+9iDLrv+wY1L+3B5S4hRVnOrP5tcEGRL4fXK/T
/nkFVqMjfUL+mhQF/rcrqCUTRgpuQC2bgs7TcgkF57m5N6UHQjAGOq9cmMHf3bK9I97R16OS0XYL
InrcWLj6AQ44KmssjgXtg1O6j9/gM88C5NfpJYeaui+/Pjf+p0dSzP4nemG+QPMrnep6/iWq5b0Z
AODvD4dXcbKrKn4cHmYUS3mwDWbAj9a1WfQAV32UKV9vmSbOR82Te4/0JjxSpG1H4UkFCEinYDDl
0WBGjtJEP5inLJR3JKU8E9s0hwWwqAi1RlIqxYkjaufRW95jlbk6L09j43VMTw7A2RJ1gVa1dpjj
h/mmWg0GzDrRtwQOXwe8NIiLx6/GPAfpszT46kEWts/XhL1R7lAjDZwBRfxLFLLHceV1EPvx2hTm
PRqo1UG7SznnLJ3M0zw0lWme6+G/eLHuT7wiq0mH9SGr3tqn+0lEqF+qO6Q+Tii1CO/uhrvOc9GO
GiT/UegP3t6vQguTESahpsZ7K+We+ww4imirpBM5R8vMl8eZsl2rBJdi7MzX+2zGXwhHRD5O1gtF
z/N/KYCUUQqkOt5BPxREAe2XRJdsqxNS5VUOA0pkjjaVbChu1GH/OpURQcWwybaidwZGumlw9Pup
iSw1tSRswcdmn68o3W8WW6bCSNAfDacFbc3C+4rXPXfxYcPnjDEYmdYYrF/6LSJS2U6r0Du9t4Jw
+opHnq8H9ZVUtxRUq082fAOYSkboqtkBc/STDsJQUFaBGpwQfwgwpT1jQgT0AjtnP5zT9Aauu13y
c5ZelsdRDZWCXkuCcO5K6quMqrcclsyXMqqxweMY6gH6+NOBu8dqwndeganEkzWJ67naSTkyeTsP
YPrGNybWBC2Dw3l7fUGtRycStMKJhvlXyClHLpIJSPXgpszApBDkjTaRzyIq4kPfWDVPhm/whqJL
gOfy6aC/c+ZnEvUh/lFWNLlFmSKQO0LJdpygK1JeP7fu4SRTdVS2Y5f9B0QXjP3viObWOxpBZ7jw
7WhT/TuEyHBEm6BVjJf1Nr7GRw4zrLA4QSkht3KWXEC6hEU0Ho7OCYW/1WhOHk2yMyKDI95tewFt
pCa6TCBMhJyONcYONXPpIrqzJED5cBmcB8Sil2FbnK1ciDrgrjhA5+ikh8zk99vrQii57ePTmMcn
J3xzCP1x+Jyw9+HHTtAWDQX1TLL4IRYuNJU2QMaAhhY2LvfrunuqP6AirotkagymH0bb8Kfkamu6
hGHC4tChgJ2wewmGHGA5zAiAOH3WG+/LIxeC7d1M1agtZ2b+amTHG3VdZXLIUNaTzuCES+/QS7hI
PnDcZzouQBxEzPq8TqECXUgzu8L5098N15LUnCvUnsQzxFoR4WNKHmRdTsJTVGEDXysjWTD152A7
5HS52qKrk1bEt+q4JEdi6PZE0rmam+Tdde0WkSNkebx/MVA06T1H8mAwWiYjeSd1fHYdyV2bve1B
HwVh4QUGLyark6IKp7Y5f5dcOzLTmH7Cxl+90uF7R4XUy8gXBFDkH6kNJs0stpPwQ1lzfhB1TXle
9ZNJRRMbemYHzrLKAzwM0P2Gmd/AZGmiCt8hbR6d1TdaTOkCZd6Wtks2A6Fo+j+zitOzWB2R3SsM
aleHi+2xaYRN1IyvqQzuKOAFEhcjxvv7wASwoObUDuVO4D3DmbcexAVX0W5xN26RszZj3Ugv9V4K
dzIxVZzI31z1Ar4TkHsWllLcE2BZQ2azxabS8dkvjHc2/nGBnCqakCGgQFLz4bCXzXVKS2qKHbMn
nQ63Frr67ZeSJMwXVqA1ynirvX6tav444LsU1CGSroHUo515VITR8/5SvptgzKDrEQUF/khCvWC0
vnAI/xhE1xZGxBdTyeBx057T54qdUy5XIkgDHRclid1TeyStO+xqTB/6sznPk0jdIpEeg26NPwbB
UnSIR4mZWGtlMAqBYYHF9hym/4x5/OEy3igRObjuwz40ebJDDZKeU2IKdE3TZBer+FEMIj6D+jTi
X8TKE3DEpP2cF2GM/mPpfkFV085ltyHFzdYNoc1B8v8EMLbokojbEun1QruwwuBmMRqDc3WFe4kW
As5SQO9+qeapTR/gaLt+IlXoSdbIvIQIua3ed8wdJ+FMzjVKVYQJduF59aXxhOjdcJvcakv5u3zE
QGV6YvyPoGFjnzob88Tn4LzUvpP6SK0VgLmxQDIx8IW1UGKQB7SVFAf2kWQUUmJjFPPK04dj1nf5
fuwdjjsN4TZUJMLlCqdAT71oxiFB4JxmTbqWa8GA1BZ4wxcuuone42TydMNTz+gWJWYPSi0D4WU1
HdUrtfU6iCWSDDCBVCl/7CfMlp6JxaLFGJwJxnt9icARGFQElzV4AWMbQ6CXmzcaPKYs4MDfvmPE
2mkfoRMAvEplWYQpCZT70fEVqIW9pCjBXP562CsVvDSkNTAFdOPDunYPlYOwzSvVJosgjdy0DDYL
syD+viJYRyY3Ho6iVXMvOdohaqs/91rc5rt5D1EUFx5sMdre4VUnwwiXsWwHYr2Ie1d3Vo09GZJy
T9B1Ah3Iw/p8nzdD1t1Q+83gjEIhT0oLnlVmNGg4r6Kph8682GwHfMQuS/2+l39Fy09l+eZ8lGiW
8/7UN1ZWLM5F7rZwKdklwjb1d5qJ/CsCjJaPBWJn7H5BaAfAHFfUnUv0CqytQ6Yi0UFoBrdM6NfM
KyboEuvJAGCLQtgA8HYVmei0fWtO2YjMSTmSg5YhP9h0Q6KyfnIcfJyL0WAPb9WxmCSBC2ZLbHIu
zwoqc7326BoofDvPWZCgj2SLV9CZwU/FsLvRTOcYjjXPjzxHeIbnnXI1ya5qjoKk+AoF5582kD7R
IJG5/lkC85ChBNa+bpVjho8OG51r9LN6uv/V1oJkbjOCzMokWCUW1HTNgrpvM7DJ7+XtkO+BCG3N
1M5zDu6+aPC0lIuBmqmzXAPrMOe5XSrvA2ltIbfvkekspGl4hrUUo6gNaPxXEO20xn+1HZiTAtIt
9uJjTdP54PhqUZV5NieaVyIjevxedg4fYch14zswsfMUnBM7EatytBRsvlgKPust9gH7Q0iwMcVl
9ggbHWPsvl2oe5de+X4TIuunEp6fgzGRPu3fh/Uph0tB5vt0NnacIVnHITHttZLBZMOLf4gjPtbF
MDVIdDpgVrzZv342B55Yixl4aXu2ucK8NZmRLHkaajZnhz7KpQ+syqRU8aq64YhLuIgWWgYAbYrj
coET7WR9tX06HRkwx4Pkj5wS4LGdaxXtNv+rtaHJKrxeXG0l9sdEt9z4/4zMVWPw9EpDwv374sl5
mTgYWTmQLmYC2f99UHxESAuHgbATqrt5e4vnzVVZ/nSu+LJI2uVnUmrmGKijdWV+dlOzmqBo7GKj
ylmQFpmRijRxfZHhfFOBBkSgMHnfWcMJBh6WLr5PYZA4dduZpUYJgX4k9J3Mo72M5qiynGT6zNe8
B1JXQptbCw2asJ1VQy+vyKAvNJb+sUnX/civ6Vtu1QyKi7xSSN71Jfabx9zN5/qAhNwOVlKUDOrc
AX+GmcJTpUxTBhc9NvCb6PZgdtKztV3mfV4wG3zhqhsiW4yZlNqvgxDrM54UCSqLDwrm65ytb4Yp
P1Vo0ifQJCM2Nr3Xmqe8JQXgxp9hQlaH3lg/hfIEKH/I0+W7pFfc+CX1F7zkgdsjxbouUvzT66gb
gLx1VFsTh/AdXCLuSKvRBpTo0Qr4OAv+GZ8C6rS8hv+qDRAmmfQ6HFhytgTcNMhL8xnab/w1Up4m
+qcrlYAdxt9ni2OkoKmeFNVpDv/j8CibKs0dGGxULqzD3z4g0UY6FrLaFWss8BUEUgwyRlBUj6gN
0FUKELB0IdD2wLOgnR6OjO+RE41NwKDFKtcO0HLKTAGHAwL+mX8zK1WeKp6/zidL4nJnSdkZbjwx
mCEU8K/JpX4aLyaBlPnhIM24cfdq3KGuZ5Ecj9hSxl/e0AqjplqSbwX32a/PDRluaIVQVx7UmQyd
xKftQ3NPy4FG6qFJdKV4vyBNsC1Orh6Vu5fQYxIrRAyL+Akwb2p53lX4E9cDEABEFpFAlSDuEhHf
6DWMZ/SzWK7KWD331YRUnYvX+xzXEgx+pxhglPW2wsQFHHtYc9IAPbAFRm2bf8A25CpF40Rhfo8s
YTvapNsDXbbOkYs630ZXBchymBInIZ6xxUWKQjdMGUhkBjJCC9EWkATpjAIBZ3fUerKhMF0AFFWs
R6gLV9GV7AKEj8DvRM1eUZrU9pst+uYIFwqWcP/9RkNTTO4IhPijP2UA7MXSYWTmBhtsKpu43A0S
tUI50W/n+nEfvTB983OwU77C4V78I1Uh1PbqXxSssNlZilCgWzWu7o3oOcjCMEHKzmqLN249bCNl
NrmjedPAK8xdX/vsUGuZw410aAvSYjCWQgkIWTVU6EL7GqXnNC8E6x0x85aqUJJo5be9t6bZXmjX
kT5Wyg4imS83pWpmiRpVm/4JmZekUYSpqpOo+yR1tZzonct2dbFWNKdr2aU3RLiMK3Et5JSQRa2x
LPk+yWXlyViEjNLpTJvFMn3POlSR/uGMWWjHJcPFm7SImwrU/z3ARxK7IUID69xew1UmVIMooXJA
lpXq3/+Gm1WaTRSA7hMYGNVMizw35EhKZ/oWib1PQObB062xrtUS7h1/+6MGBR/XT8X++bKpAxMN
ehBxZUa7FjAnaQRlDk+zcscXOolmAnTxCQwEKwNCfOpRxVK7pYaF3u1CskPp5W3ACNWDzbskjvYb
MZgkbrTlI5GaUe6OdJx7C/sPcPplgOZ4c63LdWAsasZKmSliTU/tXyi+ZEjRkMCyNKbCZTOP5ojC
9eQdHBTlxJMmx/gfKypqJU8yAZofKuBy6dpmnL1EJKoGqgQBG8jQib4xC+Bey/oO8pxG5V6hyeT5
Hw4MWkXT6FciCKPJN8WHrSsiY0srRFWi2Q3cJhob1iJGYsJ9his9C+Mlw0RNU+BtZD5EnSP4jc/v
+2vo8rc8yV8A6q/Rm7u3UkZaOVyIIQjz9Phy9N+vbKmooqp1ccDf4xLOFCLqnpe/Jngj5XLEAqBz
WPM0kBCOpA6x2Ohi+WQJuUWn72j3JlVQocbvUXd+tpWjh2TRmJdHLbQjdL4QFvToTm9xgLS/TWHq
X9D7eNeVNyqPoPZv+nZH2iUIJgfXGKJ6vku67E3Q4X0P8Vb1Otshte498ZmjC1vD04fuk6ihoZw3
Z5qcZwfegtn0yaxLrlq6nfejyk2AjC1Xi1xpTMhqwTUt4bSgzg4RAUDPpxskfXAQUngtjfFsyoJT
VbeWDEJeU5VXg5c8CEbrbp5pxzh0ZVvtml14ImbGIR01LutkGftGdjlf6B0nRckowm3+NSQUHn+X
klidCS04qBEUk7hCbxFSX7MgoSYD2AJgXFMq9Q7xcEogzc+pokSRkwChMpzQ9SbYhp9JDKmOnRSG
SA7sXJWy0r8NOsxarGUN9gaHWZSO9c+urcAmwKX4h63NVFitiIkF1vBB0otigsYJyRuR/snsS9nk
eU+2WPJqOzEdfwHBu49rEX0jul9m+AAcs4W9lDUbRf0sPsFBEHj844tOyqH6hGURQnkgUJfJHbsX
Menvywi8PaUMnSW2Ur9TNIITbD6bBBmIPf5xdW+JSe96VW5WH6U4PNJie6tTtvOVilwm3kFgqy9F
fP6tAEYlS6fIk5trxCJ7nMCW8JX3O+REaZalIBcQ9ERHrO/TDp4G4rD3XKN0nxOQJZyj4hBAiQAC
InX68OW9xfTChG7vJbNPhuLCifmPajTBpCuAOP56HGVSeUaghp+cmi8Li3jc5Y5oF76bUILLHPIk
GNHKUmPu19As4dlr10W096pGKQ/59Hvsz9vSTdxGdYGJUvd21PecdRUadTo+8WR3a37f5bivNzyR
IekXeFNr148H/8Lv+SoBJUI8XxSma8CDab8gDcDcRm9BDa75h/hrm49qLFed00DYomxHB19dnXC6
i25KFU6UivaB6qIJFGwCoo/qv67rCV1WUrZZCbKYBeyROMbMwK8maYIBPvvtr/glLV+gg1kRDnhu
qaY1bkn4qEgxdDIQpmh89mu0wyoEH2IFMEUmaf874bLwKAQKhISHstaLaFIxHQZ0SZoR6GOTawn6
ARYg5erl0YsAx9YRJG6KF93WHHl0qVE58W9Tl3O1z0g7Lh9FdDpMA+PBfa9BcSK+YLi+7NRdw3Ie
f/7mjazUDOZmniBWjB8jkSZPjMTMa1j/WJoJkdzoAExTr44on1jo8xyaNXxlQQYuvH9WBibDLKth
em07dFcDRAYJhqz+qfTDrwfbAAoaq+2DiPze7lRxSH8JL09J5DAXSJZB091wpFlYYrD3sOMBg1gx
C2lNZQqTgxA11wi6ZfqjU2b4+nybhhCUSZTXXRNRCOK4XxueFYhWzQ9rNTXIhvh3eZuXwpsALQh5
DudikkvuTb86vG0qaALQ1VLzxKbbeudQbxNfP3IbhFhpLMo/73dK+k+5FLdj+tpCTEwkLapEZb4H
a722QOfRZC/GJz4v7hfUydVkn9P2oci0x+BPctFYdBPeqyWmH4FfOgovSm1sx9v90uWhRtSCTbYy
nfypRewhLozXeGT9xEhIa5Dmm6tLaGpfY0+jrV/rCMiDwaTwnLWqiHLaiQYn4XtWbKK0n2pQmOuv
thN8xq5fVTXgf0R31CxDJWSq4613hhcP6MP4+12gGwaUGT1CYO3CCgy7HenpVBpaZSX9B4cdUFnG
xajuoNLNhp2AKviETaBA/yHRsdoG7PJoGEsGRRodeG8rmmhLLGjaSJZ3nQYjpkyCPDoCask/e5Q9
62y28OtjYzFb1JT7mNCvGIKj3u44LgBXhMgkUf4F0OMOkEXhJV+PlNp9aIxz/uqDUDNM2zIF8lxH
usxn+GjKEB8Z6fYwyecJhSirLjLA/0IyG5cOsZDinUzUVNnIBBfVuMS0QA0WFfLaBoo+ZzZ+VmDu
cLJB/5gjKDNegocIRn6ZHsMHPn2JX7Pq/Xu2u/X5Iw8i38LYfnXw7odGZIW+jewpgF584t0gvV8h
UYZUlpOQ72W+hHjWI9c2c0PfQm+KTSN0EHK8UWKuM0sml1KwEEbcNWOOG/mbgANKYZ7z1dflNih7
8cGekQX/eNkGZutEuaYvrXky5ej51u/Z75O0ZD0iohy37wmFOUfGAUxVM63hYpk00WAX8fXwCUjY
6GBJlwjcQIUPxFl5BBHnUXdSsE+AjH7sCKH+gKUEEYVJJanmb8E3IlV4V8EHvFBcf8roLCPozN3U
xUihpWuODXmXNhJt6nUMdzJZcV0XQwTfGf68eS0/RzEz7E4d88MYbF2ephfU8F4kXjSeUvdx3u9U
AlCXvrkRW1JyXDARPZhs6c2LEeoS5/u1Ddhp7ZHRWq2pPvRuohrbsOH6wlJFlkKm8cFMvuf/HpOD
MMRArxls2fqASoKT24GbQfkU60bYDOnvZyoH/0tMNKS8+KKYE/73SiOJztqu/IaKdM0IgLJU1fTV
qUH9LJp3KSRCq0loLgI3UssCFNOu7mZA9El6+6MvtX5dqNBph38aBvsiGv0JpIB0pjoSAsxvPzg3
Z3OT07PvmxoHIO3fzjfjPS6PJSMHxDUl+xztGF4+yucM5Mi8+hZggb6njxzQw0kcooUKgQRbRiWJ
yWe1UYJZoEIT/zyV5FQOb1ThTjYBj04vuFisVsnsX3EV6XK4sempTnkQHfryGxcBWuCof5WN55mx
d8tjEWeIabfGczYblXWAkqXM2d0W1iDqKa+ivgHrNi9L4t55tgoSGW8l7549m9dyx/tapSARS0td
WpPNKVjAkOtawSHLjFFZfO1u/5J1eOFLDX0h3DNBd+dly6Cizd1g4ogG6uGinQqZNujNSwP+slqG
VhnZZdjlXB2p9X7TjuugdT12Et1bTFOJiVxGUmjM6ABcxaWsy6cFnRyhXkojkqJ2hMJhLpBf9dX8
eg/qozcpiuIz20H5ik4tS1tmpXqpyHCTC1kM6ZOfbrMsPSy2Pk2OluNMsCrZ/txPIokrKtb2Ufw8
9L5Tsi5sOPxjz0D+qViwVt2kzR4RdpHO9eUUpiTqi66TgvsFtgSEffThb4CAT/Y5R90L+q1R3/Fl
+ovxn4w7uoEnNgFWyQvqwytdzwHK7gbzMbzL38XmrzicIM3lIM4K1gxltO69JZWJiZIYPIU0yni9
PyXxYSEJ9fA/A4qJPq6DRTDTu5K4xkd75JFTfEmhQi3q8Vvg6PXX6CHVxZT74gY5DGspdKyRHQYy
X66jKnukYncWQJOoklkjKWZ4K/u4RyQNJ3ixKGXOS9yW9VcDRkKbtL4fN4Sa76QfJ7k/KxmRDNJK
Ogzu8y6Txud0pJm2DgneHLhJe3PjXffVime0WO0vUMDH6QJ7ujSgi7KlYh9Gz7LD8avCBlXueo40
v9qaBsJdfGmqlFsFZICdjpPRKUCG6ceo7BZQaMWizDieqCh17OPVobDjAFG96ZrhAY6gPPgVc1CT
3VKehNrbfdiVMF2d5sINyvEf98MlBcMIygbQ/t8Zv5Y5X8lhKBcIolD0Il80YNZbmDFrC87gXsny
3yWiztz544E785QW1UoJkEpGpLnH/pAkdSZsBu83/w/UhW921HYH2WKfAn9Nh5AGi0cnyo+BB54h
KjDeji17QdoeziFPRmRSb9dO6uo04XG3FpZqxQznETwZz9WDGoFN+jwygTGqiC3QvIflU5saDo/r
mBrVwp7y1+SF//f7UqIXPYZoE+0NfCQEVFV/3OIPdCO9o6dslIP0o/sC4sesp0mVS6gGAfzGy7BG
5LpnPESFrnhmdr8rYX7Tn0LGGpgN9C/RCf/w2LMYVB5eCM1SDwSG+qQBHjF3vugw4M5rJjscuHN2
wvi+WPqmrB/k4lv9R2oTZQa5X8UZ6U65Q/KnAZUm/+MFBnIWIXa0BG46dcIr3C8bqve+Pbz+eq3J
uDUN7FAf4XCjJ1yKvxFpyaU5C9LFGZxavelIBxTThncDHL00Wnb5gbeM4cAE/ExLWiNVKghs65rH
SvDEoFT1W8HUYQAAGme/LKxEU5Ww/jPkglS5n2/uqO1VhIaNaSTzMIAfijD1zS7a8hSLV1GRJysJ
j0CmY6cU8oVqIU1qPClprae7VRDwVLDwFXqH0iBcE5ioV6+5jrZqnNN0KzufCcnteiZg5Dn0aT2y
TkYLJWt8Awm2KsVh//6l5mkL5iNlV2ejvLF+8iYm5Cg+qChgVxRSGVL13FKM3+UJuhrMbFE7NEIS
GRYYaN8KXGD9/uiPg9TXehtITx+EkJS3cP88opSckbgqcsVczqi2zdeyxKaEBAFo2M6jQ37v4bhb
ILmjxdk9kMEybT7S6MOwdZrMfjHByOqo7xCGDirytK12rYpQr/ZxV211bWyCdEWAM65r7HEaNJoB
FifJjgSBu7Q00BAD09M7vZhsZWYg1XDE7VVrbo9/E9VlH4Niid2xLgLizedREUErQsstJP/kCqgp
TjWR2W/OoDRRhK50Wb0SwbDuwhNS6WaffMxhtK4H66fp4CjLGHahNXd8lBPRcYU08k2l8exEHBzv
jGQlgWLm/gtUKnywHLuGKXsXtm9jOaMQNHMkJ65K3OdRrWV4rpAacKIn7ql6MHhr4MgFk0tXq5ar
F9+9dcibBQMCfZwRgJPORKL1n1WdhUUHWs+lGkPhadXXo76A51JVz8L3JZcS7ahWChsk4TrNQuIT
djGbJ5LST+8cHDyf+WMjy6BUl0SS/1DJacLwpfphGZ7NiKeF1R2dbOn7HvmCvcheNEUHbmP/7X87
WyiWgdQOceewAfC+vBjWvGnXQIW7HBLkeeW8jDvXo1a0tU6oDwOjeBbYUNJLOWGqAAyZn8D+sJUd
+V6vvz0MTqVf+8+s6OeR/d4Eqgl5liqqWXUgMKp1hZ+OqVhxqs2Oj4ZhA0cUK0KP6TEpV/LhTT2g
GSvwdzqDRNyQl/iEjGQKYy9R01X4kAQp2Z6IqI+V+EhzXrBMnX5cuWzTuKnH9PITj+f2MTxP4+nj
uqrow+yuf1nHN0Dhb0XLBm8KV7YJxMP4uHXmIYkNmRnzzsPRdDv4plK1xOArMDtmiIIEj+AmxPq3
dxnGdTwaCTA40gRqLd3G4e8QOPTVLYNaDrrfXsqefjDDl10ZY9J9wHCuxrtyk1rO8cWGfv3+gfHn
2KI9pmTxJuE5SzRGJJLLpL7nh9TLycOLNyq+eaBJb58tCtQ7ufbPr09gd4e5e9UhFJBUkd3SSgzX
z0Bn5KvgbvJdwV4Q2eilt573cJOF4Zo7y3TaGGsbVtqZ2RKXSu/OBUQ5/kKZEpQbADDpE9TtW3pq
LnVqNPaJ07F3zrq17S+W5ITqVaIop6A5RN+sk5Uq7vG90SjPeHx/C6FvUYnUF3H1nCn2fhSEC7E8
ifmO+1mT4e7Du1FUCd2T0prkUBePp+3v+5daYPhg/MqC/M8swbS1LWbJarA2k616RQS7c9lkV+kQ
NBoWIVbuhrITzxVN9/59w9ZOJjmyKmOdYk24y8qMkfi7esWlJctDg3LJzIowzocvS36Q4VrydCvx
iKUpSrmW5JmRM2T/pTbG+ZgX8964I9miAeDnvJo4b23azxhg73ZK4p6tSw/vhvdEkfpDf3GrrO7C
jxOU9JtiDgEA5/VMDxPBw+QdkR35UbApcikcwT9urZ5yf5KCywesNXz3Mpb6cJSSFeAYHbAe+0Ab
37yFa2i43sITl2OnXvwBAXm+Q70pcNrwYE25YT8aKlkCZ0w1xu0LVlfW+SkPBSHHbZCFH19BAhj8
S9upCIvil8zIGV9F5MTIQIuT36QZlaTc87TSYAKshghsje1t5GN5t1UX+rc3LeC8xFmN2EaRawFQ
n2DxnP5GRCJCnfIjXEzj4EDtqV6E+pzPWFiuugr+LvuGrCWkD+mAIEgMhPxhxlmTlnjhxShmTf3+
12x0nOSOqOrzp1AhH5x52wO4gvovLcGx3rPtEvgBuDKG6k8ySwIKWd0NGiKk2m7fiYbdD/3bdwu8
/Ld2G2pPMYNJ2ZXAPGvoJWiRvGDMnOlR3qXBWSpOd7Gw+hScU8ewncLa0ZPbmqmImpq7/lfN4CI1
m6q+McvFQr5VXhaQ+Gx6UZDx63Zd+QcyGSgwFKbdt/bFJuZCbAIC/dypGiOYJKmGKCTJ0CiY9wII
qZIxtZC8uaqrGiA52mfhGZyhZYQgQ78GwShz7S3Rwk0Y7ZRgsJ3mYz8ZrJy4FOEgLKAU0SWgfpO2
jXxIP4ItR/4I46gXPTGLQPfbulmK993i4N67lDLdHsWOieXR/YcnDMAP+uB5YdsxLoxDezAIYjmj
Kd5bC2OxpIEqQMb+qYj+roJJzxjuytztSpm31fEm9p0VWOR37l/d8hCIf53hdH1V5BFgTobAJNsj
mSJv2p+851p9eajHG5+iNMs3+KKyjpXQUDP1anfhHDK0zAjShU6Cpy98VykSifmSY21u2pTVy0w/
Ky6NAomZEjWrEFHP6rWD8UzGp36kt+x6pcdd2aP6tNvTyrsO3PjiMj5JI2MIjVO7aZ8QYqKmsUeB
AhN7USqWiO83rBu1wPfR/W8uMpS4rLQstrR85vJooSW/YLfNbHtm7dIEJORhG+/nVlOVyuoZWXh4
j0iTYvZAm38TtpKunD2dvh8ycy+t/uvO4osx7ZIlChsUNin7Q6k2XUpdvrGuJbLGt+BkC8edJ+ez
KcVdSI2Qf5d5/63ug0Yefzc+lEkZDsWP7cbV9fnjwpFzsGsUWkykG2wlfPmzfn1wgzo9Nn2kRCrb
NKL9OUfVe6+D40Spliygrleaq4iU20CcksgViK5pQCC6iqKEa4F2KGobSYmrqcIvQiGrUjweJGia
qGA5tIOf0p0ojygZq1BVTk5c9JeHzWyPnE98b9iD/lIlKrK8I5RUdocPwtZchBRYn5iMLf+Whc6t
OTfZSRIkpgJWncLEkzzEucFCeGYEKCUjZh9hQPGyNPYsmhgmecVHm6NqjysoSCl/DNYyKFGFmc3u
e0BJbcnuMBP5m65U2DgKtHfCLNcLQx6rKbp7XQ9xvxQqGV0QI/eYU3DxU9gVOvKcKCVb/Dr4X36v
HmBQvMIwrFMl+jElp6oRszjnUU5HqPnCEiHECLIsaHqbQ7/rY3ZWEHArDx/LmchaDgMF6Qkr+HAb
GwNM8YoesYkQSdv0hIupTEkPi0FoU22QSz5dFHlKQdL0esH/uFpOsmKsJmLdBM/JxOZqD1Mu4EJ8
0sXEtfunNSfkJ3byxgtNZQDSteiytIrGVo4fMDGfJIw9Qb1BQGCpn0vzavCm3nC1PTIAaTWD6V4W
2q9bAMwoJt8xETTd7W1AFyQrP6JLFMHNskqZbXrbla6oNO/po70NVAALpfwO7vDrm1tkTVPhgVRB
8u2FskwN5jcRn5ITfIYUUVkh6jvs63oGGVB/0UF3cbb6hbkt
`pragma protect end_protected
