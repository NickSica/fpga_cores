   input         cfg_dout0,
   input         cfg_dout1,
   input         cfg_dout2,
   input         cfg_dout3,
   input         cfg_dout4,
   input         cfg_dout5,
   input         cfg_dout6,
   input         cfg_dout7,
   input         cfg_dout8,
   input         cfg_dout9,
   input         cfg_dout10,
   input         cfg_dout11,
   input         cfg_dout12,
   input         cfg_dout13,
   input         cfg_dout14,
   input         cfg_dout15,
   input         cfg_dout16,
   input         cfg_dout17,
   input         cfg_dout18,
   input         cfg_dout19,
   input         cfg_dout20,
   input         cfg_dout21,
   input         cfg_dout22,
   input         cfg_dout23,
   input         cfg_dout24,
   input         cfg_dout25,
   input         cfg_dout26,
   input         cfg_dout27,
   input         cfg_dout28,
   input         cfg_dout29,
   input         cfg_dout30,
   input         cfg_dout31,
   input         cfg_dout32,
   input         cfg_dout33,
   input         cfg_dout34,
   input         cfg_dout35,
   input         cfg_dout36,
   input         cfg_dout37,
   input         cfg_dout38,
   input         cfg_dout39,
   input         cfg_dout40,
   input         cfg_dout41,
   input         cfg_dout42,
   input         cfg_dout43,
   input         cfg_dout44,
   input         cfg_dout45,
   input         cfg_dout46,
   input         cfg_dout47,
   input         cfg_dout48,
   input         cfg_dout49,
   input         cfg_dout50,
   input         cfg_dout51,
   input         cfg_dout52,
   input         cfg_dout53,
   input         cfg_dout54,
   input         cfg_dout55,
   input         cfg_dout56,
   input         cfg_dout57,
   input         cfg_dout58,
   input         cfg_dout59,
   input         cfg_dout60,
   input         cfg_dout61,
   input         cfg_dout62,
   input         cfg_dout63,
   input         cfg_dout64,
   input         cfg_dout65,
   input         cfg_dout66,
   input         cfg_dout67,
   input         cfg_dout68,
   input         cfg_dout69,
   input         cfg_dout70,
   input         cfg_dout71,
   input         cfg_dout72,
   input         cfg_dout73,
   input         cfg_dout74,
   input         cfg_dout75,
   input         cfg_dout76,
   input         cfg_dout77,
   input         cfg_dout78,
   input         cfg_dout79,
   input         cfg_dout80,
   input         cfg_dout81,
   input         cfg_dout82,
   input         cfg_dout83,
   input         cfg_dout84,
   input         cfg_dout85,
   input         cfg_dout86,
   input         cfg_dout87,
   input         cfg_dout88,
   input         cfg_dout89,
   input         cfg_dout90,
   input         cfg_dout91,
   input         cfg_dout92,
   input         cfg_dout93,
   input         cfg_dout94,
   input         cfg_dout95,
   input         cfg_dout96,
   input         cfg_dout97,
   input         cfg_dout98,
   input         cfg_dout99,
   input         cfg_dout100,
   input         cfg_dout101,
   input         cfg_dout102,
   input         cfg_dout103,
   input         cfg_dout104,
   input         cfg_dout105,
   input         cfg_dout106,
   input         cfg_dout107,
   input         cfg_dout108,
   input         cfg_dout109,
   input         cfg_dout110,
   input         cfg_dout111,
   input         cfg_dout112,
   input         cfg_dout113,
   input         cfg_dout114,
   input         cfg_dout115,
   input         cfg_dout116,
   input         cfg_dout117,
   input         cfg_dout118,
   input         cfg_dout119,
   input         cfg_dout120,
   input         cfg_dout121,
   input         cfg_dout122,
   input         cfg_dout123,
   input         cfg_dout124,
   input         cfg_dout125,
   input         cfg_dout126,
   input         cfg_dout127,
   input         cfg_dout128,
   input         cfg_dout129,
   input         cfg_dout130,
   input         cfg_dout131,
   input         cfg_dout132,
   input         cfg_dout133,
   input         cfg_dout134,
   input         cfg_dout135,
   input         cfg_dout136,
   input         cfg_dout137,
   input         cfg_dout138,
   input         cfg_dout139,
   input         cfg_dout140,
   input         cfg_dout141,
   input         cfg_dout142,
   input         cfg_dout143,
   input         cfg_dout144,
   input         cfg_dout145,
   input         cfg_dout146,
   input         cfg_dout147,
   input         cfg_dout148,
   input         cfg_dout149,
   input         cfg_dout150,
   input         cfg_dout151,
   input         cfg_dout152,
   input         cfg_dout153,
   input         cfg_dout154,
   input         cfg_dout155,
   input         cfg_dout156,
   input         cfg_dout157,
   input         cfg_dout158,
   input         cfg_dout159,
   input         cfg_dout160,
   input         cfg_dout161,
   input         cfg_dout162,
   input         cfg_dout163,
   input         cfg_dout164,
   input         cfg_dout165,
   input         cfg_dout166,
   input         cfg_dout167,
   input         cfg_dout168,
   input         cfg_dout169,
   input         cfg_dout170,
   input         cfg_dout171,
   input         cfg_dout172,
   input         cfg_dout173,
   input         cfg_dout174,
   input         cfg_dout175,
   input         cfg_dout176,
   input         cfg_dout177,
   input         cfg_dout178,
   input         cfg_dout179,
   input         cfg_dout180,
   input         cfg_dout181,
   input         cfg_dout182,
   input         cfg_dout183,
   input         cfg_dout184,
   input         cfg_dout185,
   input         cfg_dout186,
   input         cfg_dout187,
   input         cfg_dout188,
   input         cfg_dout189,
   input         cfg_dout190,
   input         cfg_dout191,
   input         cfg_dout192,
   input         cfg_dout193,
   input         cfg_dout194,
   input         cfg_dout195,
   input         cfg_dout196,
   input         cfg_dout197,
   input         cfg_dout198,
   input         cfg_dout199,
   input         cfg_dout200,
   input         cfg_dout201,
   input         cfg_dout202,
   input         cfg_dout203,
   input         cfg_dout204,
   input         cfg_dout205,
   input         cfg_dout206,
   input         cfg_dout207,
   input         cfg_dout208,
   input         cfg_dout209,
   input         cfg_dout210,
   input         cfg_dout211,
   input         cfg_dout212,
   input         cfg_dout213,
   input         cfg_dout214,
   input         cfg_dout215,
   input         cfg_dout216,
   input         cfg_dout217,
   input         cfg_dout218,
   input         cfg_dout219,
   input         cfg_dout220,
   input         cfg_dout221,
   input         cfg_dout222,
   input         cfg_dout223,
   input         cfg_dout224,
   input         cfg_dout225,
   input         cfg_dout226,
   input         cfg_dout227,
   input         cfg_dout228,
   input         cfg_dout229,
   input         cfg_dout230,
   input         cfg_dout231,
   input         cfg_dout232,
   input         cfg_dout233,
   input         cfg_dout234,
   input         cfg_dout235,
   input         cfg_dout236,
   input         cfg_dout237,
   input         cfg_dout238,
   input         cfg_dout239,
   input         cfg_dout240,
   input         cfg_dout241,
   input         cfg_dout242,
   input         cfg_dout243,
   input         cfg_dout244,
   input         cfg_dout245,
   input         cfg_dout246,
   input         cfg_dout247,
   input         cfg_dout248,
   input         cfg_dout249,
   input         cfg_dout250,
   input         cfg_dout251,
   input         cfg_dout252,
   input         cfg_dout253,
   input         cfg_dout254,
   input         cfg_dout255,
   input         cfg_dout256,
   input         cfg_dout257,
   input         cfg_dout258,
   input         cfg_dout259,
   input         cfg_dout260,
   input         cfg_dout261,
   input         cfg_dout262,
   input         cfg_dout263,
   input         cfg_dout264,
   input         cfg_dout265,
   input         cfg_dout266,
   input         cfg_dout267,
   input         cfg_dout268,
   input         cfg_dout269,
   input         cfg_dout270,
   input         cfg_dout271,
   input         cfg_dout272,
   input         cfg_dout273,
   input         cfg_dout274,
   input         cfg_dout275,
   input         cfg_dout276,
   input         cfg_dout277,
   input         cfg_dout278,
   input         cfg_dout279,
   input         cfg_dout280,
   input         cfg_dout281,
   input         cfg_dout282,
   input         cfg_dout283,
   input         cfg_dout284,
   input         cfg_dout285,
   input         cfg_dout286,
   input         cfg_dout287,
   input         cfg_dout288,
   input         cfg_dout289,
   input         cfg_dout290,
   input         cfg_dout291,
   input         cfg_dout292,
   input         cfg_dout293,
   input         cfg_dout294,
   input         cfg_dout295,
   input         cfg_dout296,
   input         cfg_dout297,
   input         cfg_dout298,
   input         cfg_dout299,
   input         cfg_dout300,
   input         cfg_dout301,
   input         cfg_dout302,
   input         cfg_dout303,
   input         cfg_dout304,
   input         cfg_dout305,
   input         cfg_dout306,
   input         cfg_dout307,
   input         cfg_dout308,
   input         cfg_dout309,
   input         cfg_dout310,
   input         cfg_dout311,
   input         cfg_dout312,
   input         cfg_dout313,
   input         cfg_dout314,
   input         cfg_dout315,
   input         cfg_dout316,
   input         cfg_dout317,
   input         cfg_dout318,
   input         cfg_dout319,
   input         cfg_dout320,
   input         cfg_dout321,
   input         cfg_dout322,
   input         cfg_dout323,
   input         cfg_dout324,
   input         cfg_dout325,
   input         cfg_dout326,
   input         cfg_dout327,
   input         cfg_dout328,
   input         cfg_dout329,
   input         cfg_dout330,
   input         cfg_dout331,
   input         cfg_dout332,
   input         cfg_dout333,
   input         cfg_dout334,
   input         cfg_dout335,
   input         cfg_dout336,
   input         cfg_dout337,
   input         cfg_dout338,
   input         cfg_dout339,
   input         cfg_dout340,
   input         cfg_dout341,
   input         cfg_dout342,
   input         cfg_dout343,
   input         cfg_dout344,
   input         cfg_dout345,
   input         cfg_dout346,
   input         cfg_dout347,
   input         cfg_dout348,
   input         cfg_dout349,
   input         cfg_dout350,
   input         cfg_dout351,
   input         cfg_dout352,
   input         cfg_dout353,
   input         cfg_dout354,
   input         cfg_dout355,
   input         cfg_dout356,
   input         cfg_dout357,
   input         cfg_dout358,
   input         cfg_dout359,
   input         cfg_dout360,
   input         cfg_dout361,
   input         cfg_dout362,
   input         cfg_dout363,
   input         cfg_dout364,
   input         cfg_dout365,
   input         cfg_dout366,
   input         cfg_dout367,
   input         cfg_dout368,
   input         cfg_dout369,
   input         cfg_dout370,
   input         cfg_dout371,
   input         cfg_dout372,
   input         cfg_dout373,
   input         cfg_dout374,
   input         cfg_dout375,
   input         cfg_dout376,
   input         cfg_dout377,
   input         cfg_dout378,
   input         cfg_dout379,
   input         cfg_dout380,
   input         cfg_dout381,
   input         cfg_dout382,
   input         cfg_dout383,
   input         cfg_dout384,
   input         cfg_dout385,
   input         cfg_dout386,
   input         cfg_dout387,
   input         cfg_dout388,
   input         cfg_dout389,
   input         cfg_dout390,
   input         cfg_dout391,
   input         cfg_dout392,
   input         cfg_dout393,
   input         cfg_dout394,
   input         cfg_dout395,
   input         cfg_dout396,
   input         cfg_dout397,
   input         cfg_dout398,
   input         cfg_dout399,
   input         cfg_dout400,
   input         cfg_dout401,
   input         cfg_dout402,
   input         cfg_dout403,
   input         cfg_dout404,
   input         cfg_dout405,
   input         cfg_dout406,
   input         cfg_dout407,
   input         cfg_dout408,
   input         cfg_dout409,
   input         cfg_dout410,
   input         cfg_dout411,
   input         cfg_dout412,
   input         cfg_dout413,
   input         cfg_dout414,
   input         cfg_dout415,
   input         cfg_dout416,
   input         cfg_dout417,
   input         cfg_dout418,
   input         cfg_dout419,
   input         cfg_dout420,
   input         cfg_dout421,
   input         cfg_dout422,
   input         cfg_dout423,
   input         cfg_dout424,
   input         cfg_dout425,
   input         cfg_dout426,
   input         cfg_dout427,
   input         cfg_dout428,
   input         cfg_dout429,
   input         cfg_dout430,
   input         cfg_dout431,
   input         cfg_dout432,
   input         cfg_dout433,
   input         cfg_dout434,
   input         cfg_dout435,
   input         cfg_dout436,
   input         cfg_dout437,
   input         cfg_dout438,
   input         cfg_dout439,
   input         cfg_dout440,
   input         cfg_dout441,
   input         cfg_dout442,
   input         cfg_dout443,
   input         cfg_dout444,
   input         cfg_dout445,
   input         cfg_dout446,
   input         cfg_dout447,
   input         cfg_dout448,
   input         cfg_dout449,
   input         cfg_dout450,
   input         cfg_dout451,
   input         cfg_dout452,
   input         cfg_dout453,
   input         cfg_dout454,
   input         cfg_dout455,
   input         cfg_dout456,
   input         cfg_dout457,
   input         cfg_dout458,
   input         cfg_dout459,
   input         cfg_dout460,
   input         cfg_dout461,
   input         cfg_dout462,
   input         cfg_dout463,
   input         cfg_dout464,
   input         cfg_dout465,
   input         cfg_dout466,
   input         cfg_dout467,
   input         cfg_dout468,
   input         cfg_dout469,
   input         cfg_dout470,
   input         cfg_dout471,
   input         cfg_dout472,
   input         cfg_dout473,
   input         cfg_dout474,
   input         cfg_dout475,
   input         cfg_dout476,
   input         cfg_dout477,
   input         cfg_dout478,
   input         cfg_dout479,
   input         cfg_dout480,
   input         cfg_dout481,
   input         cfg_dout482,
   input         cfg_dout483,
   input         cfg_dout484,
   input         cfg_dout485,
   input         cfg_dout486,
   input         cfg_dout487,
   input         cfg_dout488,
   input         cfg_dout489,
   input         cfg_dout490,
   input         cfg_dout491,
   input         cfg_dout492,
   input         cfg_dout493,
   input         cfg_dout494,
   input         cfg_dout495,
   input         cfg_dout496,
   input         cfg_dout497,
   input         cfg_dout498,
   input         cfg_dout499,
   input         cfg_dout500,
   input         cfg_dout501,
   input         cfg_dout502,
   input         cfg_dout503,
   input         cfg_dout504,
   input         cfg_dout505,
   input         cfg_dout506,
   input         cfg_dout507,
   input         cfg_dout508,
   input         cfg_dout509,
   input         cfg_dout510,
   input         cfg_dout511,
   input         cfg_dout512,
   input         cfg_dout513,
   input         cfg_dout514,
   input         cfg_dout515,
   input         cfg_dout516,
   input         cfg_dout517,
   input         cfg_dout518,
   input         cfg_dout519,
   input         cfg_dout520,
   input         cfg_dout521,
   input         cfg_dout522,
   input         cfg_dout523,
   input         cfg_dout524,
   input         cfg_dout525,
   input         cfg_dout526,
   input         cfg_dout527,
   input         cfg_dout528,
   input         cfg_dout529,
   input         cfg_dout530,
   input         cfg_dout531,
   input         cfg_dout532,
   input         cfg_dout533,
   input         cfg_dout534,
   input         cfg_dout535,
   input         cfg_dout536,
   input         cfg_dout537,
   input         cfg_dout538,
   input         cfg_dout539,
   input         cfg_dout540,
   input         cfg_dout541,
   input         cfg_dout542,
   input         cfg_dout543,
   input         cfg_dout544,
   input         cfg_dout545,
   input         cfg_dout546,
   input         cfg_dout547,
   input         cfg_dout548,
   input         cfg_dout549,
   input         cfg_dout550,
   input         cfg_dout551,
   input         cfg_dout552,
   input         cfg_dout553,
   input         cfg_dout554,
   input         cfg_dout555,
   input         cfg_dout556,
   input         cfg_dout557,
   input         cfg_dout558,
   input         cfg_dout559,
   input         cfg_dout560,
   input         cfg_dout561,
   input         cfg_dout562,
   input         cfg_dout563,
   input         cfg_dout564,
   input         cfg_dout565,
   input         cfg_dout566,
   input         cfg_dout567,
   input         cfg_dout568,
   input         cfg_dout569,
   input         cfg_dout570,
   input         cfg_dout571,
   input         cfg_dout572,
   input         cfg_dout573,
   input         cfg_dout574,
   input         cfg_dout575,
   input         cfg_dout576,
   input         cfg_dout577,
   input         cfg_dout578,
   input         cfg_dout579,
   input         cfg_dout580,
   input         cfg_dout581,
   input         cfg_dout582,
   input         cfg_dout583,
   input         cfg_dout584,
   input         cfg_dout585,
   input         cfg_dout586,
   input         cfg_dout587,
   input         cfg_dout588,
   input         cfg_dout589,
   input         cfg_dout590,
   input         cfg_dout591,
   input         cfg_dout592,
   input         cfg_dout593,
   input         cfg_dout594,
   input         cfg_dout595,
   input         cfg_dout596,
   input         cfg_dout597,
   input         cfg_dout598,
   input         cfg_dout599,
   input         cfg_dout600,
   input         cfg_dout601,
   input         cfg_dout602,
   input         cfg_dout603,
   input         cfg_dout604,
   input         cfg_dout605,
   input         cfg_dout606,
   input         cfg_dout607,
   input         cfg_dout608,
   input         cfg_dout609,
   input         cfg_dout610,
   input         cfg_dout611,
   input         cfg_dout612,
   input         cfg_dout613,
   input         cfg_dout614,
   input         cfg_dout615,
   input         cfg_dout616,
   input         cfg_dout617,
   input         cfg_dout618,
   input         cfg_dout619,
   input         cfg_dout620,
   input         cfg_dout621,
   input         cfg_dout622,
   input         cfg_dout623,
   input         cfg_dout624,
   input         cfg_dout625,
   input         cfg_dout626,
   input         cfg_dout627,
   input         cfg_dout628,
   input         cfg_dout629,
   input         cfg_dout630,
   input         cfg_dout631,
   input         cfg_dout632,
   input         cfg_dout633,
   input         cfg_dout634,
   input         cfg_dout635,
   input         cfg_dout636,
   input         cfg_dout637,
   input         cfg_dout638,
   input         cfg_dout639,
   input         cfg_dout640,
   input         cfg_dout641,
   input         cfg_dout642,
   input         cfg_dout643,
   input         cfg_dout644,
   input         cfg_dout645,
   input         cfg_dout646,
   input         cfg_dout647,
   input         cfg_dout648,
   input         cfg_dout649,
   input         cfg_dout650,
   input         cfg_dout651,
   input         cfg_dout652,
   input         cfg_dout653,
   input         cfg_dout654,
   input         cfg_dout655,
   input         cfg_dout656,
   input         cfg_dout657,
   input         cfg_dout658,
   input         cfg_dout659,
   input         cfg_dout660,
   input         cfg_dout661,
   input         cfg_dout662,
   input         cfg_dout663,
   input         cfg_dout664,
   input         cfg_dout665,
   input         cfg_dout666,
   input         cfg_dout667,
   input         cfg_dout668,
   input         cfg_dout669,
   input         cfg_dout670,
   input         cfg_dout671,
   input         cfg_dout672,
   input         cfg_dout673,
   input         cfg_dout674,
   input         cfg_dout675,
   input         cfg_dout676,
   input         cfg_dout677,
   input         cfg_dout678,
   input         cfg_dout679,
   input         cfg_dout680,
   input         cfg_dout681,
   input         cfg_dout682,
   input         cfg_dout683,
   input         cfg_dout684,
   input         cfg_dout685,
   input         cfg_dout686,
   input         cfg_dout687,
   input         cfg_dout688,
   input         cfg_dout689,
   input         cfg_dout690,
   input         cfg_dout691,
   input         cfg_dout692,
   input         cfg_dout693,
   input         cfg_dout694,
   input         cfg_dout695,
   input         cfg_dout696,
   input         cfg_dout697,
   input         cfg_dout698,
   input         cfg_dout699,
   input         cfg_dout700,
   input         cfg_dout701,
   input         cfg_dout702,
   input         cfg_dout703,
   input         cfg_dout704,
   input         cfg_dout705,
   input         cfg_dout706,
   input         cfg_dout707,
   input         cfg_dout708,
   input         cfg_dout709,
   input         cfg_dout710,
   input         cfg_dout711,
   input         cfg_dout712,
   input         cfg_dout713,
   input         cfg_dout714,
   input         cfg_dout715,
   input         cfg_dout716,
   input         cfg_dout717,
   input         cfg_dout718,
   input         cfg_dout719,
   input         cfg_dout720,
   input         cfg_dout721,
   input         cfg_dout722,
   input         cfg_dout723,
   input         cfg_dout724,
   input         cfg_dout725,
   input         cfg_dout726,
   input         cfg_dout727,
   input         cfg_dout728,
   input         cfg_dout729,
   input         cfg_dout730,
   input         cfg_dout731,
   input         cfg_dout732,
   input         cfg_dout733,
   input         cfg_dout734,
   input         cfg_dout735,
   input         cfg_dout736,
   input         cfg_dout737,
   input         cfg_dout738,
   input         cfg_dout739,
   input         cfg_dout740,
   input         cfg_dout741,
   input         cfg_dout742,
   input         cfg_dout743,
   input         cfg_dout744,
   input         cfg_dout745,
   input         cfg_dout746,
   input         cfg_dout747,
   input         cfg_dout748,
   input         cfg_dout749,
   input         cfg_dout750,
   input         cfg_dout751,
   input         cfg_dout752,
   input         cfg_dout753,
   input         cfg_dout754,
   input         cfg_dout755,
   input         cfg_dout756,
   input         cfg_dout757,
   input         cfg_dout758,
   input         cfg_dout759,
   input         cfg_dout760,
   input         cfg_dout761,
   input         cfg_dout762,
   input         cfg_dout763,
   input         cfg_dout764,
   input         cfg_dout765,
   input         cfg_dout766,
   input         cfg_dout767,
   input         cfg_dout768,
   input         cfg_dout769,
   input         cfg_dout770,
   input         cfg_dout771,
   input         cfg_dout772,
   input         cfg_dout773,
   input         cfg_dout774,
   input         cfg_dout775,
   input         cfg_dout776,
   input         cfg_dout777,
   input         cfg_dout778,
   input         cfg_dout779,
   input         cfg_dout780,
   input         cfg_dout781,
   input         cfg_dout782,
   input         cfg_dout783,
   input         cfg_dout784,
   input         cfg_dout785,
   input         cfg_dout786,
   input         cfg_dout787,
   input         cfg_dout788,
   input         cfg_dout789,
   input         cfg_dout790,
   input         cfg_dout791,
   input         cfg_dout792,
   input         cfg_dout793,
   input         cfg_dout794,
   input         cfg_dout795,
   input         cfg_dout796,
   input         cfg_dout797,
   input         cfg_dout798,
   input         cfg_dout799,
   input         cfg_dout800,
   input         cfg_dout801,
   input         cfg_dout802,
   input         cfg_dout803,
   input         cfg_dout804,
   input         cfg_dout805,
   input         cfg_dout806,
   input         cfg_dout807,
   input         cfg_dout808,
   input         cfg_dout809,
   input         cfg_dout810,
   input         cfg_dout811,
   input         cfg_dout812,
   input         cfg_dout813,
   input         cfg_dout814,
   input         cfg_dout815,
   input         cfg_dout816,
   input         cfg_dout817,
   input         cfg_dout818,
   input         cfg_dout819,
   input         cfg_dout820,
   input         cfg_dout821,
   input         cfg_dout822,
   input         cfg_dout823,
   input         cfg_dout824,
   input         cfg_dout825,
   input         cfg_dout826,
   input         cfg_dout827,
   input         cfg_dout828,
   input         cfg_dout829,
   input         cfg_dout830,
   input         cfg_dout831,
   input         cfg_dout832,
   input         cfg_dout833,
   input         cfg_dout834,
   input         cfg_dout835,
   input         cfg_dout836,
   input         cfg_dout837,
   input         cfg_dout838,
   input         cfg_dout839,
   input         cfg_dout840,
   input         cfg_dout841,
   input         cfg_dout842,
   input         cfg_dout843,
   input         cfg_dout844,
   input         cfg_dout845,
   input         cfg_dout846,
   input         cfg_dout847,
   input         cfg_dout848,
   input         cfg_dout849,
   input         cfg_dout850,
   input         cfg_dout851,
   input         cfg_dout852,
   input         cfg_dout853,
   input         cfg_dout854,
   input         cfg_dout855,
   input         cfg_dout856,
   input         cfg_dout857,
   input         cfg_dout858,
   input         cfg_dout859,
   input         cfg_dout860,
   input         cfg_dout861,
   input         cfg_dout862,
   input         cfg_dout863,
   input         cfg_dout864,
   input         cfg_dout865,
   input         cfg_dout866,
   input         cfg_dout867,
   input         cfg_dout868,
   input         cfg_dout869,
   input         cfg_dout870,
   input         cfg_dout871,
   input         cfg_dout872,
   input         cfg_dout873,
   input         cfg_dout874,
   input         cfg_dout875,
   input         cfg_dout876,
   input         cfg_dout877,
   input         cfg_dout878,
   input         cfg_dout879,
   input         cfg_dout880,
   input         cfg_dout881,
   input         cfg_dout882,
   input         cfg_dout883,
   input         cfg_dout884,
   input         cfg_dout885,
   input         cfg_dout886,
   input         cfg_dout887,
   input         cfg_dout888,
   input         cfg_dout889,
   input         cfg_dout890,
   input         cfg_dout891,
   input         cfg_dout892,
   input         cfg_dout893,
   input         cfg_dout894,
   input         cfg_dout895,
   input         cfg_dout896,
   input         cfg_dout897,
   input         cfg_dout898,
   input         cfg_dout899,
   input         cfg_dout900,
   input         cfg_dout901,
   input         cfg_dout902,
   input         cfg_dout903,
   input         cfg_dout904,
   input         cfg_dout905,
   input         cfg_dout906,
   input         cfg_dout907,
   input         cfg_dout908,
   input         cfg_dout909,
   input         cfg_dout910,
   input         cfg_dout911,
   input         cfg_dout912,
   input         cfg_dout913,
   input         cfg_dout914,
   input         cfg_dout915,
   input         cfg_dout916,
   input         cfg_dout917,
   input         cfg_dout918,
   input         cfg_dout919,
   input         cfg_dout920,
   input         cfg_dout921,
   input         cfg_dout922,
   input         cfg_dout923,
   input         cfg_dout924,
   input         cfg_dout925,
   input         cfg_dout926,
   input         cfg_dout927,
   input         cfg_dout928,
   input         cfg_dout929,
   input         cfg_dout930,
   input         cfg_dout931,
   input         cfg_dout932,
   input         cfg_dout933,
   input         cfg_dout934,
   input         cfg_dout935,
   input         cfg_dout936,
   input         cfg_dout937,
   input         cfg_dout938,
   input         cfg_dout939,
   input         cfg_dout940,
   input         cfg_dout941,
   input         cfg_dout942,
   input         cfg_dout943,
   input         cfg_dout944,
   input         cfg_dout945,
   input         cfg_dout946,
   input         cfg_dout947,
   input         cfg_dout948,
   input         cfg_dout949,
   input         cfg_dout950,
   input         cfg_dout951,
   input         cfg_dout952,
   input         cfg_dout953,
   input         cfg_dout954,
   input         cfg_dout955,
   input         cfg_dout956,
   input         cfg_dout957,
   input         cfg_dout958,
   input         cfg_dout959,
   input         cfg_dout960,
   input         cfg_dout961,
   input         cfg_dout962,
   input         cfg_dout963,
   input         cfg_dout964,
   input         cfg_dout965,
   input         cfg_dout966,
   input         cfg_dout967,
   input         cfg_dout968,
   input         cfg_dout969,
   input         cfg_dout970,
   input         cfg_dout971,
   input         cfg_dout972,
   input         cfg_dout973,
   input         cfg_dout974,
   input         cfg_dout975,
   input         cfg_dout976,
   input         cfg_dout977,
   input         cfg_dout978,
   input         cfg_dout979,
   input         cfg_dout980,
   input         cfg_dout981,
   input         cfg_dout982,
   input         cfg_dout983,
   input         cfg_dout984,
   input         cfg_dout985,
   input         cfg_dout986,
   input         cfg_dout987,
   input         cfg_dout988,
   input         cfg_dout989,
   input         cfg_dout990,
   input         cfg_dout991,
   input         cfg_dout992,
   input         cfg_dout993,
   input         cfg_dout994,
   input         cfg_dout995,
   input         cfg_dout996,
   input         cfg_dout997,
   input         cfg_dout998,
   input         cfg_dout999,
   input         cfg_dout1000,
   input         cfg_dout1001,
   input         cfg_dout1002,
   input         cfg_dout1003,
   input         cfg_dout1004,
   input         cfg_dout1005,
   input         cfg_dout1006,
   input         cfg_dout1007,
   input         cfg_dout1008,
   input         cfg_dout1009,
   input         cfg_dout1010,
   input         cfg_dout1011,
   input         cfg_dout1012,
   input         cfg_dout1013,
   input         cfg_dout1014,
   input         cfg_dout1015,
   input         cfg_dout1016,
   input         cfg_dout1017,
   input         cfg_dout1018,
   input         cfg_dout1019,
   input         cfg_dout1020,
   input         cfg_dout1021,
   input         cfg_dout1022,
   input         cfg_dout1023,
   input         cfg_dout1024,
   input         cfg_dout1025,
   input         cfg_dout1026,
   input         cfg_dout1027,
   input         cfg_dout1028,
   input         cfg_dout1029,
   input         cfg_dout1030,
   input         cfg_dout1031,
   input         cfg_dout1032,
   input         cfg_dout1033,
   input         cfg_dout1034,
   input         cfg_dout1035,
   input         cfg_dout1036,
   input         cfg_dout1037,
   input         cfg_dout1038,
   input         cfg_dout1039,
   input         cfg_dout1040,
   input         cfg_dout1041,
   input         cfg_dout1042,
   input         cfg_dout1043,
   input         cfg_dout1044,
   input         cfg_dout1045,
   input         cfg_dout1046,
   input         cfg_dout1047,
   input         cfg_dout1048,
   input         cfg_dout1049,
   input         cfg_dout1050,
   input         cfg_dout1051,
   input         cfg_dout1052,
   input         cfg_dout1053,
   input         cfg_dout1054,
   input         cfg_dout1055,
   input         cfg_dout1056,
   input         cfg_dout1057,
   input         cfg_dout1058,
   input         cfg_dout1059,
   input         cfg_dout1060,
   input         cfg_dout1061,
   input         cfg_dout1062,
   input         cfg_dout1063,
   input         cfg_dout1064,
   input         cfg_dout1065,
   input         cfg_dout1066,
   input         cfg_dout1067,
   input         cfg_dout1068,
   input         cfg_dout1069,
   input         cfg_dout1070,
   input         cfg_dout1071,
   input         cfg_dout1072,
   input         cfg_dout1073,
   input         cfg_dout1074,
   input         cfg_dout1075,
   input         cfg_dout1076,
   input         cfg_dout1077,
   input         cfg_dout1078,
   input         cfg_dout1079,
   input         cfg_dout1080,
   input         cfg_dout1081,
   input         cfg_dout1082,
   input         cfg_dout1083,
   input         cfg_dout1084,
   input         cfg_dout1085,
   input         cfg_dout1086,
   input         cfg_dout1087,
   input         cfg_dout1088,
   input         cfg_dout1089,
   input         cfg_dout1090,
   input         cfg_dout1091,
   input         cfg_dout1092,
   input         cfg_dout1093,
   input         cfg_dout1094,
   input         cfg_dout1095,
   input         cfg_dout1096,
   input         cfg_dout1097,
   input         cfg_dout1098,
   input         cfg_dout1099,
   input         cfg_dout1100,
   input         cfg_dout1101,
   input         cfg_dout1102,
   input         cfg_dout1103,
   input         cfg_dout1104,
   input         cfg_dout1105,
   input         cfg_dout1106,
   input         cfg_dout1107,
   input         cfg_dout1108,
   input         cfg_dout1109,
   input         cfg_dout1110,
   input         cfg_dout1111,
   input         cfg_dout1112,
   input         cfg_dout1113,
   input         cfg_dout1114,
   input         cfg_dout1115,
   input         cfg_dout1116,
   input         cfg_dout1117,
   input         cfg_dout1118,
   input         cfg_dout1119,
   input         cfg_dout1120,
   input         cfg_dout1121,
   input         cfg_dout1122,
   input         cfg_dout1123,
   input         cfg_dout1124,
   input         cfg_dout1125,
   input         cfg_dout1126,
   input         cfg_dout1127,
   input         cfg_dout1128,
   input         cfg_dout1129,
   input         cfg_dout1130,
   input         cfg_dout1131,
   input         cfg_dout1132,
   input         cfg_dout1133,
   input         cfg_dout1134,
   input         cfg_dout1135,
   input         cfg_dout1136,
   input         cfg_dout1137,
   input         cfg_dout1138,
   input         cfg_dout1139,
   input         cfg_dout1140,
   input         cfg_dout1141,
   input         cfg_dout1142,
   input         cfg_dout1143,
   input         cfg_dout1144,
   input         cfg_dout1145,
   input         cfg_dout1146,
   input         cfg_dout1147,
   input         cfg_dout1148,
   input         cfg_dout1149,
   input         cfg_dout1150,
   input         cfg_dout1151,
   input         cfg_dout1152,
   input         cfg_dout1153,
   input         cfg_dout1154,
   input         cfg_dout1155,
   input         cfg_dout1156,
   input         cfg_dout1157,
   input         cfg_dout1158,
   input         cfg_dout1159,
   input         cfg_dout1160,
   input         cfg_dout1161,
   input         cfg_dout1162,
   input         cfg_dout1163,
   input         cfg_dout1164,
   input         cfg_dout1165,
   input         cfg_dout1166,
   input         cfg_dout1167,
   input         cfg_dout1168,
   input         cfg_dout1169,
   input         cfg_dout1170,
   input         cfg_dout1171,
   input         cfg_dout1172,
   input         cfg_dout1173,
   input         cfg_dout1174,
   input         cfg_dout1175,
   input         cfg_dout1176,
   input         cfg_dout1177,
   input         cfg_dout1178,
   input         cfg_dout1179,
   input         cfg_dout1180,
   input         cfg_dout1181,
   input         cfg_dout1182,
   input         cfg_dout1183,
   input         cfg_dout1184,
   input         cfg_dout1185,
   input         cfg_dout1186,
   input         cfg_dout1187,
   input         cfg_dout1188,
   input         cfg_dout1189,
   input         cfg_dout1190,
   input         cfg_dout1191,
   input         cfg_dout1192,
   input         cfg_dout1193,
   input         cfg_dout1194,
   input         cfg_dout1195,
   input         cfg_dout1196,
   input         cfg_dout1197,
   input         cfg_dout1198,
   input         cfg_dout1199,
   input         cfg_dout1200,
   input         cfg_dout1201,
   input         cfg_dout1202,
   input         cfg_dout1203,
   input         cfg_dout1204,
   input         cfg_dout1205,
   input         cfg_dout1206,
   input         cfg_dout1207,
   input         cfg_dout1208,
   input         cfg_dout1209,
   input         cfg_dout1210,
   input         cfg_dout1211,
   input         cfg_dout1212,
   input         cfg_dout1213,
   input         cfg_dout1214,
   input         cfg_dout1215,
   input         cfg_dout1216,
   input         cfg_dout1217,
   input         cfg_dout1218,
   input         cfg_dout1219,
   input         cfg_dout1220,
   input         cfg_dout1221,
   input         cfg_dout1222,
   input         cfg_dout1223,
   input         cfg_dout1224,
   input         cfg_dout1225,
   input         cfg_dout1226,
   input         cfg_dout1227,
   input         cfg_dout1228,
   input         cfg_dout1229,
   input         cfg_dout1230,
   input         cfg_dout1231,
   input         cfg_dout1232,
   input         cfg_dout1233,
   input         cfg_dout1234,
   input         cfg_dout1235,
   input         cfg_dout1236,
   input         cfg_dout1237,
   input         cfg_dout1238,
   input         cfg_dout1239,
   input         cfg_dout1240,
   input         cfg_dout1241,
   input         cfg_dout1242,
   input         cfg_dout1243,
   input         cfg_dout1244,
   input         cfg_dout1245,
   input         cfg_dout1246,
   input         cfg_dout1247,
   input         cfg_dout1248,
   input         cfg_dout1249,
   input         cfg_dout1250,
   input         cfg_dout1251,
   input         cfg_dout1252,
   input         cfg_dout1253,
   input         cfg_dout1254,
   input         cfg_dout1255,
   input         cfg_dout1256,
   input         cfg_dout1257,
   input         cfg_dout1258,
   input         cfg_dout1259,
   input         cfg_dout1260,
   input         cfg_dout1261,
   input         cfg_dout1262,
   input         cfg_dout1263,
   input         cfg_dout1264,
   input         cfg_dout1265,
   input         cfg_dout1266,
   input         cfg_dout1267,
   input         cfg_dout1268,
   input         cfg_dout1269,
   input         cfg_dout1270,
   input         cfg_dout1271,
   input         cfg_dout1272,
   input         cfg_dout1273,
   input         cfg_dout1274,
   input         cfg_dout1275,
   input         cfg_dout1276,
   input         cfg_dout1277,
   input         cfg_dout1278,
   input         cfg_dout1279,
   input         cfg_dout1280,
   input         cfg_dout1281,
   input         cfg_dout1282,
   input         cfg_dout1283,
   input         cfg_dout1284,
   input         cfg_dout1285,
   input         cfg_dout1286,
   input         cfg_dout1287,
   input         cfg_dout1288,
   input         cfg_dout1289,
   input         cfg_dout1290,
   input         cfg_dout1291,
   input         cfg_dout1292,
   input         cfg_dout1293,
   input         cfg_dout1294,
   input         cfg_dout1295,
   input         cfg_dout1296,
   input         cfg_dout1297,
   input         cfg_dout1298,
   input         cfg_dout1299,
   input         cfg_dout1300,
   input         cfg_dout1301,
   input         cfg_dout1302,
   input         cfg_dout1303,
   input         cfg_dout1304,
   input         cfg_dout1305,
   input         cfg_dout1306,
   input         cfg_dout1307,
   input         cfg_dout1308,
   input         cfg_dout1309,
   input         cfg_dout1310,
   input         cfg_dout1311,
   input         cfg_dout1312,
   input         cfg_dout1313,
   input         cfg_dout1314,
   input         cfg_dout1315,
   input         cfg_dout1316,
   input         cfg_dout1317,
   input         cfg_dout1318,
   input         cfg_dout1319,
   input         cfg_dout1320,
   input         cfg_dout1321,
   input         cfg_dout1322,
   input         cfg_dout1323,
   input         cfg_dout1324,
   input         cfg_dout1325,
   input         cfg_dout1326,
   input         cfg_dout1327,
   input         cfg_dout1328,
   input         cfg_dout1329,
   input         cfg_dout1330,
   input         cfg_dout1331,
   input         cfg_dout1332,
   input         cfg_dout1333,
   input         cfg_dout1334,
   input         cfg_dout1335,
   input         cfg_dout1336,
   input         cfg_dout1337,
   input         cfg_dout1338,
   input         cfg_dout1339,
   input         cfg_dout1340,
   input         cfg_dout1341,
   input         cfg_dout1342,
   input         cfg_dout1343,
   input         cfg_dout1344,
   input         cfg_dout1345,
   input         cfg_dout1346,
   input         cfg_dout1347,
   input         cfg_dout1348,
   input         cfg_dout1349,
   input         cfg_dout1350,
   input         cfg_dout1351,
   input         cfg_dout1352,
   input         cfg_dout1353,
   input         cfg_dout1354,
   input         cfg_dout1355,
   input         cfg_dout1356,
   input         cfg_dout1357,
   input         cfg_dout1358,
   input         cfg_dout1359,
   input         cfg_dout1360,
   input         cfg_dout1361,
   input         cfg_dout1362,
   input         cfg_dout1363,
   input         cfg_dout1364,
   input         cfg_dout1365,
   input         cfg_dout1366,
   input         cfg_dout1367,
   input         cfg_dout1368,
   input         cfg_dout1369,
   input         cfg_dout1370,
   input         cfg_dout1371,
   input         cfg_dout1372,
   input         cfg_dout1373,
   input         cfg_dout1374,
   input         cfg_dout1375,
   input         cfg_dout1376,
   input         cfg_dout1377,
   input         cfg_dout1378,
   input         cfg_dout1379,
   input         cfg_dout1380,
   input         cfg_dout1381,
   input         cfg_dout1382,
   input         cfg_dout1383,
   input         cfg_dout1384,
   input         cfg_dout1385,
   input         cfg_dout1386,
   input         cfg_dout1387,
   input         cfg_dout1388,
   input         cfg_dout1389,
   input         cfg_dout1390,
   input         cfg_dout1391,
   input         cfg_dout1392,
   input         cfg_dout1393,
   input         cfg_dout1394,
   input         cfg_dout1395,
   input         cfg_dout1396,
   input         cfg_dout1397,
   input         cfg_dout1398,
   input         cfg_dout1399,
   input         cfg_dout1400,
   input         cfg_dout1401,
   input         cfg_dout1402,
   input         cfg_dout1403,
   input         cfg_dout1404,
   input         cfg_dout1405,
   input         cfg_dout1406,
   input         cfg_dout1407,
   input         cfg_dout1408,
   input         cfg_dout1409,
   input         cfg_dout1410,
   input         cfg_dout1411,
   input         cfg_dout1412,
   input         cfg_dout1413,
   input         cfg_dout1414,
   input         cfg_dout1415,
   input         cfg_dout1416,
   input         cfg_dout1417,
   input         cfg_dout1418,
   input         cfg_dout1419,
   input         cfg_dout1420,
   input         cfg_dout1421,
   input         cfg_dout1422,
   input         cfg_dout1423,
   input         cfg_dout1424,
   input         cfg_dout1425,
   input         cfg_dout1426,
   input         cfg_dout1427,
   input         cfg_dout1428,
   input         cfg_dout1429,
   input         cfg_dout1430,
   input         cfg_dout1431,
   input         cfg_dout1432,
   input         cfg_dout1433,
   input         cfg_dout1434,
   input         cfg_dout1435,
   input         cfg_dout1436,
   input         cfg_dout1437,
   input         cfg_dout1438,
   input         cfg_dout1439,
   input         cfg_dout1440,
   input         cfg_dout1441,
   input         cfg_dout1442,
   input         cfg_dout1443,
   input         cfg_dout1444,
   input         cfg_dout1445,
   input         cfg_dout1446,
   input         cfg_dout1447,
   input         cfg_dout1448,
   input         cfg_dout1449,
   input         cfg_dout1450,
   input         cfg_dout1451,
   input         cfg_dout1452,
   input         cfg_dout1453,
   input         cfg_dout1454,
   input         cfg_dout1455,
   input         cfg_dout1456,
   input         cfg_dout1457,
   input         cfg_dout1458,
   input         cfg_dout1459,
   input         cfg_dout1460,
   input         cfg_dout1461,
   input         cfg_dout1462,
   input         cfg_dout1463,
   input         cfg_dout1464,
   input         cfg_dout1465,
   input         cfg_dout1466,
   input         cfg_dout1467,
   input         cfg_dout1468,
   input         cfg_dout1469,
   input         cfg_dout1470,
   input         cfg_dout1471,
   input         cfg_dout1472,
   input         cfg_dout1473,
   input         cfg_dout1474,
   input         cfg_dout1475,
   input         cfg_dout1476,
   input         cfg_dout1477,
   input         cfg_dout1478,
   input         cfg_dout1479,
   input         cfg_dout1480,
   input         cfg_dout1481,
   input         cfg_dout1482,
   input         cfg_dout1483,
   input         cfg_dout1484,
   input         cfg_dout1485,
   input         cfg_dout1486,
   input         cfg_dout1487,
   input         cfg_dout1488,
   input         cfg_dout1489,
   input         cfg_dout1490,
   input         cfg_dout1491,
   input         cfg_dout1492,
   input         cfg_dout1493,
   input         cfg_dout1494,
   input         cfg_dout1495,
   input         cfg_dout1496,
   input         cfg_dout1497,
   input         cfg_dout1498,
   input         cfg_dout1499,
   input         cfg_dout1500,
   input         cfg_dout1501,
   input         cfg_dout1502,
   input         cfg_dout1503,
   input         cfg_dout1504,
   input         cfg_dout1505,
   input         cfg_dout1506,
   input         cfg_dout1507,
   input         cfg_dout1508,
   input         cfg_dout1509,
   input         cfg_dout1510,
   input         cfg_dout1511,
   input         cfg_dout1512,
   input         cfg_dout1513,
   input         cfg_dout1514,
   input         cfg_dout1515,
   input         cfg_dout1516,
   input         cfg_dout1517,
   input         cfg_dout1518,
   input         cfg_dout1519,
   input         cfg_dout1520,
   input         cfg_dout1521,
   input         cfg_dout1522,
   input         cfg_dout1523,
   input         cfg_dout1524,
   input         cfg_dout1525,
   input         cfg_dout1526,
   input         cfg_dout1527,
   input         cfg_dout1528,
   input         cfg_dout1529,
   input         cfg_dout1530,
   input         cfg_dout1531,
   input         cfg_dout1532,
   input         cfg_dout1533,
   input         cfg_dout1534,
   input         cfg_dout1535,
   input         cfg_dout1536,
   input         cfg_dout1537,
   input         cfg_dout1538,
   input         cfg_dout1539,
   input         cfg_dout1540,
   input         cfg_dout1541,
   input         cfg_dout1542,
   input         cfg_dout1543,
   input         cfg_dout1544,
   input         cfg_dout1545,
   input         cfg_dout1546,
   input         cfg_dout1547,
   input         cfg_dout1548,
   input         cfg_dout1549,
   input         cfg_dout1550,
   input         cfg_dout1551,
   input         cfg_dout1552,
   input         cfg_dout1553,
   input         cfg_dout1554,
   input         cfg_dout1555,
   input         cfg_dout1556,
   input         cfg_dout1557,
   input         cfg_dout1558,
   input         cfg_dout1559,
   input         cfg_dout1560,
   input         cfg_dout1561,
   input         cfg_dout1562,
   input         cfg_dout1563,
   input         cfg_dout1564,
   input         cfg_dout1565,
   input         cfg_dout1566,
   input         cfg_dout1567,
   input         cfg_dout1568,
   input         cfg_dout1569,
   input         cfg_dout1570,
   input         cfg_dout1571,
   input         cfg_dout1572,
   input         cfg_dout1573,
   input         cfg_dout1574,
   input         cfg_dout1575,
   input         cfg_dout1576,
   input         cfg_dout1577,
   input         cfg_dout1578,
   input         cfg_dout1579,
   input         cfg_dout1580,
   input         cfg_dout1581,
   input         cfg_dout1582,
   input         cfg_dout1583,
   input         cfg_dout1584,
   input         cfg_dout1585,
   input         cfg_dout1586,
   input         cfg_dout1587,
   input         cfg_dout1588,
   input         cfg_dout1589,
   input         cfg_dout1590,
   input         cfg_dout1591,
   input         cfg_dout1592,
   input         cfg_dout1593,
   input         cfg_dout1594,
   input         cfg_dout1595,
   input         cfg_dout1596,
   input         cfg_dout1597,
   input         cfg_dout1598,
   input         cfg_dout1599,
   input         cfg_dout1600,
   input         cfg_dout1601,
   input         cfg_dout1602,
   input         cfg_dout1603,
   input         cfg_dout1604,
   input         cfg_dout1605,
   input         cfg_dout1606,
   input         cfg_dout1607,
   input         cfg_dout1608,
   input         cfg_dout1609,
   input         cfg_dout1610,
   input         cfg_dout1611,
   input         cfg_dout1612,
   input         cfg_dout1613,
   input         cfg_dout1614,
   input         cfg_dout1615,
   input         cfg_dout1616,
   input         cfg_dout1617,
   input         cfg_dout1618,
   input         cfg_dout1619,
   input         cfg_dout1620,
   input         cfg_dout1621,
   input         cfg_dout1622,
   input         cfg_dout1623,
   input         cfg_dout1624,
   input         cfg_dout1625,
   input         cfg_dout1626,
   input         cfg_dout1627,
   input         cfg_dout1628,
   input         cfg_dout1629,
   input         cfg_dout1630,
   input         cfg_dout1631,
   input         cfg_dout1632,
   input         cfg_dout1633,
   input         cfg_dout1634,
   input         cfg_dout1635,
   input         cfg_dout1636,
   input         cfg_dout1637,
   input         cfg_dout1638,
   input         cfg_dout1639,
   input         cfg_dout1640,
   input         cfg_dout1641,
   input         cfg_dout1642,
   input         cfg_dout1643,
   input         cfg_dout1644,
   input         cfg_dout1645,
   input         cfg_dout1646,
   input         cfg_dout1647,
   input         cfg_dout1648,
   input         cfg_dout1649,
   input         cfg_dout1650,
   input         cfg_dout1651,
   input         cfg_dout1652,
   input         cfg_dout1653,
   input         cfg_dout1654,
   input         cfg_dout1655,
   input         cfg_dout1656,
   input         cfg_dout1657,
   input         cfg_dout1658,
   input         cfg_dout1659,
   input         cfg_dout1660,
   input         cfg_dout1661,
   input         cfg_dout1662,
   input         cfg_dout1663,
   input         cfg_dout1664,
   input         cfg_dout1665,
   input         cfg_dout1666,
   input         cfg_dout1667,
   input         cfg_dout1668,
   input         cfg_dout1669,
   input         cfg_dout1670,
   input         cfg_dout1671,
   input         cfg_dout1672,
   input         cfg_dout1673,
   input         cfg_dout1674,
   input         cfg_dout1675,
   input         cfg_dout1676,
   input         cfg_dout1677,
   input         cfg_dout1678,
   input         cfg_dout1679,
   input         cfg_dout1680,
   input         cfg_dout1681,
   input         cfg_dout1682,
   input         cfg_dout1683,
   input         cfg_dout1684,
   input         cfg_dout1685,
   input         cfg_dout1686,
   input         cfg_dout1687,
   input         cfg_dout1688,
   input         cfg_dout1689,
   input         cfg_dout1690,
   input         cfg_dout1691,
   input         cfg_dout1692,
   input         cfg_dout1693,
   input         cfg_dout1694,
   input         cfg_dout1695,
   input         cfg_dout1696,
   input         cfg_dout1697,
   input         cfg_dout1698,
   input         cfg_dout1699,
   input         cfg_dout1700,
   input         cfg_dout1701,
   input         cfg_dout1702,
   input         cfg_dout1703,
   input         cfg_dout1704,
   input         cfg_dout1705,
   input         cfg_dout1706,
   input         cfg_dout1707,
   input         cfg_dout1708,
   input         cfg_dout1709,
   input         cfg_dout1710,
   input         cfg_dout1711,
   input         cfg_dout1712,
   input         cfg_dout1713,
   input         cfg_dout1714,
   input         cfg_dout1715,
   input         cfg_dout1716,
   input         cfg_dout1717,
   input         cfg_dout1718,
   input         cfg_dout1719,
   input         cfg_dout1720,
   input         cfg_dout1721,
   input         cfg_dout1722,
   input         cfg_dout1723,
   input         cfg_dout1724,
   input         cfg_dout1725,
   input         cfg_dout1726,
   input         cfg_dout1727,
   input         cfg_dout1728,
   input         cfg_dout1729,
   input         cfg_dout1730,
   input         cfg_dout1731,
   input         cfg_dout1732,
   input         cfg_dout1733,
   input         cfg_dout1734,
   input         cfg_dout1735,
   input         cfg_dout1736,
   input         cfg_dout1737,
   input         cfg_dout1738,
   input         cfg_dout1739,
   input         cfg_dout1740,
   input         cfg_dout1741,
   input         cfg_dout1742,
   input         cfg_dout1743,
   input         cfg_dout1744,
   input         cfg_dout1745,
   input         cfg_dout1746,
   input         cfg_dout1747,
   input         cfg_dout1748,
   input         cfg_dout1749,
   input         cfg_dout1750,
   input         cfg_dout1751,
   input         cfg_dout1752,
   input         cfg_dout1753,
   input         cfg_dout1754,
   input         cfg_dout1755,
   input         cfg_dout1756,
   input         cfg_dout1757,
   input         cfg_dout1758,
   input         cfg_dout1759,
   input         cfg_dout1760,
   input         cfg_dout1761,
   input         cfg_dout1762,
   input         cfg_dout1763,
   input         cfg_dout1764,
   input         cfg_dout1765,
   input         cfg_dout1766,
   input         cfg_dout1767,
   input         cfg_dout1768,
   input         cfg_dout1769,
   input         cfg_dout1770,
   input         cfg_dout1771,
   input         cfg_dout1772,
   input         cfg_dout1773,
   input         cfg_dout1774,
   input         cfg_dout1775,
   input         cfg_dout1776,
   input         cfg_dout1777,
   input         cfg_dout1778,
   input         cfg_dout1779,
   input         cfg_dout1780,
   input         cfg_dout1781,
   input         cfg_dout1782,
   input         cfg_dout1783,
   input         cfg_dout1784,
   input         cfg_dout1785,
   input         cfg_dout1786,
   input         cfg_dout1787,
   input         cfg_dout1788,
   input         cfg_dout1789,
   input         cfg_dout1790,
   input         cfg_dout1791,
   input         cfg_dout1792,
   input         cfg_dout1793,
   input         cfg_dout1794,
   input         cfg_dout1795,
   input         cfg_dout1796,
   input         cfg_dout1797,
   input         cfg_dout1798,
   input         cfg_dout1799,
   input         cfg_dout1800,
   input         cfg_dout1801,
   input         cfg_dout1802,
   input         cfg_dout1803,
   input         cfg_dout1804,
   input         cfg_dout1805,
   input         cfg_dout1806,
   input         cfg_dout1807,
   input         cfg_dout1808,
   input         cfg_dout1809,
   input         cfg_dout1810,
   input         cfg_dout1811,
   input         cfg_dout1812,
   input         cfg_dout1813,
   input         cfg_dout1814,
   input         cfg_dout1815,
   input         cfg_dout1816,
   input         cfg_dout1817,
   input         cfg_dout1818,
   input         cfg_dout1819,
   input         cfg_dout1820,
   input         cfg_dout1821,
   input         cfg_dout1822,
   input         cfg_dout1823,
   input         cfg_dout1824,
   input         cfg_dout1825,
   input         cfg_dout1826,
   input         cfg_dout1827,
   input         cfg_dout1828,
   input         cfg_dout1829,
   input         cfg_dout1830,
   input         cfg_dout1831,
   input         cfg_dout1832,
   input         cfg_dout1833,
   input         cfg_dout1834,
   input         cfg_dout1835,
   input         cfg_dout1836,
   input         cfg_dout1837,
   input         cfg_dout1838,
   input         cfg_dout1839,
   input         cfg_dout1840,
   input         cfg_dout1841,
   input         cfg_dout1842,
   input         cfg_dout1843,
   input         cfg_dout1844,
   input         cfg_dout1845,
   input         cfg_dout1846,
   input         cfg_dout1847,
   input         cfg_dout1848,
   input         cfg_dout1849,
   input         cfg_dout1850,
   input         cfg_dout1851,
   input         cfg_dout1852,
   input         cfg_dout1853,
   input         cfg_dout1854,
   input         cfg_dout1855,
   input         cfg_dout1856,
   input         cfg_dout1857,
   input         cfg_dout1858,
   input         cfg_dout1859,
   input         cfg_dout1860,
   input         cfg_dout1861,
   input         cfg_dout1862,
   input         cfg_dout1863,
   input         cfg_dout1864,
   input         cfg_dout1865,
   input         cfg_dout1866,
   input         cfg_dout1867,
   input         cfg_dout1868,
   input         cfg_dout1869,
   input         cfg_dout1870,
   input         cfg_dout1871,
   input         cfg_dout1872,
   input         cfg_dout1873,
   input         cfg_dout1874,
   input         cfg_dout1875,
   input         cfg_dout1876,
   input         cfg_dout1877,
   input         cfg_dout1878,
   input         cfg_dout1879,
   input         cfg_dout1880,
   input         cfg_dout1881,
   input         cfg_dout1882,
   input         cfg_dout1883,
   input         cfg_dout1884,
   input         cfg_dout1885,
   input         cfg_dout1886,
   input         cfg_dout1887,
   input         cfg_dout1888,
   input         cfg_dout1889,
   input         cfg_dout1890,
   input         cfg_dout1891,
   input         cfg_dout1892,
   input         cfg_dout1893,
   input         cfg_dout1894,
   input         cfg_dout1895,
   input         cfg_dout1896,
   input         cfg_dout1897,
   input         cfg_dout1898,
   input         cfg_dout1899,
   input         cfg_dout1900,
   input         cfg_dout1901,
   input         cfg_dout1902,
   input         cfg_dout1903,
   input         cfg_dout1904,
   input         cfg_dout1905,
   input         cfg_dout1906,
   input         cfg_dout1907,
   input         cfg_dout1908,
   input         cfg_dout1909,
   input         cfg_dout1910,
   input         cfg_dout1911,
   input         cfg_dout1912,
   input         cfg_dout1913,
   input         cfg_dout1914,
   input         cfg_dout1915,
   input         cfg_dout1916,
   input         cfg_dout1917,
   input         cfg_dout1918,
   input         cfg_dout1919,
   input         cfg_dout1920,
   input         cfg_dout1921,
   input         cfg_dout1922,
   input         cfg_dout1923,
   input         cfg_dout1924,
   input         cfg_dout1925,
   input         cfg_dout1926,
   input         cfg_dout1927,
   input         cfg_dout1928,
   input         cfg_dout1929,
   input         cfg_dout1930,
   input         cfg_dout1931,
   input         cfg_dout1932,
   input         cfg_dout1933,
   input         cfg_dout1934,
   input         cfg_dout1935,
   input         cfg_dout1936,
   input         cfg_dout1937,
   input         cfg_dout1938,
   input         cfg_dout1939,
   input         cfg_dout1940,
   input         cfg_dout1941,
   input         cfg_dout1942,
   input         cfg_dout1943,
   input         cfg_dout1944,
   input         cfg_dout1945,
   input         cfg_dout1946,
   input         cfg_dout1947,
   input         cfg_dout1948,
   input         cfg_dout1949,
   input         cfg_dout1950,
   input         cfg_dout1951,
   input         cfg_dout1952,
   input         cfg_dout1953,
   input         cfg_dout1954,
   input         cfg_dout1955,
   input         cfg_dout1956,
   input         cfg_dout1957,
   input         cfg_dout1958,
   input         cfg_dout1959,
   input         cfg_dout1960,
   input         cfg_dout1961,
   input         cfg_dout1962,
   input         cfg_dout1963,
   input         cfg_dout1964,
   input         cfg_dout1965,
   input         cfg_dout1966,
   input         cfg_dout1967,
   input         cfg_dout1968,
   input         cfg_dout1969,
   input         cfg_dout1970,
   input         cfg_dout1971,
   input         cfg_dout1972,
   input         cfg_dout1973,
   input         cfg_dout1974,
   input         cfg_dout1975,
   input         cfg_dout1976,
   input         cfg_dout1977,
   input         cfg_dout1978,
   input         cfg_dout1979,
   input         cfg_dout1980,
   input         cfg_dout1981,
   input         cfg_dout1982,
   input         cfg_dout1983,
   input         cfg_dout1984,
   input         cfg_dout1985,
   input         cfg_dout1986,
   input         cfg_dout1987,
   input         cfg_dout1988,
   input         cfg_dout1989,
   input         cfg_dout1990,
   input         cfg_dout1991,
   input         cfg_dout1992,
   input         cfg_dout1993,
   input         cfg_dout1994,
   input         cfg_dout1995,
   input         cfg_dout1996,
   input         cfg_dout1997,
   input         cfg_dout1998,
   input         cfg_dout1999,
   input         cfg_dout2000,
   input         cfg_dout2001,
   input         cfg_dout2002,
   input         cfg_dout2003,
   input         cfg_dout2004,
   input         cfg_dout2005,
   input         cfg_dout2006,
   input         cfg_dout2007,
   input         cfg_dout2008,
   input         cfg_dout2009,
   input         cfg_dout2010,
   input         cfg_dout2011,
   input         cfg_dout2012,
   input         cfg_dout2013,
   input         cfg_dout2014,
   input         cfg_dout2015,
   input         cfg_dout2016,
   input         cfg_dout2017,
   input         cfg_dout2018,
   input         cfg_dout2019,
   input         cfg_dout2020,
   input         cfg_dout2021,
   input         cfg_dout2022,
   input         cfg_dout2023,
   input         cfg_dout2024,
   input         cfg_dout2025,
   input         cfg_dout2026,
   input         cfg_dout2027,
   input         cfg_dout2028,
   input         cfg_dout2029,
   input         cfg_dout2030,
   input         cfg_dout2031,
   input         cfg_dout2032,
   input         cfg_dout2033,
   input         cfg_dout2034,
   input         cfg_dout2035,
   input         cfg_dout2036,
   input         cfg_dout2037,
   input         cfg_dout2038,
   input         cfg_dout2039,
   input         cfg_dout2040,
   input         cfg_dout2041,
   input         cfg_dout2042,
   input         cfg_dout2043,
   input         cfg_dout2044,
   input         cfg_dout2045,
   input         cfg_dout2046,
   input         cfg_dout2047,
   input         cfg_dout2048,
   input         cfg_dout2049,
   input         cfg_dout2050,
   input         cfg_dout2051,
   input         cfg_dout2052,
   input         cfg_dout2053,
   input         cfg_dout2054,
   input         cfg_dout2055,
   input         cfg_dout2056,
   input         cfg_dout2057,
   input         cfg_dout2058,
   input         cfg_dout2059,
   input         cfg_dout2060,
   input         cfg_dout2061,
   input         cfg_dout2062,
   input         cfg_dout2063,
   input         cfg_dout2064,
   input         cfg_dout2065,
   input         cfg_dout2066,
   input         cfg_dout2067,
   input         cfg_dout2068,
   input         cfg_dout2069,
   input         cfg_dout2070,
   input         cfg_dout2071,
   input         cfg_dout2072,
   input         cfg_dout2073,
   input         cfg_dout2074,
   input         cfg_dout2075,
   input         cfg_dout2076,
   input         cfg_dout2077,
   input         cfg_dout2078,
   input         cfg_dout2079,
   input         cfg_dout2080,
   input         cfg_dout2081,
   input         cfg_dout2082,
   input         cfg_dout2083,
   input         cfg_dout2084,
   input         cfg_dout2085,
   input         cfg_dout2086,
   input         cfg_dout2087,
   input         cfg_dout2088,
   input         cfg_dout2089,
   input         cfg_dout2090,
   input         cfg_dout2091,
   input         cfg_dout2092,
   input         cfg_dout2093,
   input         cfg_dout2094,
   input         cfg_dout2095,
   input         cfg_dout2096,
   input         cfg_dout2097,
   input         cfg_dout2098,
   input         cfg_dout2099,
   input         cfg_dout2100,
   input         cfg_dout2101,
   input         cfg_dout2102,
   input         cfg_dout2103,
   input         cfg_dout2104,
   input         cfg_dout2105,
   input         cfg_dout2106,
   input         cfg_dout2107,
   input         cfg_dout2108,
   input         cfg_dout2109,
   input         cfg_dout2110,
   input         cfg_dout2111,
   input         cfg_dout2112,
   input         cfg_dout2113,
   input         cfg_dout2114,
   input         cfg_dout2115,
   input         cfg_dout2116,
   input         cfg_dout2117,
   input         cfg_dout2118,
   input         cfg_dout2119,
   input         cfg_dout2120,
   input         cfg_dout2121,
   input         cfg_dout2122,
   input         cfg_dout2123,
   input         cfg_dout2124,
   input         cfg_dout2125,
   input         cfg_dout2126,
   input         cfg_dout2127,
   input         cfg_dout2128,
   input         cfg_dout2129,
   input         cfg_dout2130,
   input         cfg_dout2131,
   input         cfg_dout2132,
   input         cfg_dout2133,
   input         cfg_dout2134,
   input         cfg_dout2135,
   input         cfg_dout2136,
   input         cfg_dout2137,
   input         cfg_dout2138,
   input         cfg_dout2139,
   input         cfg_dout2140,
   input         cfg_dout2141,
   input         cfg_dout2142,
   input         cfg_dout2143,
   input         cfg_dout2144,
   input         cfg_dout2145,
   input         cfg_dout2146,
   input         cfg_dout2147,
   input         cfg_dout2148,
   input         cfg_dout2149,
   input         cfg_dout2150,
   input         cfg_dout2151,
   input         cfg_dout2152,
   input         cfg_dout2153,
   input         cfg_dout2154,
   input         cfg_dout2155,
   input         cfg_dout2156,
   input         cfg_dout2157,
   input         cfg_dout2158,
   input         cfg_dout2159,
   input         cfg_dout2160,
   input         cfg_dout2161,
   input         cfg_dout2162,
   input         cfg_dout2163,
   input         cfg_dout2164,
   input         cfg_dout2165,
   input         cfg_dout2166,
   input         cfg_dout2167,
   input         cfg_dout2168,
   input         cfg_dout2169,
   input         cfg_dout2170,
   input         cfg_dout2171,
   input         cfg_dout2172,
   input         cfg_dout2173,
   input         cfg_dout2174,
   input         cfg_dout2175,
   input         cfg_dout2176,
   input         cfg_dout2177,
   input         cfg_dout2178,
   input         cfg_dout2179,
   input         cfg_dout2180,
   input         cfg_dout2181,
   input         cfg_dout2182,
   input         cfg_dout2183,
   input         cfg_dout2184,
   input         cfg_dout2185,
   input         cfg_dout2186,
   input         cfg_dout2187,
   input         cfg_dout2188,
   input         cfg_dout2189,
   input         cfg_dout2190,
   input         cfg_dout2191,
   input         cfg_dout2192,
   input         cfg_dout2193,
   input         cfg_dout2194,
   input         cfg_dout2195,
   input         cfg_dout2196,
   input         cfg_dout2197,
   input         cfg_dout2198,
   input         cfg_dout2199,
   input         cfg_dout2200,
   input         cfg_dout2201,
   input         cfg_dout2202,
   input         cfg_dout2203,
   input         cfg_dout2204,
   input         cfg_dout2205,
   input         cfg_dout2206,
   input         cfg_dout2207,
   input         cfg_dout2208,
   input         cfg_dout2209,
   input         cfg_dout2210,
   input         cfg_dout2211,
   input         cfg_dout2212,
   input         cfg_dout2213,
   input         cfg_dout2214,
   input         cfg_dout2215,
   input         cfg_dout2216,
   input         cfg_dout2217,
   input         cfg_dout2218,
   input         cfg_dout2219,
   input         cfg_dout2220,
   input         cfg_dout2221,
   input         cfg_dout2222,
   input         cfg_dout2223,
   input         cfg_dout2224,
   input         cfg_dout2225,
   input         cfg_dout2226,
   input         cfg_dout2227,
   input         cfg_dout2228,
   input         cfg_dout2229,
   input         cfg_dout2230,
   input         cfg_dout2231,
   input         cfg_dout2232,
   input         cfg_dout2233,
   input         cfg_dout2234,
   input         cfg_dout2235,
   input         cfg_dout2236,
   input         cfg_dout2237,
   input         cfg_dout2238,
   input         cfg_dout2239,
   input         cfg_dout2240,
   input         cfg_dout2241,
   input         cfg_dout2242,
   input         cfg_dout2243,
   input         cfg_dout2244,
   input         cfg_dout2245,
   input         cfg_dout2246,
   input         cfg_dout2247,
   input         cfg_dout2248,
   input         cfg_dout2249,
   input         cfg_dout2250,
   input         cfg_dout2251,
   input         cfg_dout2252,
   input         cfg_dout2253,
   input         cfg_dout2254,
   input         cfg_dout2255,
   input         cfg_dout2256,
   input         cfg_dout2257,
   input         cfg_dout2258,
   input         cfg_dout2259,
   input         cfg_dout2260,
   input         cfg_dout2261,
   input         cfg_dout2262,
   input         cfg_dout2263,
   input         cfg_dout2264,
   input         cfg_dout2265,
   input         cfg_dout2266,
   input         cfg_dout2267,
   input         cfg_dout2268,
   input         cfg_dout2269,
   input         cfg_dout2270,
   input         cfg_dout2271,
   input         cfg_dout2272,
   input         cfg_dout2273,
   input         cfg_dout2274,
   input         cfg_dout2275,
   input         cfg_dout2276,
   input         cfg_dout2277,
   input         cfg_dout2278,
   input         cfg_dout2279,
   input         cfg_dout2280,
   input         cfg_dout2281,
   input         cfg_dout2282,
   input         cfg_dout2283,
   input         cfg_dout2284,
   input         cfg_dout2285,
   input         cfg_dout2286,
   input         cfg_dout2287,
   input         cfg_dout2288,
   input         cfg_dout2289,
   input         cfg_dout2290,
   input         cfg_dout2291,
   input         cfg_dout2292,
   input         cfg_dout2293,
   input         cfg_dout2294,
   input         cfg_dout2295,
   input         cfg_dout2296,
   input         cfg_dout2297,
   input         cfg_dout2298,
   input         cfg_dout2299,
   input         cfg_dout2300,
   input         cfg_dout2301,
   input         cfg_dout2302,
   input         cfg_dout2303,
   input         cfg_dout2304,
   input         cfg_dout2305,
   input         cfg_dout2306,
   input         cfg_dout2307,
   input         cfg_dout2308,
   input         cfg_dout2309,
   input         cfg_dout2310,
   input         cfg_dout2311,
   input         cfg_dout2312,
   input         cfg_dout2313,
   input         cfg_dout2314,
   input         cfg_dout2315,
   input         cfg_dout2316,
   input         cfg_dout2317,
   input         cfg_dout2318,
   input         cfg_dout2319,
   input         cfg_dout2320,
   input         cfg_dout2321,
   input         cfg_dout2322,
   input         cfg_dout2323,
   input         cfg_dout2324,
   input         cfg_dout2325,
   input         cfg_dout2326,
   input         cfg_dout2327,
   input         cfg_dout2328,
   input         cfg_dout2329,
   input         cfg_dout2330,
   input         cfg_dout2331,
   input         cfg_dout2332,
   input         cfg_dout2333,
   input         cfg_dout2334,
   input         cfg_dout2335,
   input         cfg_dout2336,
   input         cfg_dout2337,
   input         cfg_dout2338,
   input         cfg_dout2339,
   input         cfg_dout2340,
   input         cfg_dout2341,
   input         cfg_dout2342,
   input         cfg_dout2343,
   input         cfg_dout2344,
   input         cfg_dout2345,
   input         cfg_dout2346,
   input         cfg_dout2347,
   input         cfg_dout2348,
   input         cfg_dout2349,
   input         cfg_dout2350,
   input         cfg_dout2351,
   input         cfg_dout2352,
   input         cfg_dout2353,
   input         cfg_dout2354,
   input         cfg_dout2355,
   input         cfg_dout2356,
   input         cfg_dout2357,
   input         cfg_dout2358,
   input         cfg_dout2359,
   input         cfg_dout2360,
   input         cfg_dout2361,
   input         cfg_dout2362,
   input         cfg_dout2363,
   input         cfg_dout2364,
   input         cfg_dout2365,
   input         cfg_dout2366,
   input         cfg_dout2367,
   input         cfg_dout2368,
   input         cfg_dout2369,
   input         cfg_dout2370,
   input         cfg_dout2371,
   input         cfg_dout2372,
   input         cfg_dout2373,
   input         cfg_dout2374,
   input         cfg_dout2375,
   input         cfg_dout2376,
   input         cfg_dout2377,
   input         cfg_dout2378,
   input         cfg_dout2379,
   input         cfg_dout2380,
   input         cfg_dout2381,
   input         cfg_dout2382,
   input         cfg_dout2383,
   input         cfg_dout2384,
   input         cfg_dout2385,
   input         cfg_dout2386,
   input         cfg_dout2387,
   input         cfg_dout2388,
   input         cfg_dout2389,
   input         cfg_dout2390,
   input         cfg_dout2391,
   input         cfg_dout2392,
   input         cfg_dout2393,
   input         cfg_dout2394,
   input         cfg_dout2395,
   input         cfg_dout2396,
   input         cfg_dout2397,
   input         cfg_dout2398,
   input         cfg_dout2399,
   input         cfg_dout2400,
   input         cfg_dout2401,
   input         cfg_dout2402,
   input         cfg_dout2403,
   input         cfg_dout2404,
   input         cfg_dout2405,
   input         cfg_dout2406,
   input         cfg_dout2407,
   input         cfg_dout2408,
   input         cfg_dout2409,
   input         cfg_dout2410,
   input         cfg_dout2411,
   input         cfg_dout2412,
   input         cfg_dout2413,
   input         cfg_dout2414,
   input         cfg_dout2415,
   input         cfg_dout2416,
   input         cfg_dout2417,
   input         cfg_dout2418,
   input         cfg_dout2419,
   input         cfg_dout2420,
   input         cfg_dout2421,
   input         cfg_dout2422,
   input         cfg_dout2423,
   input         cfg_dout2424,
   input         cfg_dout2425,
   input         cfg_dout2426,
   input         cfg_dout2427,
   input         cfg_dout2428,
   input         cfg_dout2429,
   input         cfg_dout2430,
   input         cfg_dout2431,
   input         cfg_dout2432,
   input         cfg_dout2433,
   input         cfg_dout2434,
   input         cfg_dout2435,
   input         cfg_dout2436,
   input         cfg_dout2437,
   input         cfg_dout2438,
   input         cfg_dout2439,
   input         cfg_dout2440,
   input         cfg_dout2441,
   input         cfg_dout2442,
   input         cfg_dout2443,
   input         cfg_dout2444,
   input         cfg_dout2445,
   input         cfg_dout2446,
   input         cfg_dout2447,
   input         cfg_dout2448,
   input         cfg_dout2449,
   input         cfg_dout2450,
   input         cfg_dout2451,
   input         cfg_dout2452,
   input         cfg_dout2453,
   input         cfg_dout2454,
   input         cfg_dout2455,
   input         cfg_dout2456,
   input         cfg_dout2457,
   input         cfg_dout2458,
   input         cfg_dout2459,
   input         cfg_dout2460,
   input         cfg_dout2461,
   input         cfg_dout2462,
   input         cfg_dout2463,
   input         cfg_dout2464,
   input         cfg_dout2465,
   input         cfg_dout2466,
   input         cfg_dout2467,
   input         cfg_dout2468,
   input         cfg_dout2469,
   input         cfg_dout2470,
   input         cfg_dout2471,
   input         cfg_dout2472,
   input         cfg_dout2473,
   input         cfg_dout2474,
   input         cfg_dout2475,
   input         cfg_dout2476,
   input         cfg_dout2477,
   input         cfg_dout2478,
   input         cfg_dout2479,
   input         cfg_dout2480,
   input         cfg_dout2481,
   input         cfg_dout2482,
   input         cfg_dout2483,
   input         cfg_dout2484,
   input         cfg_dout2485,
   input         cfg_dout2486,
   input         cfg_dout2487,
   input         cfg_dout2488,
   input         cfg_dout2489,
   input         cfg_dout2490,
   input         cfg_dout2491,
   input         cfg_dout2492,
   input         cfg_dout2493,
   input         cfg_dout2494,
   input         cfg_dout2495,
   input         cfg_dout2496,
   input         cfg_dout2497,
   input         cfg_dout2498,
   input         cfg_dout2499,
   input         cfg_dout2500,
   input         cfg_dout2501,
   input         cfg_dout2502,
   input         cfg_dout2503,
   input         cfg_dout2504,
   input         cfg_dout2505,
   input         cfg_dout2506,
   input         cfg_dout2507,
   input         cfg_dout2508,
   input         cfg_dout2509,
   input         cfg_dout2510,
   input         cfg_dout2511,
   input         cfg_dout2512,
   input         cfg_dout2513,
   input         cfg_dout2514,
   input         cfg_dout2515,
   input         cfg_dout2516,
   input         cfg_dout2517,
   input         cfg_dout2518,
   input         cfg_dout2519,
   input         cfg_dout2520,
   input         cfg_dout2521,
   input         cfg_dout2522,
   input         cfg_dout2523,
   input         cfg_dout2524,
   input         cfg_dout2525,
   input         cfg_dout2526,
   input         cfg_dout2527,
   input         cfg_dout2528,
   input         cfg_dout2529,
   input         cfg_dout2530,
   input         cfg_dout2531,
   input         cfg_dout2532,
   input         cfg_dout2533,
   input         cfg_dout2534,
   input         cfg_dout2535,
   input         cfg_dout2536,
   input         cfg_dout2537,
   input         cfg_dout2538,
   input         cfg_dout2539,
   input         cfg_dout2540,
   input         cfg_dout2541,
   input         cfg_dout2542,
   input         cfg_dout2543,
   input         cfg_dout2544,
   input         cfg_dout2545,
   input         cfg_dout2546,
   input         cfg_dout2547,
   input         cfg_dout2548,
   input         cfg_dout2549,
   input         cfg_dout2550,
   input         cfg_dout2551,
   input         cfg_dout2552,
   input         cfg_dout2553,
   input         cfg_dout2554,
   input         cfg_dout2555,
   input         cfg_dout2556,
   input         cfg_dout2557,
   input         cfg_dout2558,
   input         cfg_dout2559,
   input         cfg_dout2560,
   input         cfg_dout2561,
   input         cfg_dout2562,
   input         cfg_dout2563,
   input         cfg_dout2564,
   input         cfg_dout2565,
   input         cfg_dout2566,
   input         cfg_dout2567,
   input         cfg_dout2568,
   input         cfg_dout2569,
   input         cfg_dout2570,
   input         cfg_dout2571,
   input         cfg_dout2572,
   input         cfg_dout2573,
   input         cfg_dout2574,
   input         cfg_dout2575,
   input         cfg_dout2576,
   input         cfg_dout2577,
   input         cfg_dout2578,
   input         cfg_dout2579,
   input         cfg_dout2580,
   input         cfg_dout2581,
   input         cfg_dout2582,
   input         cfg_dout2583,
   input         cfg_dout2584,
   input         cfg_dout2585,
   input         cfg_dout2586,
   input         cfg_dout2587,
   input         cfg_dout2588,
   input         cfg_dout2589,
   input         cfg_dout2590,
   input         cfg_dout2591,
   input         cfg_dout2592,
   input         cfg_dout2593,
   input         cfg_dout2594,
   input         cfg_dout2595,
   input         cfg_dout2596,
   input         cfg_dout2597,
   input         cfg_dout2598,
   input         cfg_dout2599,
   input         cfg_dout2600,
   input         cfg_dout2601,
   input         cfg_dout2602,
   input         cfg_dout2603,
   input         cfg_dout2604,
   input         cfg_dout2605,
   input         cfg_dout2606,
   input         cfg_dout2607,
   input         cfg_dout2608,
   input         cfg_dout2609,
   input         cfg_dout2610,
   input         cfg_dout2611,
   input         cfg_dout2612,
   input         cfg_dout2613,
   input         cfg_dout2614,
   input         cfg_dout2615,
   input         cfg_dout2616,
   input         cfg_dout2617,
   input         cfg_dout2618,
   input         cfg_dout2619,
   input         cfg_dout2620,
   input         cfg_dout2621,
   input         cfg_dout2622,
   input         cfg_dout2623,
   input         cfg_dout2624,
   input         cfg_dout2625,
   input         cfg_dout2626,
   input         cfg_dout2627,
   input         cfg_dout2628,
   input         cfg_dout2629,
   input         cfg_dout2630,
   input         cfg_dout2631,
   input         cfg_dout2632,
   input         cfg_dout2633,
   input         cfg_dout2634,
   input         cfg_dout2635,
   input         cfg_dout2636,
   input         cfg_dout2637,
   input         cfg_dout2638,
   input         cfg_dout2639,
   input         cfg_dout2640,
   input         cfg_dout2641,
   input         cfg_dout2642,
   input         cfg_dout2643,
   input         cfg_dout2644,
   input         cfg_dout2645,
   input         cfg_dout2646,
   input         cfg_dout2647,
   input         cfg_dout2648,
   input         cfg_dout2649,
   input         cfg_dout2650,
   input         cfg_dout2651,
   input         cfg_dout2652,
   input         cfg_dout2653,
   input         cfg_dout2654,
   input         cfg_dout2655,
   input         cfg_dout2656,
   input         cfg_dout2657,
   input         cfg_dout2658,
   input         cfg_dout2659,
   input         cfg_dout2660,
   input         cfg_dout2661,
   input         cfg_dout2662,
   input         cfg_dout2663,
   input         cfg_dout2664,
   input         cfg_dout2665,
   input         cfg_dout2666,
   input         cfg_dout2667,
   input         cfg_dout2668,
   input         cfg_dout2669,
   input         cfg_dout2670,
   input         cfg_dout2671,
   input         cfg_dout2672,
   input         cfg_dout2673,
   input         cfg_dout2674,
   input         cfg_dout2675,
   input         cfg_dout2676,
   input         cfg_dout2677,
   input         cfg_dout2678,
   input         cfg_dout2679,
   input         cfg_dout2680,
   input         cfg_dout2681,
   input         cfg_dout2682,
   input         cfg_dout2683,
   input         cfg_dout2684,
   input         cfg_dout2685,
   input         cfg_dout2686,
   input         cfg_dout2687,
   input         cfg_dout2688,
   input         cfg_dout2689,
   input         cfg_dout2690,
   input         cfg_dout2691,
   input         cfg_dout2692,
   input         cfg_dout2693,
   input         cfg_dout2694,
   input         cfg_dout2695,
   input         cfg_dout2696,
   input         cfg_dout2697,
   input         cfg_dout2698,
   input         cfg_dout2699,
   input         cfg_dout2700,
   input         cfg_dout2701,
   input         cfg_dout2702,
   input         cfg_dout2703,
   input         cfg_dout2704,
   input         cfg_dout2705,
   input         cfg_dout2706,
   input         cfg_dout2707,
   input         cfg_dout2708,
   input         cfg_dout2709,
   input         cfg_dout2710,
   input         cfg_dout2711,
   input         cfg_dout2712,
   input         cfg_dout2713,
   input         cfg_dout2714,
   input         cfg_dout2715,
   input         cfg_dout2716,
   input         cfg_dout2717,
   input         cfg_dout2718,
   input         cfg_dout2719,
   input         cfg_dout2720,
   input         cfg_dout2721,
   input         cfg_dout2722,
   input         cfg_dout2723,
   input         cfg_dout2724,
   input         cfg_dout2725,
   input         cfg_dout2726,
   input         cfg_dout2727,
   input         cfg_dout2728,
   input         cfg_dout2729,
   input         cfg_dout2730,
   input         cfg_dout2731,
   input         cfg_dout2732,
   input         cfg_dout2733,
   input         cfg_dout2734,
   input         cfg_dout2735,
   input         cfg_dout2736,
   input         cfg_dout2737,
   input         cfg_dout2738,
   input         cfg_dout2739,
   input         cfg_dout2740,
   input         cfg_dout2741,
   input         cfg_dout2742,
   input         cfg_dout2743,
   input         cfg_dout2744,
   input         cfg_dout2745,
   input         cfg_dout2746,
   input         cfg_dout2747,
   input         cfg_dout2748,
   input         cfg_dout2749,
   input         cfg_dout2750,
   input         cfg_dout2751,
   input         cfg_dout2752,
   input         cfg_dout2753,
   input         cfg_dout2754,
   input         cfg_dout2755,
   input         cfg_dout2756,
   input         cfg_dout2757,
   input         cfg_dout2758,
   input         cfg_dout2759,
   input         cfg_dout2760,
   input         cfg_dout2761,
   input         cfg_dout2762,
   input         cfg_dout2763,
   input         cfg_dout2764,
   input         cfg_dout2765,
   input         cfg_dout2766,
   input         cfg_dout2767,
   input         cfg_dout2768,
   input         cfg_dout2769,
   input         cfg_dout2770,
   input         cfg_dout2771,
   input         cfg_dout2772,
   input         cfg_dout2773,
   input         cfg_dout2774,
   input         cfg_dout2775,
   input         cfg_dout2776,
   input         cfg_dout2777,
   input         cfg_dout2778,
   input         cfg_dout2779,
   input         cfg_dout2780,
   input         cfg_dout2781,
   input         cfg_dout2782,
   input         cfg_dout2783,
   input         cfg_dout2784,
   input         cfg_dout2785,
   input         cfg_dout2786,
   input         cfg_dout2787,
   input         cfg_dout2788,
   input         cfg_dout2789,
   input         cfg_dout2790,
   input         cfg_dout2791,
   input         cfg_dout2792,
   input         cfg_dout2793,
   input         cfg_dout2794,
   input         cfg_dout2795,
   input         cfg_dout2796,
   input         cfg_dout2797,
   input         cfg_dout2798,
   input         cfg_dout2799,
   input         cfg_dout2800,
   input         cfg_dout2801,
   input         cfg_dout2802,
   input         cfg_dout2803,
   input         cfg_dout2804,
   input         cfg_dout2805,
   input         cfg_dout2806,
   input         cfg_dout2807,
   input         cfg_dout2808,
   input         cfg_dout2809,
   input         cfg_dout2810,
   input         cfg_dout2811,
   input         cfg_dout2812,
   input         cfg_dout2813,
   input         cfg_dout2814,
   input         cfg_dout2815,
   input         cfg_dout2816,
   input         cfg_dout2817,
   input         cfg_dout2818,
   input         cfg_dout2819,
   input         cfg_dout2820,
   input         cfg_dout2821,
   input         cfg_dout2822,
   input         cfg_dout2823,
   input         cfg_dout2824,
   input         cfg_dout2825,
   input         cfg_dout2826,
   input         cfg_dout2827,
   input         cfg_dout2828,
   input         cfg_dout2829,
   input         cfg_dout2830,
   input         cfg_dout2831,
   input         cfg_dout2832,
   input         cfg_dout2833,
   input         cfg_dout2834,
   input         cfg_dout2835,
   input         cfg_dout2836,
   input         cfg_dout2837,
   input         cfg_dout2838,
   input         cfg_dout2839,
   input         cfg_dout2840,
   input         cfg_dout2841,
   input         cfg_dout2842,
   input         cfg_dout2843,
   input         cfg_dout2844,
   input         cfg_dout2845,
   input         cfg_dout2846,
   input         cfg_dout2847,
   input         cfg_dout2848,
   input         cfg_dout2849,
   input         cfg_dout2850,
   input         cfg_dout2851,
   input         cfg_dout2852,
   input         cfg_dout2853,
   input         cfg_dout2854,
   input         cfg_dout2855,
   input         cfg_dout2856,
   input         cfg_dout2857,
   input         cfg_dout2858,
   input         cfg_dout2859,
   input         cfg_dout2860,
   input         cfg_dout2861,
   input         cfg_dout2862,
   input         cfg_dout2863,
   input         cfg_dout2864,
   input         cfg_dout2865,
   input         cfg_dout2866,
   input         cfg_dout2867,
   input         cfg_dout2868,
   input         cfg_dout2869,
   input         cfg_dout2870,
   input         cfg_dout2871,
   input         cfg_dout2872,
   input         cfg_dout2873,
   input         cfg_dout2874,
   input         cfg_dout2875,
   input         cfg_dout2876,
   input         cfg_dout2877,
   input         cfg_dout2878,
   input         cfg_dout2879,
   input         cfg_dout2880,
   input         cfg_dout2881,
   input         cfg_dout2882,
   input         cfg_dout2883,
   input         cfg_dout2884,
   input         cfg_dout2885,
   input         cfg_dout2886,
   input         cfg_dout2887,
   input         cfg_dout2888,
   input         cfg_dout2889,
   input         cfg_dout2890,
   input         cfg_dout2891,
   input         cfg_dout2892,
   input         cfg_dout2893,
   input         cfg_dout2894,
   input         cfg_dout2895,
   input         cfg_dout2896,
   input         cfg_dout2897,
   input         cfg_dout2898,
   input         cfg_dout2899,
   input         cfg_dout2900,
   input         cfg_dout2901,
   input         cfg_dout2902,
   input         cfg_dout2903,
   input         cfg_dout2904,
   input         cfg_dout2905,
   input         cfg_dout2906,
   input         cfg_dout2907,
   input         cfg_dout2908,
   input         cfg_dout2909,
   input         cfg_dout2910,
   input         cfg_dout2911,
   input         cfg_dout2912,
   input         cfg_dout2913,
   input         cfg_dout2914,
   input         cfg_dout2915,
   input         cfg_dout2916,
   input         cfg_dout2917,
   input         cfg_dout2918,
   input         cfg_dout2919,
   input         cfg_dout2920,
   input         cfg_dout2921,
   input         cfg_dout2922,
   input         cfg_dout2923,
   input         cfg_dout2924,
   input         cfg_dout2925,
   input         cfg_dout2926,
   input         cfg_dout2927,
   input         cfg_dout2928,
   input         cfg_dout2929,
   input         cfg_dout2930,
   input         cfg_dout2931,
   input         cfg_dout2932,
   input         cfg_dout2933,
   input         cfg_dout2934,
   input         cfg_dout2935,
   input         cfg_dout2936,
   input         cfg_dout2937,
   input         cfg_dout2938,
   input         cfg_dout2939,
   input         cfg_dout2940,
   input         cfg_dout2941,
   input         cfg_dout2942,
   input         cfg_dout2943,
   input         cfg_dout2944,
   input         cfg_dout2945,
   input         cfg_dout2946,
   input         cfg_dout2947,
   input         cfg_dout2948,
   input         cfg_dout2949,
   input         cfg_dout2950,
   input         cfg_dout2951,
   input         cfg_dout2952,
   input         cfg_dout2953,
   input         cfg_dout2954,
   input         cfg_dout2955,
   input         cfg_dout2956,
   input         cfg_dout2957,
   input         cfg_dout2958,
   input         cfg_dout2959,
   input         cfg_dout2960,
   input         cfg_dout2961,
   input         cfg_dout2962,
   input         cfg_dout2963,
   input         cfg_dout2964,
   input         cfg_dout2965,
   input         cfg_dout2966,
   input         cfg_dout2967,
   input         cfg_dout2968,
   input         cfg_dout2969,
   input         cfg_dout2970,
   input         cfg_dout2971,
   input         cfg_dout2972,
   input         cfg_dout2973,
   input         cfg_dout2974,
   input         cfg_dout2975,
   input         cfg_dout2976,
   input         cfg_dout2977,
   input         cfg_dout2978,
   input         cfg_dout2979,
   input         cfg_dout2980,
   input         cfg_dout2981,
   input         cfg_dout2982,
   input         cfg_dout2983,
   input         cfg_dout2984,
   input         cfg_dout2985,
   input         cfg_dout2986,
   input         cfg_dout2987,
   input         cfg_dout2988,
   input         cfg_dout2989,
   input         cfg_dout2990,
   input         cfg_dout2991,
   input         cfg_dout2992,
   input         cfg_dout2993,
   input         cfg_dout2994,
   input         cfg_dout2995,
   input         cfg_dout2996,
   input         cfg_dout2997,
   input         cfg_dout2998,
   input         cfg_dout2999,
   input         cfg_dout3000,
   input         cfg_dout3001,
   input         cfg_dout3002,
   input         cfg_dout3003,
   input         cfg_dout3004,
   input         cfg_dout3005,
   input         cfg_dout3006,
   input         cfg_dout3007,
   input         cfg_dout3008,
   input         cfg_dout3009,
   input         cfg_dout3010,
   input         cfg_dout3011,
   input         cfg_dout3012,
   input         cfg_dout3013,
   input         cfg_dout3014,
   input         cfg_dout3015,
   input         cfg_dout3016,
   input         cfg_dout3017,
   input         cfg_dout3018,
   input         cfg_dout3019,
   input         cfg_dout3020,
   input         cfg_dout3021,
   input         cfg_dout3022,
   input         cfg_dout3023,
   input         cfg_dout3024,
   input         cfg_dout3025,
   input         cfg_dout3026,
   input         cfg_dout3027,
   input         cfg_dout3028,
   input         cfg_dout3029,
   input         cfg_dout3030,
   input         cfg_dout3031,
   input         cfg_dout3032,
   input         cfg_dout3033,
   input         cfg_dout3034,
   input         cfg_dout3035,
   input         cfg_dout3036,
   input         cfg_dout3037,
   input         cfg_dout3038,
   input         cfg_dout3039,
   input         cfg_dout3040,
   input         cfg_dout3041,
   input         cfg_dout3042,
   input         cfg_dout3043,
   input         cfg_dout3044,
   input         cfg_dout3045,
   input         cfg_dout3046,
   input         cfg_dout3047,
   input         cfg_dout3048,
   input         cfg_dout3049,
   input         cfg_dout3050,
   input         cfg_dout3051,
   input         cfg_dout3052,
   input         cfg_dout3053,
   input         cfg_dout3054,
   input         cfg_dout3055,
   input         cfg_dout3056,
   input         cfg_dout3057,
   input         cfg_dout3058,
   input         cfg_dout3059,
   input         cfg_dout3060,
   input         cfg_dout3061,
   input         cfg_dout3062,
   input         cfg_dout3063,
   input         cfg_dout3064,
   input         cfg_dout3065,
   input         cfg_dout3066,
   input         cfg_dout3067,
   input         cfg_dout3068,
   input         cfg_dout3069,
   input         cfg_dout3070,
   input         cfg_dout3071,
   input         cfg_dout3072,
   input         cfg_dout3073,
   input         cfg_dout3074,
   input         cfg_dout3075,
   input         cfg_dout3076,
   input         cfg_dout3077,
   input         cfg_dout3078,
   input         cfg_dout3079,
   input         cfg_dout3080,
   input         cfg_dout3081,
   input         cfg_dout3082,
   input         cfg_dout3083,
   input         cfg_dout3084,
   input         cfg_dout3085,
   input         cfg_dout3086,
   input         cfg_dout3087,
   input         cfg_dout3088,
   input         cfg_dout3089,
   input         cfg_dout3090,
   input         cfg_dout3091,
   input         cfg_dout3092,
   input         cfg_dout3093,
   input         cfg_dout3094,
   input         cfg_dout3095,
   input         cfg_dout3096,
   input         cfg_dout3097,
   input         cfg_dout3098,
   input         cfg_dout3099,
   input         cfg_dout3100,
   input         cfg_dout3101,
   input         cfg_dout3102,
   input         cfg_dout3103,
   input         cfg_dout3104,
   input         cfg_dout3105,
   input         cfg_dout3106,
   input         cfg_dout3107,
   input         cfg_dout3108,
   input         cfg_dout3109,
   input         cfg_dout3110,
   input         cfg_dout3111,
   input         cfg_dout3112,
   input         cfg_dout3113,
   input         cfg_dout3114,
   input         cfg_dout3115,
   input         cfg_dout3116,
   input         cfg_dout3117,
   input         cfg_dout3118,
   input         cfg_dout3119,
   input         cfg_dout3120,
   input         cfg_dout3121,
   input         cfg_dout3122,
   input         cfg_dout3123,
   input         cfg_dout3124,
   input         cfg_dout3125,
   input         cfg_dout3126,
   input         cfg_dout3127,
   input         cfg_dout3128,
   input         cfg_dout3129,
   input         cfg_dout3130,
   input         cfg_dout3131,
   input         cfg_dout3132,
   input         cfg_dout3133,
   input         cfg_dout3134,
   input         cfg_dout3135,
   input         cfg_dout3136,
   input         cfg_dout3137,
   input         cfg_dout3138,
   input         cfg_dout3139,
   input         cfg_dout3140,
   input         cfg_dout3141,
   input         cfg_dout3142,
   input         cfg_dout3143,
   input         cfg_dout3144,
   input         cfg_dout3145,
   input         cfg_dout3146,
   input         cfg_dout3147,
   input         cfg_dout3148,
   input         cfg_dout3149,
   input         cfg_dout3150,
   input         cfg_dout3151,
   input         cfg_dout3152,
   input         cfg_dout3153,
   input         cfg_dout3154,
   input         cfg_dout3155,
   input         cfg_dout3156,
   input         cfg_dout3157,
   input         cfg_dout3158,
   input         cfg_dout3159,
   input         cfg_dout3160,
   input         cfg_dout3161,
   input         cfg_dout3162,
   input         cfg_dout3163,
   input         cfg_dout3164,
   input         cfg_dout3165,
   input         cfg_dout3166,
   input         cfg_dout3167,
   input         cfg_dout3168,
   input         cfg_dout3169,
   input         cfg_dout3170,
   input         cfg_dout3171,
   input         cfg_dout3172,
   input         cfg_dout3173,
   input         cfg_dout3174,
   input         cfg_dout3175,
   input         cfg_dout3176,
   input         cfg_dout3177,
   input         cfg_dout3178,
   input         cfg_dout3179,
   input         cfg_dout3180,
   input         cfg_dout3181,
   input         cfg_dout3182,
   input         cfg_dout3183,
   input         cfg_dout3184,
   input         cfg_dout3185,
   input         cfg_dout3186,
   input         cfg_dout3187,
   input         cfg_dout3188,
   input         cfg_dout3189,
   input         cfg_dout3190,
   input         cfg_dout3191,
   input         cfg_dout3192,
   input         cfg_dout3193,
   input         cfg_dout3194,
   input         cfg_dout3195,
   input         cfg_dout3196,
   input         cfg_dout3197,
   input         cfg_dout3198,
   input         cfg_dout3199,
   input         cfg_dout3200,
   input         cfg_dout3201,
   input         cfg_dout3202,
   input         cfg_dout3203,
   input         cfg_dout3204,
   input         cfg_dout3205,
   input         cfg_dout3206,
   input         cfg_dout3207,
   input         cfg_dout3208,
   input         cfg_dout3209,
   input         cfg_dout3210,
   input         cfg_dout3211,
   input         cfg_dout3212,
   input         cfg_dout3213,
   input         cfg_dout3214,
   input         cfg_dout3215,
   input         cfg_dout3216,
   input         cfg_dout3217,
   input         cfg_dout3218,
   input         cfg_dout3219,
   input         cfg_dout3220,
   input         cfg_dout3221,
   input         cfg_dout3222,
   input         cfg_dout3223,
   input         cfg_dout3224,
   input         cfg_dout3225,
   input         cfg_dout3226,
   input         cfg_dout3227,
   input         cfg_dout3228,
   input         cfg_dout3229,
   input         cfg_dout3230,
   input         cfg_dout3231,
   input         cfg_dout3232,
   input         cfg_dout3233,
   input         cfg_dout3234,
   input         cfg_dout3235,
   input         cfg_dout3236,
   input         cfg_dout3237,
   input         cfg_dout3238,
   input         cfg_dout3239,
   input         cfg_dout3240,
   input         cfg_dout3241,
   input         cfg_dout3242,
   input         cfg_dout3243,
   input         cfg_dout3244,
   input         cfg_dout3245,
   input         cfg_dout3246,
   input         cfg_dout3247,
   input         cfg_dout3248,
   input         cfg_dout3249,
   input         cfg_dout3250,
   input         cfg_dout3251,
   input         cfg_dout3252,
   input         cfg_dout3253,
   input         cfg_dout3254,
   input         cfg_dout3255,
   input         cfg_dout3256,
   input         cfg_dout3257,
   input         cfg_dout3258,
   input         cfg_dout3259,
   input         cfg_dout3260,
   input         cfg_dout3261,
   input         cfg_dout3262,
   input         cfg_dout3263,
   input         cfg_dout3264,
   input         cfg_dout3265,
   input         cfg_dout3266,
   input         cfg_dout3267,
   input         cfg_dout3268,
   input         cfg_dout3269,
   input         cfg_dout3270,
   input         cfg_dout3271,
   input         cfg_dout3272,
   input         cfg_dout3273,
   input         cfg_dout3274,
   input         cfg_dout3275,
   input         cfg_dout3276,
   input         cfg_dout3277,
   input         cfg_dout3278,
   input         cfg_dout3279,
   input         cfg_dout3280,
   input         cfg_dout3281,
   input         cfg_dout3282,
   input         cfg_dout3283,
   input         cfg_dout3284,
   input         cfg_dout3285,
   input         cfg_dout3286,
   input         cfg_dout3287,
   input         cfg_dout3288,
   input         cfg_dout3289,
   input         cfg_dout3290,
   input         cfg_dout3291,
   input         cfg_dout3292,
   input         cfg_dout3293,
   input         cfg_dout3294,
   input         cfg_dout3295,
   input         cfg_dout3296,
   input         cfg_dout3297,
   input         cfg_dout3298,
   input         cfg_dout3299,
   input         cfg_dout3300,
   input         cfg_dout3301,
   input         cfg_dout3302,
   input         cfg_dout3303,
   input         cfg_dout3304,
   input         cfg_dout3305,
   input         cfg_dout3306,
   input         cfg_dout3307,
   input         cfg_dout3308,
   input         cfg_dout3309,
   input         cfg_dout3310,
   input         cfg_dout3311,
   input         cfg_dout3312,
   input         cfg_dout3313,
   input         cfg_dout3314,
   input         cfg_dout3315,
   input         cfg_dout3316,
   input         cfg_dout3317,
   input         cfg_dout3318,
   input         cfg_dout3319,
   input         cfg_dout3320,
   input         cfg_dout3321,
   input         cfg_dout3322,
   input         cfg_dout3323,
   input         cfg_dout3324,
   input         cfg_dout3325,
   input         cfg_dout3326,
   input         cfg_dout3327,
   input         cfg_dout3328,
   input         cfg_dout3329,
   input         cfg_dout3330,
   input         cfg_dout3331,
   input         cfg_dout3332,
   input         cfg_dout3333,
   input         cfg_dout3334,
   input         cfg_dout3335,
   input         cfg_dout3336,
   input         cfg_dout3337,
   input         cfg_dout3338,
   input         cfg_dout3339,
   input         cfg_dout3340,
   input         cfg_dout3341,
   input         cfg_dout3342,
   input         cfg_dout3343,
   input         cfg_dout3344,
   input         cfg_dout3345,
   input         cfg_dout3346,
   input         cfg_dout3347,
   input         cfg_dout3348,
   input         cfg_dout3349,
   input         cfg_dout3350,
   input         cfg_dout3351,
   input         cfg_dout3352,
   input         cfg_dout3353,
   input         cfg_dout3354,
   input         cfg_dout3355,
   input         cfg_dout3356,
   input         cfg_dout3357,
   input         cfg_dout3358,
   input         cfg_dout3359,
   input         cfg_dout3360,
   input         cfg_dout3361,
   input         cfg_dout3362,
   input         cfg_dout3363,
   input         cfg_dout3364,
   input         cfg_dout3365,
   input         cfg_dout3366,
   input         cfg_dout3367,
   input         cfg_dout3368,
   input         cfg_dout3369,
   input         cfg_dout3370,
   input         cfg_dout3371,
   input         cfg_dout3372,
   input         cfg_dout3373,
   input         cfg_dout3374,
   input         cfg_dout3375,
   input         cfg_dout3376,
   input         cfg_dout3377,
   input         cfg_dout3378,
   input         cfg_dout3379,
   input         cfg_dout3380,
   input         cfg_dout3381,
   input         cfg_dout3382,
   input         cfg_dout3383,
   input         cfg_dout3384,
   input         cfg_dout3385,
   input         cfg_dout3386,
   input         cfg_dout3387,
   input         cfg_dout3388,
   input         cfg_dout3389,
   input         cfg_dout3390,
   input         cfg_dout3391,
   input         cfg_dout3392,
   input         cfg_dout3393,
   input         cfg_dout3394,
   input         cfg_dout3395,
   input         cfg_dout3396,
   input         cfg_dout3397,
   input         cfg_dout3398,
   input         cfg_dout3399,
   input         cfg_dout3400,
   input         cfg_dout3401,
   input         cfg_dout3402,
   input         cfg_dout3403,
   input         cfg_dout3404,
   input         cfg_dout3405,
   input         cfg_dout3406,
   input         cfg_dout3407,
   input         cfg_dout3408,
   input         cfg_dout3409,
   input         cfg_dout3410,
   input         cfg_dout3411,
   input         cfg_dout3412,
   input         cfg_dout3413,
   input         cfg_dout3414,
   input         cfg_dout3415,
   input         cfg_dout3416,
   input         cfg_dout3417,
   input         cfg_dout3418,
   input         cfg_dout3419,
   input         cfg_dout3420,
   input         cfg_dout3421,
   input         cfg_dout3422,
   input         cfg_dout3423,
   input         cfg_dout3424,
   input         cfg_dout3425,
   input         cfg_dout3426,
   input         cfg_dout3427,
   input         cfg_dout3428,
   input         cfg_dout3429,
   input         cfg_dout3430,
   input         cfg_dout3431,
   input         cfg_dout3432,
   input         cfg_dout3433,
   input         cfg_dout3434,
   input         cfg_dout3435,
   input         cfg_dout3436,
   input         cfg_dout3437,
   input         cfg_dout3438,
   input         cfg_dout3439,
   input         cfg_dout3440,
   input         cfg_dout3441,
   input         cfg_dout3442,
   input         cfg_dout3443,
   input         cfg_dout3444,
   input         cfg_dout3445,
   input         cfg_dout3446,
   input         cfg_dout3447,
   input         cfg_dout3448,
   input         cfg_dout3449,
   input         cfg_dout3450,
   input         cfg_dout3451,
   input         cfg_dout3452,
   input         cfg_dout3453,
   input         cfg_dout3454,
   input         cfg_dout3455,
   input         cfg_dout3456,
   input         cfg_dout3457,
   input         cfg_dout3458,
   input         cfg_dout3459,
   input         cfg_dout3460,
   input         cfg_dout3461,
   input         cfg_dout3462,
   input         cfg_dout3463,
   input         cfg_dout3464,
   input         cfg_dout3465,
   input         cfg_dout3466,
   input         cfg_dout3467,
   input         cfg_dout3468,
   input         cfg_dout3469,
   input         cfg_dout3470,
   input         cfg_dout3471,
   input         cfg_dout3472,
   input         cfg_dout3473,
   input         cfg_dout3474,
   input         cfg_dout3475,
   input         cfg_dout3476,
   input         cfg_dout3477,
   input         cfg_dout3478,
   input         cfg_dout3479,
   input         cfg_dout3480,
   input         cfg_dout3481,
   input         cfg_dout3482,
   input         cfg_dout3483,
   input         cfg_dout3484,
   input         cfg_dout3485,
   input         cfg_dout3486,
   input         cfg_dout3487,
   input         cfg_dout3488,
   input         cfg_dout3489,
   input         cfg_dout3490,
   input         cfg_dout3491,
   input         cfg_dout3492,
   input         cfg_dout3493,
   input         cfg_dout3494,
   input         cfg_dout3495,
   input         cfg_dout3496,
   input         cfg_dout3497,
   input         cfg_dout3498,
   input         cfg_dout3499,
   input         cfg_dout3500,
   input         cfg_dout3501,
   input         cfg_dout3502,
   input         cfg_dout3503,
   input         cfg_dout3504,
   input         cfg_dout3505,
   input         cfg_dout3506,
   input         cfg_dout3507,
   input         cfg_dout3508,
   input         cfg_dout3509,
   input         cfg_dout3510,
   input         cfg_dout3511,
   input         cfg_dout3512,
   input         cfg_dout3513,
   input         cfg_dout3514,
   input         cfg_dout3515,
   input         cfg_dout3516,
   input         cfg_dout3517,
   input         cfg_dout3518,
   input         cfg_dout3519,
   input         cfg_dout3520,
   input         cfg_dout3521,
   input         cfg_dout3522,
   input         cfg_dout3523,
   input         cfg_dout3524,
   input         cfg_dout3525,
   input         cfg_dout3526,
   input         cfg_dout3527,
   input         cfg_dout3528,
   input         cfg_dout3529,
   input         cfg_dout3530,
   input         cfg_dout3531,
   input         cfg_dout3532,
   input         cfg_dout3533,
   input         cfg_dout3534,
   input         cfg_dout3535,
   input         cfg_dout3536,
   input         cfg_dout3537,
   input         cfg_dout3538,
   input         cfg_dout3539,
   input         cfg_dout3540,
   input         cfg_dout3541,
   input         cfg_dout3542,
   input         cfg_dout3543,
   input         cfg_dout3544,
   input         cfg_dout3545,
   input         cfg_dout3546,
   input         cfg_dout3547,
   input         cfg_dout3548,
   input         cfg_dout3549,
   input         cfg_dout3550,
   input         cfg_dout3551,
   input         cfg_dout3552,
   input         cfg_dout3553,
   input         cfg_dout3554,
   input         cfg_dout3555,
   input         cfg_dout3556,
   input         cfg_dout3557,
   input         cfg_dout3558,
   input         cfg_dout3559,
   input         cfg_dout3560,
   input         cfg_dout3561,
   input         cfg_dout3562,
   input         cfg_dout3563,
   input         cfg_dout3564,
   input         cfg_dout3565,
   input         cfg_dout3566,
   input         cfg_dout3567,
   input         cfg_dout3568,
   input         cfg_dout3569,
   input         cfg_dout3570,
   input         cfg_dout3571,
   input         cfg_dout3572,
   input         cfg_dout3573,
   input         cfg_dout3574,
   input         cfg_dout3575,
   input         cfg_dout3576,
   input         cfg_dout3577,
   input         cfg_dout3578,
   input         cfg_dout3579,
   input         cfg_dout3580,
   input         cfg_dout3581,
   input         cfg_dout3582,
   input         cfg_dout3583,
   input         cfg_dout3584,
   input         cfg_dout3585,
   input         cfg_dout3586,
   input         cfg_dout3587,
   input         cfg_dout3588,
   input         cfg_dout3589,
   input         cfg_dout3590,
   input         cfg_dout3591,
   input         cfg_dout3592,
   input         cfg_dout3593,
   input         cfg_dout3594,
   input         cfg_dout3595,
   input         cfg_dout3596,
   input         cfg_dout3597,
   input         cfg_dout3598,
   input         cfg_dout3599,
   input         cfg_dout3600,
   input         cfg_dout3601,
   input         cfg_dout3602,
   input         cfg_dout3603,
   input         cfg_dout3604,
   input         cfg_dout3605,
   input         cfg_dout3606,
   input         cfg_dout3607,
   input         cfg_dout3608,
   input         cfg_dout3609,
   input         cfg_dout3610,
   input         cfg_dout3611,
   input         cfg_dout3612,
   input         cfg_dout3613,
   input         cfg_dout3614,
   input         cfg_dout3615,
   input         cfg_dout3616,
   input         cfg_dout3617,
   input         cfg_dout3618,
   input         cfg_dout3619,
   input         cfg_dout3620,
   input         cfg_dout3621,
   input         cfg_dout3622,
   input         cfg_dout3623,
   input         cfg_dout3624,
   input         cfg_dout3625,
   input         cfg_dout3626,
   input         cfg_dout3627,
   input         cfg_dout3628,
   input         cfg_dout3629,
   input         cfg_dout3630,
   input         cfg_dout3631,
   input         cfg_dout3632,
   input         cfg_dout3633,
   input         cfg_dout3634,
   input         cfg_dout3635,
   input         cfg_dout3636,
   input         cfg_dout3637,
   input         cfg_dout3638,
   input         cfg_dout3639,
   input         cfg_dout3640,
   input         cfg_dout3641,
   input         cfg_dout3642,
   input         cfg_dout3643,
   input         cfg_dout3644,
   input         cfg_dout3645,
   input         cfg_dout3646,
   input         cfg_dout3647,
   input         cfg_dout3648,
   input         cfg_dout3649,
   input         cfg_dout3650,
   input         cfg_dout3651,
   input         cfg_dout3652,
   input         cfg_dout3653,
   input         cfg_dout3654,
   input         cfg_dout3655,
   input         cfg_dout3656,
   input         cfg_dout3657,
   input         cfg_dout3658,
   input         cfg_dout3659,
   input         cfg_dout3660,
   input         cfg_dout3661,
   input         cfg_dout3662,
   input         cfg_dout3663,
   input         cfg_dout3664,
   input         cfg_dout3665,
   input         cfg_dout3666,
   input         cfg_dout3667,
   input         cfg_dout3668,
   input         cfg_dout3669,
   input         cfg_dout3670,
   input         cfg_dout3671,
   input         cfg_dout3672,
   input         cfg_dout3673,
   input         cfg_dout3674,
   input         cfg_dout3675,
   input         cfg_dout3676,
   input         cfg_dout3677,
   input         cfg_dout3678,
   input         cfg_dout3679,
   input         cfg_dout3680,
   input         cfg_dout3681,
   input         cfg_dout3682,
   input         cfg_dout3683,
   input         cfg_dout3684,
   input         cfg_dout3685,
   input         cfg_dout3686,
   input         cfg_dout3687,
   input         cfg_dout3688,
   input         cfg_dout3689,
   input         cfg_dout3690,
   input         cfg_dout3691,
   input         cfg_dout3692,
   input         cfg_dout3693,
   input         cfg_dout3694,
   input         cfg_dout3695,
   input         cfg_dout3696,
   input         cfg_dout3697,
   input         cfg_dout3698,
   input         cfg_dout3699,
   input         cfg_dout3700,
   input         cfg_dout3701,
   input         cfg_dout3702,
   input         cfg_dout3703,
   input         cfg_dout3704,
   input         cfg_dout3705,
   input         cfg_dout3706,
   input         cfg_dout3707,
   input         cfg_dout3708,
   input         cfg_dout3709,
   input         cfg_dout3710,
   input         cfg_dout3711,
   input         cfg_dout3712,
   input         cfg_dout3713,
   input         cfg_dout3714,
   input         cfg_dout3715,
   input         cfg_dout3716,
   input         cfg_dout3717,
   input         cfg_dout3718,
   input         cfg_dout3719,
   input         cfg_dout3720,
   input         cfg_dout3721,
   input         cfg_dout3722,
   input         cfg_dout3723,
   input         cfg_dout3724,
   input         cfg_dout3725,
   input         cfg_dout3726,
   input         cfg_dout3727,
   input         cfg_dout3728,
   input         cfg_dout3729,
   input         cfg_dout3730,
   input         cfg_dout3731,
   input         cfg_dout3732,
   input         cfg_dout3733,
   input         cfg_dout3734,
   input         cfg_dout3735,
   input         cfg_dout3736,
   input         cfg_dout3737,
   input         cfg_dout3738,
   input         cfg_dout3739,
   input         cfg_dout3740,
   input         cfg_dout3741,
   input         cfg_dout3742,
   input         cfg_dout3743,
   input         cfg_dout3744,
   input         cfg_dout3745,
   input         cfg_dout3746,
   input         cfg_dout3747,
   input         cfg_dout3748,
   input         cfg_dout3749,
   input         cfg_dout3750,
   input         cfg_dout3751,
   input         cfg_dout3752,
   input         cfg_dout3753,
   input         cfg_dout3754,
   input         cfg_dout3755,
   input         cfg_dout3756,
   input         cfg_dout3757,
   input         cfg_dout3758,
   input         cfg_dout3759,
   input         cfg_dout3760,
   input         cfg_dout3761,
   input         cfg_dout3762,
   input         cfg_dout3763,
   input         cfg_dout3764,
   input         cfg_dout3765,
   input         cfg_dout3766,
   input         cfg_dout3767,
   input         cfg_dout3768,
   input         cfg_dout3769,
   input         cfg_dout3770,
   input         cfg_dout3771,
   input         cfg_dout3772,
   input         cfg_dout3773,
   input         cfg_dout3774,
   input         cfg_dout3775,
   input         cfg_dout3776,
   input         cfg_dout3777,
   input         cfg_dout3778,
   input         cfg_dout3779,
   input         cfg_dout3780,
   input         cfg_dout3781,
   input         cfg_dout3782,
   input         cfg_dout3783,
   input         cfg_dout3784,
   input         cfg_dout3785,
   input         cfg_dout3786,
   input         cfg_dout3787,
   input         cfg_dout3788,
   input         cfg_dout3789,
   input         cfg_dout3790,
   input         cfg_dout3791,
   input         cfg_dout3792,
   input         cfg_dout3793,
   input         cfg_dout3794,
   input         cfg_dout3795,
   input         cfg_dout3796,
   input         cfg_dout3797,
   input         cfg_dout3798,
   input         cfg_dout3799,
   input         cfg_dout3800,
   input         cfg_dout3801,
   input         cfg_dout3802,
   input         cfg_dout3803,
   input         cfg_dout3804,
   input         cfg_dout3805,
   input         cfg_dout3806,
   input         cfg_dout3807,
   input         cfg_dout3808,
   input         cfg_dout3809,
   input         cfg_dout3810,
   input         cfg_dout3811,
   input         cfg_dout3812,
   input         cfg_dout3813,
   input         cfg_dout3814,
   input         cfg_dout3815,
   input         cfg_dout3816,
   input         cfg_dout3817,
   input         cfg_dout3818,
   input         cfg_dout3819,
   input         cfg_dout3820,
   input         cfg_dout3821,
   input         cfg_dout3822,
   input         cfg_dout3823,
   input         cfg_dout3824,
   input         cfg_dout3825,
   input         cfg_dout3826,
   input         cfg_dout3827,
   input         cfg_dout3828,
   input         cfg_dout3829,
   input         cfg_dout3830,
   input         cfg_dout3831,
   input         cfg_dout3832,
   input         cfg_dout3833,
   input         cfg_dout3834,
   input         cfg_dout3835,
   input         cfg_dout3836,
   input         cfg_dout3837,
   input         cfg_dout3838,
   input         cfg_dout3839,
   input         cfg_dout3840,
   input         cfg_dout3841,
   input         cfg_dout3842,
   input         cfg_dout3843,
   input         cfg_dout3844,
   input         cfg_dout3845,
   input         cfg_dout3846,
   input         cfg_dout3847,
   input         cfg_dout3848,
   input         cfg_dout3849,
   input         cfg_dout3850,
   input         cfg_dout3851,
   input         cfg_dout3852,
   input         cfg_dout3853,
   input         cfg_dout3854,
   input         cfg_dout3855,
   input         cfg_dout3856,
   input         cfg_dout3857,
   input         cfg_dout3858,
   input         cfg_dout3859,
   input         cfg_dout3860,
   input         cfg_dout3861,
   input         cfg_dout3862,
   input         cfg_dout3863,
   input         cfg_dout3864,
   input         cfg_dout3865,
   input         cfg_dout3866,
   input         cfg_dout3867,
   input         cfg_dout3868,
   input         cfg_dout3869,
   input         cfg_dout3870,
   input         cfg_dout3871,
   input         cfg_dout3872,
   input         cfg_dout3873,
   input         cfg_dout3874,
   input         cfg_dout3875,
   input         cfg_dout3876,
   input         cfg_dout3877,
   input         cfg_dout3878,
   input         cfg_dout3879,
   input         cfg_dout3880,
   input         cfg_dout3881,
   input         cfg_dout3882,
   input         cfg_dout3883,
   input         cfg_dout3884,
   input         cfg_dout3885,
   input         cfg_dout3886,
   input         cfg_dout3887,
   input         cfg_dout3888,
   input         cfg_dout3889,
   input         cfg_dout3890,
   input         cfg_dout3891,
   input         cfg_dout3892,
   input         cfg_dout3893,
   input         cfg_dout3894,
   input         cfg_dout3895,
   input         cfg_dout3896,
   input         cfg_dout3897,
   input         cfg_dout3898,
   input         cfg_dout3899,
   input         cfg_dout3900,
   input         cfg_dout3901,
   input         cfg_dout3902,
   input         cfg_dout3903,
   input         cfg_dout3904,
   input         cfg_dout3905,
   input         cfg_dout3906,
   input         cfg_dout3907,
   input         cfg_dout3908,
   input         cfg_dout3909,
   input         cfg_dout3910,
   input         cfg_dout3911,
   input         cfg_dout3912,
   input         cfg_dout3913,
   input         cfg_dout3914,
   input         cfg_dout3915,
   input         cfg_dout3916,
   input         cfg_dout3917,
   input         cfg_dout3918,
   input         cfg_dout3919,
   input         cfg_dout3920,
   input         cfg_dout3921,
   input         cfg_dout3922,
   input         cfg_dout3923,
   input         cfg_dout3924,
   input         cfg_dout3925,
   input         cfg_dout3926,
   input         cfg_dout3927,
   input         cfg_dout3928,
   input         cfg_dout3929,
   input         cfg_dout3930,
   input         cfg_dout3931,
   input         cfg_dout3932,
   input         cfg_dout3933,
   input         cfg_dout3934,
   input         cfg_dout3935,
   input         cfg_dout3936,
   input         cfg_dout3937,
   input         cfg_dout3938,
   input         cfg_dout3939,
   input         cfg_dout3940,
   input         cfg_dout3941,
   input         cfg_dout3942,
   input         cfg_dout3943,
   input         cfg_dout3944,
   input         cfg_dout3945,
   input         cfg_dout3946,
   input         cfg_dout3947,
   input         cfg_dout3948,
   input         cfg_dout3949,
   input         cfg_dout3950,
   input         cfg_dout3951,
   input         cfg_dout3952,
   input         cfg_dout3953,
   input         cfg_dout3954,
   input         cfg_dout3955,
   input         cfg_dout3956,
   input         cfg_dout3957,
   input         cfg_dout3958,
   input         cfg_dout3959,
   input         cfg_dout3960,
   input         cfg_dout3961,
   input         cfg_dout3962,
   input         cfg_dout3963,
   input         cfg_dout3964,
   input         cfg_dout3965,
   input         cfg_dout3966,
   input         cfg_dout3967,
   input         cfg_dout3968,
   input         cfg_dout3969,
   input         cfg_dout3970,
   input         cfg_dout3971,
   input         cfg_dout3972,
   input         cfg_dout3973,
   input         cfg_dout3974,
   input         cfg_dout3975,
   input         cfg_dout3976,
   input         cfg_dout3977,
   input         cfg_dout3978,
   input         cfg_dout3979,
   input         cfg_dout3980,
   input         cfg_dout3981,
   input         cfg_dout3982,
   input         cfg_dout3983,
   input         cfg_dout3984,
   input         cfg_dout3985,
   input         cfg_dout3986,
   input         cfg_dout3987,
   input         cfg_dout3988,
   input         cfg_dout3989,
   input         cfg_dout3990,
   input         cfg_dout3991,
   input         cfg_dout3992,
   input         cfg_dout3993,
   input         cfg_dout3994,
   input         cfg_dout3995,
   input         cfg_dout3996,
   input         cfg_dout3997,
   input         cfg_dout3998,
   input         cfg_dout3999,
   input         cfg_dout4000,
   input         cfg_dout4001,
   input         cfg_dout4002,
   input         cfg_dout4003,
   input         cfg_dout4004,
   input         cfg_dout4005,
   input         cfg_dout4006,
   input         cfg_dout4007,
   input         cfg_dout4008,
   input         cfg_dout4009,
   input         cfg_dout4010,
   input         cfg_dout4011,
   input         cfg_dout4012,
   input         cfg_dout4013,
   input         cfg_dout4014,
   input         cfg_dout4015,
   input         cfg_dout4016,
   input         cfg_dout4017,
   input         cfg_dout4018,
   input         cfg_dout4019,
   input         cfg_dout4020,
   input         cfg_dout4021,
   input         cfg_dout4022,
   input         cfg_dout4023,
   input         cfg_dout4024,
   input         cfg_dout4025,
   input         cfg_dout4026,
   input         cfg_dout4027,
   input         cfg_dout4028,
   input         cfg_dout4029,
   input         cfg_dout4030,
   input         cfg_dout4031,
   input         cfg_dout4032,
   input         cfg_dout4033,
   input         cfg_dout4034,
   input         cfg_dout4035,
   input         cfg_dout4036,
   input         cfg_dout4037,
   input         cfg_dout4038,
   input         cfg_dout4039,
   input         cfg_dout4040,
   input         cfg_dout4041,
   input         cfg_dout4042,
   input         cfg_dout4043,
   input         cfg_dout4044,
   input         cfg_dout4045,
   input         cfg_dout4046,
   input         cfg_dout4047,
   input         cfg_dout4048,
   input         cfg_dout4049,
   input         cfg_dout4050,
   input         cfg_dout4051,
   input         cfg_dout4052,
   input         cfg_dout4053,
   input         cfg_dout4054,
   input         cfg_dout4055,
   input         cfg_dout4056,
   input         cfg_dout4057,
   input         cfg_dout4058,
   input         cfg_dout4059,
   input         cfg_dout4060,
   input         cfg_dout4061,
   input         cfg_dout4062,
   input         cfg_dout4063,
   input         cfg_dout4064,
   input         cfg_dout4065,
   input         cfg_dout4066,
   input         cfg_dout4067,
   input         cfg_dout4068,
   input         cfg_dout4069,
   input         cfg_dout4070,
   input         cfg_dout4071,
   input         cfg_dout4072,
   input         cfg_dout4073,
   input         cfg_dout4074,
   input         cfg_dout4075,
   input         cfg_dout4076,
   input         cfg_dout4077,
   input         cfg_dout4078,
   input         cfg_dout4079,
   input         cfg_dout4080,
   input         cfg_dout4081,
   input         cfg_dout4082,
   input         cfg_dout4083,
   input         cfg_dout4084,
   input         cfg_dout4085,
   input         cfg_dout4086,
   input         cfg_dout4087,
   input         cfg_dout4088,
   input         cfg_dout4089,
   input         cfg_dout4090,
   input         cfg_dout4091,
   input         cfg_dout4092,
   input         cfg_dout4093,
   input         cfg_dout4094,
   input         cfg_dout4095,
   input         cfg_dout4096,
   input         cfg_dout4097,
   input         cfg_dout4098,
   input         cfg_dout4099,
   input         cfg_dout4100,
   input         cfg_dout4101,
   input         cfg_dout4102,
   input         cfg_dout4103,
   input         cfg_dout4104,
   input         cfg_dout4105,
   input         cfg_dout4106,
   input         cfg_dout4107,
   input         cfg_dout4108,
   input         cfg_dout4109,
   input         cfg_dout4110,
   input         cfg_dout4111,
   input         cfg_dout4112,
   input         cfg_dout4113,
   input         cfg_dout4114,
   input         cfg_dout4115,
   input         cfg_dout4116,
   input         cfg_dout4117,
   input         cfg_dout4118,
   input         cfg_dout4119,
   input         cfg_dout4120,
   input         cfg_dout4121,
   input         cfg_dout4122,
   input         cfg_dout4123,
   input         cfg_dout4124,
   input         cfg_dout4125,
   input         cfg_dout4126,
   input         cfg_dout4127,
   input         cfg_dout4128,
   input         cfg_dout4129,
   input         cfg_dout4130,
   input         cfg_dout4131,
   input         cfg_dout4132,
   input         cfg_dout4133,
   input         cfg_dout4134,
   input         cfg_dout4135,
   input         cfg_dout4136,
   input         cfg_dout4137,
   input         cfg_dout4138,
   input         cfg_dout4139,
   input         cfg_dout4140,
   input         cfg_dout4141,
   input         cfg_dout4142,
   input         cfg_dout4143,
   input         cfg_dout4144,
   input         cfg_dout4145,
   input         cfg_dout4146,
   input         cfg_dout4147,
   input         cfg_dout4148,
   input         cfg_dout4149,
   input         cfg_dout4150,
   input         cfg_dout4151,
   input         cfg_dout4152,
   input         cfg_dout4153,
   input         cfg_dout4154,
   input         cfg_dout4155,
   input         cfg_dout4156,
   input         cfg_dout4157,
   input         cfg_dout4158,
   input         cfg_dout4159,
   input         cfg_dout4160,
   input         cfg_dout4161,
   input         cfg_dout4162,
   input         cfg_dout4163,
   input         cfg_dout4164,
   input         cfg_dout4165,
   input         cfg_dout4166,
   input         cfg_dout4167,
   input         cfg_dout4168,
   input         cfg_dout4169,
   input         cfg_dout4170,
   input         cfg_dout4171,
   input         cfg_dout4172,
   input         cfg_dout4173,
   input         cfg_dout4174,
   input         cfg_dout4175,
   input         cfg_dout4176,
   input         cfg_dout4177,
   input         cfg_dout4178,
   input         cfg_dout4179,
   input         cfg_dout4180,
   input         cfg_dout4181,
   input         cfg_dout4182,
   input         cfg_dout4183,
   input         cfg_dout4184,
   input         cfg_dout4185,
   input         cfg_dout4186,
   input         cfg_dout4187,
   input         cfg_dout4188,
   input         cfg_dout4189,
   input         cfg_dout4190,
   input         cfg_dout4191,
   input         cfg_dout4192,
   input         cfg_dout4193,
   input         cfg_dout4194,
   input         cfg_dout4195,
   input         cfg_dout4196,
   input         cfg_dout4197,
   input         cfg_dout4198,
   input         cfg_dout4199,
   input         cfg_dout4200,
   input         cfg_dout4201,
   input         cfg_dout4202,
   input         cfg_dout4203,
   input         cfg_dout4204,
   input         cfg_dout4205,
   input         cfg_dout4206,
   input         cfg_dout4207,
   input         cfg_dout4208,
   input         cfg_dout4209,
   input         cfg_dout4210,
   input         cfg_dout4211,
   input         cfg_dout4212,
   input         cfg_dout4213,
   input         cfg_dout4214,
   input         cfg_dout4215,
   input         cfg_dout4216,
   input         cfg_dout4217,
   input         cfg_dout4218,
   input         cfg_dout4219,
   input         cfg_dout4220,
   input         cfg_dout4221,
   input         cfg_dout4222,
   input         cfg_dout4223,
   input         cfg_dout4224,
   input         cfg_dout4225,
   input         cfg_dout4226,
   input         cfg_dout4227,
   input         cfg_dout4228,
   input         cfg_dout4229,
   input         cfg_dout4230,
   input         cfg_dout4231,
   input         cfg_dout4232,
   input         cfg_dout4233,
   input         cfg_dout4234,
   input         cfg_dout4235,
   input         cfg_dout4236,
   input         cfg_dout4237,
   input         cfg_dout4238,
   input         cfg_dout4239,
   input         cfg_dout4240,
   input         cfg_dout4241,
   input         cfg_dout4242,
   input         cfg_dout4243,
   input         cfg_dout4244,
   input         cfg_dout4245,
   input         cfg_dout4246,
   input         cfg_dout4247,
   input         cfg_dout4248,
   input         cfg_dout4249,
   input         cfg_dout4250,
   input         cfg_dout4251,
   input         cfg_dout4252,
   input         cfg_dout4253,
   input         cfg_dout4254,
   input         cfg_dout4255,
   input         cfg_dout4256,
   input         cfg_dout4257,
   input         cfg_dout4258,
   input         cfg_dout4259,
   input         cfg_dout4260,
   input         cfg_dout4261,
   input         cfg_dout4262,
   input         cfg_dout4263,
   input         cfg_dout4264,
   input         cfg_dout4265,
   input         cfg_dout4266,
   input         cfg_dout4267,
   input         cfg_dout4268,
   input         cfg_dout4269,
   input         cfg_dout4270,
   input         cfg_dout4271,
   input         cfg_dout4272,
   input         cfg_dout4273,
   input         cfg_dout4274,
   input         cfg_dout4275,
   input         cfg_dout4276,
   input         cfg_dout4277,
   input         cfg_dout4278,
   input         cfg_dout4279,
   input         cfg_dout4280,
   input         cfg_dout4281,
   input         cfg_dout4282,
   input         cfg_dout4283,
   input         cfg_dout4284,
   input         cfg_dout4285,
   input         cfg_dout4286,
   input         cfg_dout4287,
   input         cfg_dout4288,
   input         cfg_dout4289,
   input         cfg_dout4290,
   input         cfg_dout4291,
   input         cfg_dout4292,
   input         cfg_dout4293,
   input         cfg_dout4294,
   input         cfg_dout4295,
   input         cfg_dout4296,
   input         cfg_dout4297,
   input         cfg_dout4298,
   input         cfg_dout4299,
   input         cfg_dout4300,
   input         cfg_dout4301,
   input         cfg_dout4302,
   input         cfg_dout4303,
   input         cfg_dout4304,
   input         cfg_dout4305,
   input         cfg_dout4306,
   input         cfg_dout4307,
   input         cfg_dout4308,
   input         cfg_dout4309,
   input         cfg_dout4310,
   input         cfg_dout4311,
   input         cfg_dout4312,
   input         cfg_dout4313,
   input         cfg_dout4314,
   input         cfg_dout4315,
   input         cfg_dout4316,
   input         cfg_dout4317,
   input         cfg_dout4318,
   input         cfg_dout4319,
   input         cfg_dout4320,
   input         cfg_dout4321,
   input         cfg_dout4322,
   input         cfg_dout4323,
   input         cfg_dout4324,
   input         cfg_dout4325,
   input         cfg_dout4326,
   input         cfg_dout4327,
   input         cfg_dout4328,
   input         cfg_dout4329,
   input         cfg_dout4330,
   input         cfg_dout4331,
   input         cfg_dout4332,
   input         cfg_dout4333,
   input         cfg_dout4334,
   input         cfg_dout4335,
   input         cfg_dout4336,
   input         cfg_dout4337,
   input         cfg_dout4338,
   input         cfg_dout4339,
   input         cfg_dout4340,
   input         cfg_dout4341,
   input         cfg_dout4342,
   input         cfg_dout4343,
   input         cfg_dout4344,
   input         cfg_dout4345,
   input         cfg_dout4346,
   input         cfg_dout4347,
   input         cfg_dout4348,
   input         cfg_dout4349,
   input         cfg_dout4350,
   input         cfg_dout4351,
   input         cfg_dout4352,
   input         cfg_dout4353,
   input         cfg_dout4354,
   input         cfg_dout4355,
   input         cfg_dout4356,
   input         cfg_dout4357,
   input         cfg_dout4358,
   input         cfg_dout4359,
   input         cfg_dout4360,
   input         cfg_dout4361,
   input         cfg_dout4362,
   input         cfg_dout4363,
   input         cfg_dout4364,
   input         cfg_dout4365,
   input         cfg_dout4366,
   input         cfg_dout4367,
   input         cfg_dout4368,
   input         cfg_dout4369,
   input         cfg_dout4370,
   input         cfg_dout4371,
   input         cfg_dout4372,
   input         cfg_dout4373,
   input         cfg_dout4374,
   input         cfg_dout4375,
   input         cfg_dout4376,
   input         cfg_dout4377,
   input         cfg_dout4378,
   input         cfg_dout4379,
   input         cfg_dout4380,
   input         cfg_dout4381,
   input         cfg_dout4382,
   input         cfg_dout4383,
   input         cfg_dout4384,
   input         cfg_dout4385,
   input         cfg_dout4386,
   input         cfg_dout4387,
   input         cfg_dout4388,
   input         cfg_dout4389,
   input         cfg_dout4390,
   input         cfg_dout4391,
   input         cfg_dout4392,
   input         cfg_dout4393,
   input         cfg_dout4394,
   input         cfg_dout4395,
   input         cfg_dout4396,
   input         cfg_dout4397,
   input         cfg_dout4398,
   input         cfg_dout4399,
   input         cfg_dout4400,
   input         cfg_dout4401,
   input         cfg_dout4402,
   input         cfg_dout4403,
   input         cfg_dout4404,
   input         cfg_dout4405,
   input         cfg_dout4406,
   input         cfg_dout4407,
   input         cfg_dout4408,
   input         cfg_dout4409,
   input         cfg_dout4410,
   input         cfg_dout4411,
   input         cfg_dout4412,
   input         cfg_dout4413,
   input         cfg_dout4414,
   input         cfg_dout4415,
   input         cfg_dout4416,
   input         cfg_dout4417,
   input         cfg_dout4418,
   input         cfg_dout4419,
   input         cfg_dout4420,
   input         cfg_dout4421,
   input         cfg_dout4422,
   input         cfg_dout4423,
   input         cfg_dout4424,
   input         cfg_dout4425,
   input         cfg_dout4426,
   input         cfg_dout4427,
   input         cfg_dout4428,
   input         cfg_dout4429,
   input         cfg_dout4430,
   input         cfg_dout4431,
   input         cfg_dout4432,
   input         cfg_dout4433,
   input         cfg_dout4434,
   input         cfg_dout4435,
   input         cfg_dout4436,
   input         cfg_dout4437,
   input         cfg_dout4438,
   input         cfg_dout4439,
   input         cfg_dout4440,
   input         cfg_dout4441,
   input         cfg_dout4442,
   input         cfg_dout4443,
   input         cfg_dout4444,
   input         cfg_dout4445,
   input         cfg_dout4446,
   input         cfg_dout4447,
   input         cfg_dout4448,
   input         cfg_dout4449,
   input         cfg_dout4450,
   input         cfg_dout4451,
   input         cfg_dout4452,
   input         cfg_dout4453,
   input         cfg_dout4454,
   input         cfg_dout4455,
   input         cfg_dout4456,
   input         cfg_dout4457,
   input         cfg_dout4458,
   input         cfg_dout4459,
   input         cfg_dout4460,
   input         cfg_dout4461,
   input         cfg_dout4462,
   input         cfg_dout4463,
   input         cfg_dout4464,
   input         cfg_dout4465,
   input         cfg_dout4466,
   input         cfg_dout4467,
   input         cfg_dout4468,
   input         cfg_dout4469,
   input         cfg_dout4470,
   input         cfg_dout4471,
   input         cfg_dout4472,
   input         cfg_dout4473,
   input         cfg_dout4474,
   input         cfg_dout4475,
   input         cfg_dout4476,
   input         cfg_dout4477,
   input         cfg_dout4478,
   input         cfg_dout4479,
   input         cfg_dout4480,
   input         cfg_dout4481,
   input         cfg_dout4482,
   input         cfg_dout4483,
   input         cfg_dout4484,
   input         cfg_dout4485,
   input         cfg_dout4486,
   input         cfg_dout4487,
   input         cfg_dout4488,
   input         cfg_dout4489,
   input         cfg_dout4490,
   input         cfg_dout4491,
   input         cfg_dout4492,
   input         cfg_dout4493,
   input         cfg_dout4494,
   input         cfg_dout4495,
   input         cfg_dout4496,
   input         cfg_dout4497,
   input         cfg_dout4498,
   input         cfg_dout4499,
   input         cfg_dout4500,
   input         cfg_dout4501,
   input         cfg_dout4502,
   input         cfg_dout4503,
   input         cfg_dout4504,
   input         cfg_dout4505,
   input         cfg_dout4506,
   input         cfg_dout4507,
   input         cfg_dout4508,
   input         cfg_dout4509,
   input         cfg_dout4510,
   input         cfg_dout4511,
   input         cfg_dout4512,
   input         cfg_dout4513,
   input         cfg_dout4514,
   input         cfg_dout4515,
   input         cfg_dout4516,
   input         cfg_dout4517,
   input         cfg_dout4518,
   input         cfg_dout4519,
   input         cfg_dout4520,
   input         cfg_dout4521,
   input         cfg_dout4522,
   input         cfg_dout4523,
   input         cfg_dout4524,
   input         cfg_dout4525,
   input         cfg_dout4526,
   input         cfg_dout4527,
   input         cfg_dout4528,
   input         cfg_dout4529,
   input         cfg_dout4530,
   input         cfg_dout4531,
   input         cfg_dout4532,
   input         cfg_dout4533,
   input         cfg_dout4534,
   input         cfg_dout4535,
   input         cfg_dout4536,
   input         cfg_dout4537,
   input         cfg_dout4538,
   input         cfg_dout4539,
   input         cfg_dout4540,
   input         cfg_dout4541,
   input         cfg_dout4542,
   input         cfg_dout4543,
   input         cfg_dout4544,
   input         cfg_dout4545,
   input         cfg_dout4546,
   input         cfg_dout4547,
   input         cfg_dout4548,
   input         cfg_dout4549,
   input         cfg_dout4550,
   input         cfg_dout4551,
   input         cfg_dout4552,
   input         cfg_dout4553,
   input         cfg_dout4554,
   input         cfg_dout4555,
   input         cfg_dout4556,
   input         cfg_dout4557,
   input         cfg_dout4558,
   input         cfg_dout4559,
   input         cfg_dout4560,
   input         cfg_dout4561,
   input         cfg_dout4562,
   input         cfg_dout4563,
   input         cfg_dout4564,
   input         cfg_dout4565,
   input         cfg_dout4566,
   input         cfg_dout4567,
   input         cfg_dout4568,
   input         cfg_dout4569,
   input         cfg_dout4570,
   input         cfg_dout4571,
   input         cfg_dout4572,
   input         cfg_dout4573,
   input         cfg_dout4574,
   input         cfg_dout4575,
   input         cfg_dout4576,
   input         cfg_dout4577,
   input         cfg_dout4578,
   input         cfg_dout4579,
   input         cfg_dout4580,
   input         cfg_dout4581,
   input         cfg_dout4582,
   input         cfg_dout4583,
   input         cfg_dout4584,
   input         cfg_dout4585,
   input         cfg_dout4586,
   input         cfg_dout4587,
   input         cfg_dout4588,
   input         cfg_dout4589,
   input         cfg_dout4590,
   input         cfg_dout4591,
   input         cfg_dout4592,
   input         cfg_dout4593,
   input         cfg_dout4594,
   input         cfg_dout4595,
   input         cfg_dout4596,
   input         cfg_dout4597,
   input         cfg_dout4598,
   input         cfg_dout4599,
   input         cfg_dout4600,
   input         cfg_dout4601,
   input         cfg_dout4602,
   input         cfg_dout4603,
   input         cfg_dout4604,
   input         cfg_dout4605,
   input         cfg_dout4606,
   input         cfg_dout4607,
   input         cfg_dout4608,
   input         cfg_dout4609,
   input         cfg_dout4610,
   input         cfg_dout4611,
   input         cfg_dout4612,
   input         cfg_dout4613,
   input         cfg_dout4614,
   input         cfg_dout4615,
   input         cfg_dout4616,
   input         cfg_dout4617,
   input         cfg_dout4618,
   input         cfg_dout4619,
   input         cfg_dout4620,
   input         cfg_dout4621,
   input         cfg_dout4622,
   input         cfg_dout4623,
   input         cfg_dout4624,
   input         cfg_dout4625,
   input         cfg_dout4626,
   input         cfg_dout4627,
   input         cfg_dout4628,
   input         cfg_dout4629,
   input         cfg_dout4630,
   input         cfg_dout4631,
   input         cfg_dout4632,
   input         cfg_dout4633,
   input         cfg_dout4634,
   input         cfg_dout4635,
   input         cfg_dout4636,
   input         cfg_dout4637,
   input         cfg_dout4638,
   input         cfg_dout4639,
   input         cfg_dout4640,
   input         cfg_dout4641,
   input         cfg_dout4642,
   input         cfg_dout4643,
   input         cfg_dout4644,
   input         cfg_dout4645,
   input         cfg_dout4646,
   input         cfg_dout4647,
   input         cfg_dout4648,
   input         cfg_dout4649,
   input         cfg_dout4650,
   input         cfg_dout4651,
   input         cfg_dout4652,
   input         cfg_dout4653,
   input         cfg_dout4654,
   input         cfg_dout4655,
   input         cfg_dout4656,
   input         cfg_dout4657,
   input         cfg_dout4658,
   input         cfg_dout4659,
   input         cfg_dout4660,
   input         cfg_dout4661,
   input         cfg_dout4662,
   input         cfg_dout4663,
   input         cfg_dout4664,
   input         cfg_dout4665,
   input         cfg_dout4666,
   input         cfg_dout4667,
   input         cfg_dout4668,
   input         cfg_dout4669,
   input         cfg_dout4670,
   input         cfg_dout4671,
   input         cfg_dout4672,
   input         cfg_dout4673,
   input         cfg_dout4674,
   input         cfg_dout4675,
   input         cfg_dout4676,
   input         cfg_dout4677,
   input         cfg_dout4678,
   input         cfg_dout4679,
   input         cfg_dout4680,
   input         cfg_dout4681,
   input         cfg_dout4682,
   input         cfg_dout4683,
   input         cfg_dout4684,
   input         cfg_dout4685,
   input         cfg_dout4686,
   input         cfg_dout4687,
   input         cfg_dout4688,
   input         cfg_dout4689,
   input         cfg_dout4690,
   input         cfg_dout4691,
   input         cfg_dout4692,
   input         cfg_dout4693,
   input         cfg_dout4694,
   input         cfg_dout4695,
   input         cfg_dout4696,
   input         cfg_dout4697,
   input         cfg_dout4698,
   input         cfg_dout4699,
   input         cfg_dout4700,
   input         cfg_dout4701,
   input         cfg_dout4702,
   input         cfg_dout4703,
   input         cfg_dout4704,
   input         cfg_dout4705,
   input         cfg_dout4706,
   input         cfg_dout4707,
   input         cfg_dout4708,
   input         cfg_dout4709,
   input         cfg_dout4710,
   input         cfg_dout4711,
   input         cfg_dout4712,
   input         cfg_dout4713,
   input         cfg_dout4714,
   input         cfg_dout4715,
   input         cfg_dout4716,
   input         cfg_dout4717,
   input         cfg_dout4718,
   input         cfg_dout4719,
   input         cfg_dout4720,
   input         cfg_dout4721,
   input         cfg_dout4722,
   input         cfg_dout4723,
   input         cfg_dout4724,
   input         cfg_dout4725,
   input         cfg_dout4726,
   input         cfg_dout4727,
   input         cfg_dout4728,
   input         cfg_dout4729,
   input         cfg_dout4730,
   input         cfg_dout4731,
   input         cfg_dout4732,
   input         cfg_dout4733,
   input         cfg_dout4734,
   input         cfg_dout4735,
   input         cfg_dout4736,
   input         cfg_dout4737,
   input         cfg_dout4738,
   input         cfg_dout4739,
   input         cfg_dout4740,
   input         cfg_dout4741,
   input         cfg_dout4742,
   input         cfg_dout4743,
   input         cfg_dout4744,
   input         cfg_dout4745,
   input         cfg_dout4746,
   input         cfg_dout4747,
   input         cfg_dout4748,
   input         cfg_dout4749,
   input         cfg_dout4750,
   input         cfg_dout4751,
   input         cfg_dout4752,
   input         cfg_dout4753,
   input         cfg_dout4754,
   input         cfg_dout4755,
   input         cfg_dout4756,
   input         cfg_dout4757,
   input         cfg_dout4758,
   input         cfg_dout4759,
   input         cfg_dout4760,
   input         cfg_dout4761,
   input         cfg_dout4762,
   input         cfg_dout4763,
   input         cfg_dout4764,
   input         cfg_dout4765,
   input         cfg_dout4766,
   input         cfg_dout4767,
   input         cfg_dout4768,
   input         cfg_dout4769,
   input         cfg_dout4770,
   input         cfg_dout4771,
   input         cfg_dout4772,
   input         cfg_dout4773,
   input         cfg_dout4774,
   input         cfg_dout4775,
   input         cfg_dout4776,
   input         cfg_dout4777,
   input         cfg_dout4778,
   input         cfg_dout4779,
   input         cfg_dout4780,
   input         cfg_dout4781,
   input         cfg_dout4782,
   input         cfg_dout4783,
   input         cfg_dout4784,
   input         cfg_dout4785,
   input         cfg_dout4786,
   input         cfg_dout4787,
   input         cfg_dout4788,
   input         cfg_dout4789,
   input         cfg_dout4790,
   input         cfg_dout4791,
   input         cfg_dout4792,
   input         cfg_dout4793,
   input         cfg_dout4794,
   input         cfg_dout4795,
   input         cfg_dout4796,
   input         cfg_dout4797,
   input         cfg_dout4798,
   input         cfg_dout4799,
   input         cfg_dout4800,
   input         cfg_dout4801,
   input         cfg_dout4802,
   input         cfg_dout4803,
   input         cfg_dout4804,
   input         cfg_dout4805,
   input         cfg_dout4806,
   input         cfg_dout4807,
   input         cfg_dout4808,
   input         cfg_dout4809,
   input         cfg_dout4810,
   input         cfg_dout4811,
   input         cfg_dout4812,
   input         cfg_dout4813,
   input         cfg_dout4814,
   input         cfg_dout4815,
   input         cfg_dout4816,
   input         cfg_dout4817,
   input         cfg_dout4818,
   input         cfg_dout4819,
   input         cfg_dout4820,
   input         cfg_dout4821,
   input         cfg_dout4822,
   input         cfg_dout4823,
   input         cfg_dout4824,
   input         cfg_dout4825,
   input         cfg_dout4826,
   input         cfg_dout4827,
   input         cfg_dout4828,
   input         cfg_dout4829,
   input         cfg_dout4830,
   input         cfg_dout4831,
   input         cfg_dout4832,
   input         cfg_dout4833,
   input         cfg_dout4834,
   input         cfg_dout4835,
   input         cfg_dout4836,
   input         cfg_dout4837,
   input         cfg_dout4838,
   input         cfg_dout4839,
   input         cfg_dout4840,
   input         cfg_dout4841,
   input         cfg_dout4842,
   input         cfg_dout4843,
   input         cfg_dout4844,
   input         cfg_dout4845,
   input         cfg_dout4846,
   input         cfg_dout4847,
   input         cfg_dout4848,
   input         cfg_dout4849,
   input         cfg_dout4850,
   input         cfg_dout4851,
   input         cfg_dout4852,
   input         cfg_dout4853,
   input         cfg_dout4854,
   input         cfg_dout4855,
   input         cfg_dout4856,
   input         cfg_dout4857,
   input         cfg_dout4858,
   input         cfg_dout4859,
   input         cfg_dout4860,
   input         cfg_dout4861,
   input         cfg_dout4862,
   input         cfg_dout4863,
   input         cfg_dout4864,
   input         cfg_dout4865,
   input         cfg_dout4866,
   input         cfg_dout4867,
   input         cfg_dout4868,
   input         cfg_dout4869,
   input         cfg_dout4870,
   input         cfg_dout4871,
   input         cfg_dout4872,
   input         cfg_dout4873,
   input         cfg_dout4874,
   input         cfg_dout4875,
   input         cfg_dout4876,
   input         cfg_dout4877,
   input         cfg_dout4878,
   input         cfg_dout4879,
   input         cfg_dout4880,
   input         cfg_dout4881,
   input         cfg_dout4882,
   input         cfg_dout4883,
   input         cfg_dout4884,
   input         cfg_dout4885,
   input         cfg_dout4886,
   input         cfg_dout4887,
   input         cfg_dout4888,
   input         cfg_dout4889,
   input         cfg_dout4890,
   input         cfg_dout4891,
   input         cfg_dout4892,
   input         cfg_dout4893,
   input         cfg_dout4894,
   input         cfg_dout4895,
   input         cfg_dout4896,
   input         cfg_dout4897,
   input         cfg_dout4898,
   input         cfg_dout4899,
   input         cfg_dout4900,
   input         cfg_dout4901,
   input         cfg_dout4902,
   input         cfg_dout4903,
   input         cfg_dout4904,
   input         cfg_dout4905,
   input         cfg_dout4906,
   input         cfg_dout4907,
   input         cfg_dout4908,
   input         cfg_dout4909,
   input         cfg_dout4910,
   input         cfg_dout4911,
   input         cfg_dout4912,
   input         cfg_dout4913,
   input         cfg_dout4914,
   input         cfg_dout4915,
   input         cfg_dout4916,
   input         cfg_dout4917,
   input         cfg_dout4918,
   input         cfg_dout4919,
   input         cfg_dout4920,
   input         cfg_dout4921,
   input         cfg_dout4922,
   input         cfg_dout4923,
   input         cfg_dout4924,
   input         cfg_dout4925,
   input         cfg_dout4926,
   input         cfg_dout4927,
   input         cfg_dout4928,
   input         cfg_dout4929,
   input         cfg_dout4930,
   input         cfg_dout4931,
   input         cfg_dout4932,
   input         cfg_dout4933,
   input         cfg_dout4934,
   input         cfg_dout4935,
   input         cfg_dout4936,
   input         cfg_dout4937,
   input         cfg_dout4938,
   input         cfg_dout4939,
   input         cfg_dout4940,
   input         cfg_dout4941,
   input         cfg_dout4942,
   input         cfg_dout4943,
   input         cfg_dout4944,
   input         cfg_dout4945,
   input         cfg_dout4946,
   input         cfg_dout4947,
   input         cfg_dout4948,
   input         cfg_dout4949,
   input         cfg_dout4950,
   input         cfg_dout4951,
   input         cfg_dout4952,
   input         cfg_dout4953,
   input         cfg_dout4954,
   input         cfg_dout4955,
   input         cfg_dout4956,
   input         cfg_dout4957,
   input         cfg_dout4958,
   input         cfg_dout4959,
   input         cfg_dout4960,
   input         cfg_dout4961,
   input         cfg_dout4962,
   input         cfg_dout4963,
   input         cfg_dout4964,
   input         cfg_dout4965,
   input         cfg_dout4966,
   input         cfg_dout4967,
   input         cfg_dout4968,
   input         cfg_dout4969,
   input         cfg_dout4970,
   input         cfg_dout4971,
   input         cfg_dout4972,
   input         cfg_dout4973,
   input         cfg_dout4974,
   input         cfg_dout4975,
   input         cfg_dout4976,
   input         cfg_dout4977,
   input         cfg_dout4978,
   input         cfg_dout4979,
   input         cfg_dout4980,
   input         cfg_dout4981,
   input         cfg_dout4982,
   input         cfg_dout4983,
   input         cfg_dout4984,
   input         cfg_dout4985,
   input         cfg_dout4986,
   input         cfg_dout4987,
   input         cfg_dout4988,
   input         cfg_dout4989,
   input         cfg_dout4990,
   input         cfg_dout4991,
   input         cfg_dout4992,
   input         cfg_dout4993,
   input         cfg_dout4994,
   input         cfg_dout4995,
   input         cfg_dout4996,
   input         cfg_dout4997,
   input         cfg_dout4998,
   input         cfg_dout4999,
   input         cfg_dout5000,
   input         cfg_dout5001,
   input         cfg_dout5002,
   input         cfg_dout5003,
   input         cfg_dout5004,
   input         cfg_dout5005,
   input         cfg_dout5006,
   input         cfg_dout5007,
   input         cfg_dout5008,
   input         cfg_dout5009,
   input         cfg_dout5010,
   input         cfg_dout5011,
   input         cfg_dout5012,
   input         cfg_dout5013,
   input         cfg_dout5014,
   input         cfg_dout5015,
   input         cfg_dout5016,
   input         cfg_dout5017,
   input         cfg_dout5018,
   input         cfg_dout5019,
   input         cfg_dout5020,
   input         cfg_dout5021,
   input         cfg_dout5022,
   input         cfg_dout5023,
   input         cfg_dout5024,
   input         cfg_dout5025,
   input         cfg_dout5026,
   input         cfg_dout5027,
   input         cfg_dout5028,
   input         cfg_dout5029,
   input         cfg_dout5030,
   input         cfg_dout5031,
   input         cfg_dout5032,
   input         cfg_dout5033,
   input         cfg_dout5034,
   input         cfg_dout5035,
   input         cfg_dout5036,
   input         cfg_dout5037,
   input         cfg_dout5038,
   input         cfg_dout5039,
   input         cfg_dout5040,
   input         cfg_dout5041,
   input         cfg_dout5042,
   input         cfg_dout5043,
   input         cfg_dout5044,
   input         cfg_dout5045,
   input         cfg_dout5046,
   input         cfg_dout5047,
   input         cfg_dout5048,
   input         cfg_dout5049,
   input         cfg_dout5050,
   input         cfg_dout5051,
   input         cfg_dout5052,
   input         cfg_dout5053,
   input         cfg_dout5054,
   input         cfg_dout5055,
   input         cfg_dout5056,
   input         cfg_dout5057,
   input         cfg_dout5058,
   input         cfg_dout5059,
   input         cfg_dout5060,
   input         cfg_dout5061,
   input         cfg_dout5062,
   input         cfg_dout5063,
   input         cfg_dout5064,
   input         cfg_dout5065,
   input         cfg_dout5066,
   input         cfg_dout5067,
   input         cfg_dout5068,
   input         cfg_dout5069,
   input         cfg_dout5070,
   input         cfg_dout5071,
   input         cfg_dout5072,
   input         cfg_dout5073,
   input         cfg_dout5074,
   input         cfg_dout5075,
   input         cfg_dout5076,
   input         cfg_dout5077,
   input         cfg_dout5078,
   input         cfg_dout5079,
   input         cfg_dout5080,
   input         cfg_dout5081,
   input         cfg_dout5082,
   input         cfg_dout5083,
   input         cfg_dout5084,
   input         cfg_dout5085,
   input         cfg_dout5086,
   input         cfg_dout5087,
   input         cfg_dout5088,
   input         cfg_dout5089,
   input         cfg_dout5090,
   input         cfg_dout5091,
   input         cfg_dout5092,
   input         cfg_dout5093,
   input         cfg_dout5094,
   input         cfg_dout5095,
   input         cfg_dout5096,
   input         cfg_dout5097,
   input         cfg_dout5098,
   input         cfg_dout5099,
   input         cfg_dout5100,
   input         cfg_dout5101,
   input         cfg_dout5102,
   input         cfg_dout5103,
   input         cfg_dout5104,
   input         cfg_dout5105,
   input         cfg_dout5106,
   input         cfg_dout5107,
   input         cfg_dout5108,
   input         cfg_dout5109,
   input         cfg_dout5110,
   input         cfg_dout5111,
   input         cfg_dout5112,
   input         cfg_dout5113,
   input         cfg_dout5114,
   input         cfg_dout5115,
   input         cfg_dout5116,
   input         cfg_dout5117,
   input         cfg_dout5118,
   input         cfg_dout5119,
   input         cfg_dout5120,
   input         cfg_dout5121,
   input         cfg_dout5122,
   input         cfg_dout5123,
   input         cfg_dout5124,
   input         cfg_dout5125,
   input         cfg_dout5126,
   input         cfg_dout5127,
   input         cfg_dout5128,
   input         cfg_dout5129,
   input         cfg_dout5130,
   input         cfg_dout5131,
   input         cfg_dout5132,
   input         cfg_dout5133,
   input         cfg_dout5134,
   input         cfg_dout5135,
   input         cfg_dout5136,
   input         cfg_dout5137,
   input         cfg_dout5138,
   input         cfg_dout5139,
   input         cfg_dout5140,
   input         cfg_dout5141,
   input         cfg_dout5142,
   input         cfg_dout5143,
   input         cfg_dout5144,
   input         cfg_dout5145,
   input         cfg_dout5146,
   input         cfg_dout5147,
   input         cfg_dout5148,
   input         cfg_dout5149,
   input         cfg_dout5150,
   input         cfg_dout5151,
   input         cfg_dout5152,
   input         cfg_dout5153,
   input         cfg_dout5154,
   input         cfg_dout5155,
   input         cfg_dout5156,
   input         cfg_dout5157,
   input         cfg_dout5158,
   input         cfg_dout5159,
   input         cfg_dout5160,
   input         cfg_dout5161,
   input         cfg_dout5162,
   input         cfg_dout5163,
   input         cfg_dout5164,
   input         cfg_dout5165,
   input         cfg_dout5166,
   input         cfg_dout5167,
   input         cfg_dout5168,
   input         cfg_dout5169,
   input         cfg_dout5170,
   input         cfg_dout5171,
   input         cfg_dout5172,
   input         cfg_dout5173,
   input         cfg_dout5174,
   input         cfg_dout5175,
   input         cfg_dout5176,
   input         cfg_dout5177,
   input         cfg_dout5178,
   input         cfg_dout5179,
   input         cfg_dout5180,
   input         cfg_dout5181,
   input         cfg_dout5182,
   input         cfg_dout5183,
   input         cfg_dout5184,
   input         cfg_dout5185,
   input         cfg_dout5186,
   input         cfg_dout5187,
   input         cfg_dout5188,
   input         cfg_dout5189,
   input         cfg_dout5190,
   input         cfg_dout5191,
   input         cfg_dout5192,
   input         cfg_dout5193,
   input         cfg_dout5194,
   input         cfg_dout5195,
   input         cfg_dout5196,
   input         cfg_dout5197,
   input         cfg_dout5198,
   input         cfg_dout5199,
   input         cfg_dout5200,
   input         cfg_dout5201,
   input         cfg_dout5202,
   input         cfg_dout5203,
   input         cfg_dout5204,
   input         cfg_dout5205,
   input         cfg_dout5206,
   input         cfg_dout5207,
   input         cfg_dout5208,
   input         cfg_dout5209,
   input         cfg_dout5210,
   input         cfg_dout5211,
   input         cfg_dout5212,
   input         cfg_dout5213,
   input         cfg_dout5214,
   input         cfg_dout5215,
   input         cfg_dout5216,
   input         cfg_dout5217,
   input         cfg_dout5218,
   input         cfg_dout5219,
   input         cfg_dout5220,
   input         cfg_dout5221,
   input         cfg_dout5222,
   input         cfg_dout5223,
   input         cfg_dout5224,
   input         cfg_dout5225,
   input         cfg_dout5226,
   input         cfg_dout5227,
   input         cfg_dout5228,
   input         cfg_dout5229,
   input         cfg_dout5230,
   input         cfg_dout5231,
   input         cfg_dout5232,
   input         cfg_dout5233,
   input         cfg_dout5234,
   input         cfg_dout5235,
   input         cfg_dout5236,
   input         cfg_dout5237,
   input         cfg_dout5238,
   input         cfg_dout5239,
   input         cfg_dout5240,
   input         cfg_dout5241,
   input         cfg_dout5242,
   input         cfg_dout5243,
   input         cfg_dout5244,
   input         cfg_dout5245,
   input         cfg_dout5246,
   input         cfg_dout5247,
   input         cfg_dout5248,
   input         cfg_dout5249,
   input         cfg_dout5250,
   input         cfg_dout5251,
   input         cfg_dout5252,
   input         cfg_dout5253,
   input         cfg_dout5254,
   input         cfg_dout5255,
   input         cfg_dout5256,
   input         cfg_dout5257,
   input         cfg_dout5258,
   input         cfg_dout5259,
   input         cfg_dout5260,
   input         cfg_dout5261,
   input         cfg_dout5262,
   input         cfg_dout5263,
   input         cfg_dout5264,
   input         cfg_dout5265,
   input         cfg_dout5266,
   input         cfg_dout5267,
   input         cfg_dout5268,
   input         cfg_dout5269,
   input         cfg_dout5270,
   input         cfg_dout5271,
   input         cfg_dout5272,
   input         cfg_dout5273,
   input         cfg_dout5274,
   input         cfg_dout5275,
   input         cfg_dout5276,
   input         cfg_dout5277,
   input         cfg_dout5278,
   input         cfg_dout5279,
   input         cfg_dout5280,
   input         cfg_dout5281,
   input         cfg_dout5282,
   input         cfg_dout5283,
   input         cfg_dout5284,
   input         cfg_dout5285,
   input         cfg_dout5286,
   input         cfg_dout5287,
   input         cfg_dout5288,
   input         cfg_dout5289,
   input         cfg_dout5290,
   input         cfg_dout5291,
   input         cfg_dout5292,
   input         cfg_dout5293,
   input         cfg_dout5294,
   input         cfg_dout5295,
   input         cfg_dout5296,
   input         cfg_dout5297,
   input         cfg_dout5298,
   input         cfg_dout5299,
   input         cfg_dout5300,
   input         cfg_dout5301,
   input         cfg_dout5302,
   input         cfg_dout5303,
   input         cfg_dout5304,
   input         cfg_dout5305,
   input         cfg_dout5306,
   input         cfg_dout5307,
   input         cfg_dout5308,
   input         cfg_dout5309,
   input         cfg_dout5310,
   input         cfg_dout5311,
   input         cfg_dout5312,
   input         cfg_dout5313,
   input         cfg_dout5314,
   input         cfg_dout5315,
   input         cfg_dout5316,
   input         cfg_dout5317,
   input         cfg_dout5318,
   input         cfg_dout5319,
   input         cfg_dout5320,
   input         cfg_dout5321,
   input         cfg_dout5322,
   input         cfg_dout5323,
   input         cfg_dout5324,
   input         cfg_dout5325,
   input         cfg_dout5326,
   input         cfg_dout5327,
   input         cfg_dout5328,
   input         cfg_dout5329,
   input         cfg_dout5330,
   input         cfg_dout5331,
   input         cfg_dout5332,
   input         cfg_dout5333,
   input         cfg_dout5334,
   input         cfg_dout5335,
   input         cfg_dout5336,
   input         cfg_dout5337,
   input         cfg_dout5338,
   input         cfg_dout5339,
   input         cfg_dout5340,
   input         cfg_dout5341,
   input         cfg_dout5342,
   input         cfg_dout5343,
   input         cfg_dout5344,
   input         cfg_dout5345,
   input         cfg_dout5346,
   input         cfg_dout5347,
   input         cfg_dout5348,
   input         cfg_dout5349,
   input         cfg_dout5350,
   input         cfg_dout5351,
   input         cfg_dout5352,
   input         cfg_dout5353,
   input         cfg_dout5354,
   input         cfg_dout5355,
   input         cfg_dout5356,
   input         cfg_dout5357,
   input         cfg_dout5358,
   input         cfg_dout5359,
   input         cfg_dout5360,
   input         cfg_dout5361,
   input         cfg_dout5362,
   input         cfg_dout5363,
   input         cfg_dout5364,
   input         cfg_dout5365,
   input         cfg_dout5366,
   input         cfg_dout5367,
   input         cfg_dout5368,
   input         cfg_dout5369,
   input         cfg_dout5370,
   input         cfg_dout5371,
   input         cfg_dout5372,
   input         cfg_dout5373,
   input         cfg_dout5374,
   input         cfg_dout5375,
   input         cfg_dout5376,
   input         cfg_dout5377,
   input         cfg_dout5378,
   input         cfg_dout5379,
   input         cfg_dout5380,
   input         cfg_dout5381,
   input         cfg_dout5382,
   input         cfg_dout5383,
   input         cfg_dout5384,
   input         cfg_dout5385,
   input         cfg_dout5386,
   input         cfg_dout5387,
   input         cfg_dout5388,
   input         cfg_dout5389,
   input         cfg_dout5390,
   input         cfg_dout5391,
   input         cfg_dout5392,
   input         cfg_dout5393,
   input         cfg_dout5394,
   input         cfg_dout5395,
   input         cfg_dout5396,
   input         cfg_dout5397,
   input         cfg_dout5398,
   input         cfg_dout5399,
   input         cfg_dout5400,
   input         cfg_dout5401,
   input         cfg_dout5402,
   input         cfg_dout5403,
   input         cfg_dout5404,
   input         cfg_dout5405,
   input         cfg_dout5406,
   input         cfg_dout5407,
   input         cfg_dout5408,
   input         cfg_dout5409,
   input         cfg_dout5410,
   input         cfg_dout5411,
   input         cfg_dout5412,
   input         cfg_dout5413,
   input         cfg_dout5414,
   input         cfg_dout5415,
   input         cfg_dout5416,
   input         cfg_dout5417,
   input         cfg_dout5418,
   input         cfg_dout5419,
   input         cfg_dout5420,
   input         cfg_dout5421,
   input         cfg_dout5422,
   input         cfg_dout5423,
   input         cfg_dout5424,
   input         cfg_dout5425,
   input         cfg_dout5426,
   input         cfg_dout5427,
   input         cfg_dout5428,
   input         cfg_dout5429,
   input         cfg_dout5430,
   input         cfg_dout5431,
   input         cfg_dout5432,
   input         cfg_dout5433,
   input         cfg_dout5434,
   input         cfg_dout5435,
   input         cfg_dout5436,
   input         cfg_dout5437,
   input         cfg_dout5438,
   input         cfg_dout5439,
   input         cfg_dout5440,
   input         cfg_dout5441,
   input         cfg_dout5442,
   input         cfg_dout5443,
   input         cfg_dout5444,
   input         cfg_dout5445,
   input         cfg_dout5446,
   input         cfg_dout5447,
   input         cfg_dout5448,
   input         cfg_dout5449,
   input         cfg_dout5450,
   input         cfg_dout5451,
   input         cfg_dout5452,
   input         cfg_dout5453,
   input         cfg_dout5454,
   input         cfg_dout5455,
   input         cfg_dout5456,
   input         cfg_dout5457,
   input         cfg_dout5458,
   input         cfg_dout5459,
   input         cfg_dout5460,
   input         cfg_dout5461,
   input         cfg_dout5462,
   input         cfg_dout5463,
   input         cfg_dout5464,
   input         cfg_dout5465,
   input         cfg_dout5466,
   input         cfg_dout5467,
   input         cfg_dout5468,
   input         cfg_dout5469,
   input         cfg_dout5470,
   input         cfg_dout5471,
   input         cfg_dout5472,
   input         cfg_dout5473,
   input         cfg_dout5474,
   input         cfg_dout5475,
   input         cfg_dout5476,
   input         cfg_dout5477,
   input         cfg_dout5478,
   input         cfg_dout5479,
   input         cfg_dout5480,
   input         cfg_dout5481,
   input         cfg_dout5482,
   input         cfg_dout5483,
   input         cfg_dout5484,
   input         cfg_dout5485,
   input         cfg_dout5486,
   input         cfg_dout5487,
   input         cfg_dout5488,
   input         cfg_dout5489,
   input         cfg_dout5490,
   input         cfg_dout5491,
   input         cfg_dout5492,
   input         cfg_dout5493,
   input         cfg_dout5494,
   input         cfg_dout5495,
   input         cfg_dout5496,
   input         cfg_dout5497,
   input         cfg_dout5498,
   input         cfg_dout5499,
   input         cfg_dout5500,
   input         cfg_dout5501,
   input         cfg_dout5502,
   input         cfg_dout5503,
   input         cfg_dout5504,
   input         cfg_dout5505,
   input         cfg_dout5506,
   input         cfg_dout5507,
   input         cfg_dout5508,
   input         cfg_dout5509,
   input         cfg_dout5510,
   input         cfg_dout5511,
   input         cfg_dout5512,
   input         cfg_dout5513,
   input         cfg_dout5514,
   input         cfg_dout5515,
   input         cfg_dout5516,
   input         cfg_dout5517,
   input         cfg_dout5518,
   input         cfg_dout5519,
   input         cfg_dout5520,
   input         cfg_dout5521,
   input         cfg_dout5522,
   input         cfg_dout5523,
   input         cfg_dout5524,
   input         cfg_dout5525,
   input         cfg_dout5526,
   input         cfg_dout5527,
   input         cfg_dout5528,
   input         cfg_dout5529,
   input         cfg_dout5530,
   input         cfg_dout5531,
   input         cfg_dout5532,
   input         cfg_dout5533,
   input         cfg_dout5534,
   input         cfg_dout5535,
   input         cfg_dout5536,
   input         cfg_dout5537,
   input         cfg_dout5538,
   input         cfg_dout5539,
   input         cfg_dout5540,
   input         cfg_dout5541,
   input         cfg_dout5542,
   input         cfg_dout5543,
   input         cfg_dout5544,
   input         cfg_dout5545,
   input         cfg_dout5546,
   input         cfg_dout5547,
   input         cfg_dout5548,
   input         cfg_dout5549,
   input         cfg_dout5550,
   input         cfg_dout5551,
   input         cfg_dout5552,
   input         cfg_dout5553,
   input         cfg_dout5554,
   input         cfg_dout5555,
   input         cfg_dout5556,
   input         cfg_dout5557,
   input         cfg_dout5558,
   input         cfg_dout5559,
   input         cfg_dout5560,
   input         cfg_dout5561,
   input         cfg_dout5562,
   input         cfg_dout5563,
   input         cfg_dout5564,
   input         cfg_dout5565,
   input         cfg_dout5566,
   input         cfg_dout5567,
   input         cfg_dout5568,
   input         cfg_dout5569,
   input         cfg_dout5570,
   input         cfg_dout5571,
   input         cfg_dout5572,
   input         cfg_dout5573,
   input         cfg_dout5574,
   input         cfg_dout5575,
   input         cfg_dout5576,
   input         cfg_dout5577,
   input         cfg_dout5578,
   input         cfg_dout5579,
   input         cfg_dout5580,
   input         cfg_dout5581,
   input         cfg_dout5582,
   input         cfg_dout5583,
   input         cfg_dout5584,
   input         cfg_dout5585,
   input         cfg_dout5586,
   input         cfg_dout5587,
   input         cfg_dout5588,
   input         cfg_dout5589,
   input         cfg_dout5590,
   input         cfg_dout5591,
   input         cfg_dout5592,
   input         cfg_dout5593,
   input         cfg_dout5594,
   input         cfg_dout5595,
   input         cfg_dout5596,
   input         cfg_dout5597,
   input         cfg_dout5598,
   input         cfg_dout5599,
   input         cfg_dout5600,
   input         cfg_dout5601,
   input         cfg_dout5602,
   input         cfg_dout5603,
   input         cfg_dout5604,
   input         cfg_dout5605,
   input         cfg_dout5606,
   input         cfg_dout5607,
   input         cfg_dout5608,
   input         cfg_dout5609,
   input         cfg_dout5610,
   input         cfg_dout5611,
   input         cfg_dout5612,
   input         cfg_dout5613,
   input         cfg_dout5614,
   input         cfg_dout5615,
   input         cfg_dout5616,
   input         cfg_dout5617,
   input         cfg_dout5618,
   input         cfg_dout5619,
   input         cfg_dout5620,
   input         cfg_dout5621,
   input         cfg_dout5622,
   input         cfg_dout5623,
   input         cfg_dout5624,
   input         cfg_dout5625,
   input         cfg_dout5626,
   input         cfg_dout5627,
   input         cfg_dout5628,
   input         cfg_dout5629,
   input         cfg_dout5630,
   input         cfg_dout5631,
   input         cfg_dout5632,
   input         cfg_dout5633,
   input         cfg_dout5634,
   input         cfg_dout5635,
   input         cfg_dout5636,
   input         cfg_dout5637,
   input         cfg_dout5638,
   input         cfg_dout5639,
   input         cfg_dout5640,
   input         cfg_dout5641,
   input         cfg_dout5642,
   input         cfg_dout5643,
   input         cfg_dout5644,
   input         cfg_dout5645,
   input         cfg_dout5646,
   input         cfg_dout5647,
   input         cfg_dout5648,
   input         cfg_dout5649,
   input         cfg_dout5650,
   input         cfg_dout5651,
   input         cfg_dout5652,
   input         cfg_dout5653,
   input         cfg_dout5654,
   input         cfg_dout5655,
   input         cfg_dout5656,
   input         cfg_dout5657,
   input         cfg_dout5658,
   input         cfg_dout5659,
   input         cfg_dout5660,
   input         cfg_dout5661,
   input         cfg_dout5662,
   input         cfg_dout5663,
   input         cfg_dout5664,
   input         cfg_dout5665,
   input         cfg_dout5666,
   input         cfg_dout5667,
   input         cfg_dout5668,
   input         cfg_dout5669,
   input         cfg_dout5670,
   input         cfg_dout5671,
   input         cfg_dout5672,
   input         cfg_dout5673,
   input         cfg_dout5674,
   input         cfg_dout5675,
   input         cfg_dout5676,
   input         cfg_dout5677,
   input         cfg_dout5678,
   input         cfg_dout5679,
   input         cfg_dout5680,
   input         cfg_dout5681,
   input         cfg_dout5682,
   input         cfg_dout5683,
   input         cfg_dout5684,
   input         cfg_dout5685,
   input         cfg_dout5686,
   input         cfg_dout5687,
   input         cfg_dout5688,
   input         cfg_dout5689,
   input         cfg_dout5690,
   input         cfg_dout5691,
   input         cfg_dout5692,
   input         cfg_dout5693,
   input         cfg_dout5694,
   input         cfg_dout5695,
   input         cfg_dout5696,
   input         cfg_dout5697,
   input         cfg_dout5698,
   input         cfg_dout5699,
   input         cfg_dout5700,
   input         cfg_dout5701,
   input         cfg_dout5702,
   input         cfg_dout5703,
   input         cfg_dout5704,
   input         cfg_dout5705,
   input         cfg_dout5706,
   input         cfg_dout5707,
   input         cfg_dout5708,
   input         cfg_dout5709,
   input         cfg_dout5710,
   input         cfg_dout5711,
   input         cfg_dout5712,
   input         cfg_dout5713,
   input         cfg_dout5714,
   input         cfg_dout5715,
   input         cfg_dout5716,
   input         cfg_dout5717,
   input         cfg_dout5718,
   input         cfg_dout5719,
   input         cfg_dout5720,
   input         cfg_dout5721,
   input         cfg_dout5722,
   input         cfg_dout5723,
   input         cfg_dout5724,
   input         cfg_dout5725,
   input         cfg_dout5726,
   input         cfg_dout5727,
   input         cfg_dout5728,
   input         cfg_dout5729,
   input         cfg_dout5730,
   input         cfg_dout5731,
   input         cfg_dout5732,
   input         cfg_dout5733,
   input         cfg_dout5734,
   input         cfg_dout5735,
   input         cfg_dout5736,
   input         cfg_dout5737,
   input         cfg_dout5738,
   input         cfg_dout5739,
   input         cfg_dout5740,
   input         cfg_dout5741,
   input         cfg_dout5742,
   input         cfg_dout5743,
   input         cfg_dout5744,
   input         cfg_dout5745,
   input         cfg_dout5746,
   input         cfg_dout5747,
   input         cfg_dout5748,
   input         cfg_dout5749,
   input         cfg_dout5750,
   input         cfg_dout5751,
   input         cfg_dout5752,
   input         cfg_dout5753,
   input         cfg_dout5754,
   input         cfg_dout5755,
   input         cfg_dout5756,
   input         cfg_dout5757,
   input         cfg_dout5758,
   input         cfg_dout5759,
   input         cfg_dout5760,
   input         cfg_dout5761,
   input         cfg_dout5762,
   input         cfg_dout5763,
   input         cfg_dout5764,
   input         cfg_dout5765,
   input         cfg_dout5766,
   input         cfg_dout5767,
   input         cfg_dout5768,
   input         cfg_dout5769,
   input         cfg_dout5770,
   input         cfg_dout5771,
   input         cfg_dout5772,
   input         cfg_dout5773,
   input         cfg_dout5774,
   input         cfg_dout5775,
   input         cfg_dout5776,
   input         cfg_dout5777,
   input         cfg_dout5778,
   input         cfg_dout5779,
   input         cfg_dout5780,
   input         cfg_dout5781,
   input         cfg_dout5782,
   input         cfg_dout5783,
   input         cfg_dout5784,
   input         cfg_dout5785,
   input         cfg_dout5786,
   input         cfg_dout5787,
   input         cfg_dout5788,
   input         cfg_dout5789,
   input         cfg_dout5790,
   input         cfg_dout5791,
   input         cfg_dout5792,
   input         cfg_dout5793,
   input         cfg_dout5794,
   input         cfg_dout5795,
   input         cfg_dout5796,
   input         cfg_dout5797,
   input         cfg_dout5798,
   input         cfg_dout5799,
   input         cfg_dout5800,
   input         cfg_dout5801,
   input         cfg_dout5802,
   input         cfg_dout5803,
   input         cfg_dout5804,
   input         cfg_dout5805,
   input         cfg_dout5806,
   input         cfg_dout5807,
   input         cfg_dout5808,
   input         cfg_dout5809,
   input         cfg_dout5810,
   input         cfg_dout5811,
   input         cfg_dout5812,
   input         cfg_dout5813,
   input         cfg_dout5814,
   input         cfg_dout5815,
   input         cfg_dout5816,
   input         cfg_dout5817,
   input         cfg_dout5818,
   input         cfg_dout5819,
   input         cfg_dout5820,
   input         cfg_dout5821,
   input         cfg_dout5822,
   input         cfg_dout5823,
   input         cfg_dout5824,
   input         cfg_dout5825,
   input         cfg_dout5826,
   input         cfg_dout5827,
   input         cfg_dout5828,
   input         cfg_dout5829,
   input         cfg_dout5830,
   input         cfg_dout5831,
   input         cfg_dout5832,
   input         cfg_dout5833,
   input         cfg_dout5834,
   input         cfg_dout5835,
   input         cfg_dout5836,
   input         cfg_dout5837,
   input         cfg_dout5838,
   input         cfg_dout5839,
   input         cfg_dout5840,
   input         cfg_dout5841,
   input         cfg_dout5842,
   input         cfg_dout5843,
   input         cfg_dout5844,
   input         cfg_dout5845,
   input         cfg_dout5846,
   input         cfg_dout5847,
   input         cfg_dout5848,
   input         cfg_dout5849,
   input         cfg_dout5850,
   input         cfg_dout5851,
   input         cfg_dout5852,
   input         cfg_dout5853,
   input         cfg_dout5854,
   input         cfg_dout5855,
   input         cfg_dout5856,
   input         cfg_dout5857,
   input         cfg_dout5858,
   input         cfg_dout5859,
   input         cfg_dout5860,
   input         cfg_dout5861,
   input         cfg_dout5862,
   input         cfg_dout5863,
   input         cfg_dout5864,
   input         cfg_dout5865,
   input         cfg_dout5866,
   input         cfg_dout5867,
   input         cfg_dout5868,
   input         cfg_dout5869,
   input         cfg_dout5870,
   input         cfg_dout5871,
   input         cfg_dout5872,
   input         cfg_dout5873,
   input         cfg_dout5874,
   input         cfg_dout5875,
   input         cfg_dout5876,
   input         cfg_dout5877,
   input         cfg_dout5878,
   input         cfg_dout5879,
   input         cfg_dout5880,
   input         cfg_dout5881,
   input         cfg_dout5882,
   input         cfg_dout5883,
   input         cfg_dout5884,
   input         cfg_dout5885,
   input         cfg_dout5886,
   input         cfg_dout5887,
   input         cfg_dout5888,
   input         cfg_dout5889,
   input         cfg_dout5890,
   input         cfg_dout5891,
   input         cfg_dout5892,
   input         cfg_dout5893,
   input         cfg_dout5894,
   input         cfg_dout5895,
   input         cfg_dout5896,
   input         cfg_dout5897,
   input         cfg_dout5898,
   input         cfg_dout5899,
   input         cfg_dout5900,
   input         cfg_dout5901,
   input         cfg_dout5902,
   input         cfg_dout5903,
   input         cfg_dout5904,
   input         cfg_dout5905,
   input         cfg_dout5906,
   input         cfg_dout5907,
   input         cfg_dout5908,
   input         cfg_dout5909,
   input         cfg_dout5910,
   input         cfg_dout5911,
   input         cfg_dout5912,
   input         cfg_dout5913,
   input         cfg_dout5914,
   input         cfg_dout5915,
   input         cfg_dout5916,
   input         cfg_dout5917,
   input         cfg_dout5918,
   input         cfg_dout5919,
   input         cfg_dout5920,
   input         cfg_dout5921,
   input         cfg_dout5922,
   input         cfg_dout5923,
   input         cfg_dout5924,
   input         cfg_dout5925,
   input         cfg_dout5926,
   input         cfg_dout5927,
   input         cfg_dout5928,
   input         cfg_dout5929,
   input         cfg_dout5930,
   input         cfg_dout5931,
   input         cfg_dout5932,
   input         cfg_dout5933,
   input         cfg_dout5934,
   input         cfg_dout5935,
   input         cfg_dout5936,
   input         cfg_dout5937,
   input         cfg_dout5938,
   input         cfg_dout5939,
   input         cfg_dout5940,
   input         cfg_dout5941,
   input         cfg_dout5942,
   input         cfg_dout5943,
   input         cfg_dout5944,
   input         cfg_dout5945,
   input         cfg_dout5946,
   input         cfg_dout5947,
   input         cfg_dout5948,
   input         cfg_dout5949,
   input         cfg_dout5950,
   input         cfg_dout5951,
   input         cfg_dout5952,
   input         cfg_dout5953,
   input         cfg_dout5954,
   input         cfg_dout5955,
   input         cfg_dout5956,
   input         cfg_dout5957,
   input         cfg_dout5958,
   input         cfg_dout5959,
   input         cfg_dout5960,
   input         cfg_dout5961,
   input         cfg_dout5962,
   input         cfg_dout5963,
   input         cfg_dout5964,
   input         cfg_dout5965,
   input         cfg_dout5966,
   input         cfg_dout5967,
   input         cfg_dout5968,
   input         cfg_dout5969,
   input         cfg_dout5970,
   input         cfg_dout5971,
   input         cfg_dout5972,
   input         cfg_dout5973,
   input         cfg_dout5974,
   input         cfg_dout5975,
   input         cfg_dout5976,
   input         cfg_dout5977,
   input         cfg_dout5978,
   input         cfg_dout5979,
   input         cfg_dout5980,
   input         cfg_dout5981,
   input         cfg_dout5982,
   input         cfg_dout5983,
   input         cfg_dout5984,
   input         cfg_dout5985,
   input         cfg_dout5986,
   input         cfg_dout5987,
   input         cfg_dout5988,
   input         cfg_dout5989,
   input         cfg_dout5990,
   input         cfg_dout5991,
   input         cfg_dout5992,
   input         cfg_dout5993,
   input         cfg_dout5994,
   input         cfg_dout5995,
   input         cfg_dout5996,
   input         cfg_dout5997,
   input         cfg_dout5998,
   input         cfg_dout5999,
   input         cfg_dout6000,
   input         cfg_dout6001,
   input         cfg_dout6002,
   input         cfg_dout6003,
   input         cfg_dout6004,
   input         cfg_dout6005,
   input         cfg_dout6006,
   input         cfg_dout6007,
   input         cfg_dout6008,
   input         cfg_dout6009,
   input         cfg_dout6010,
   input         cfg_dout6011,
   input         cfg_dout6012,
   input         cfg_dout6013,
   input         cfg_dout6014,
   input         cfg_dout6015,
   input         cfg_dout6016,
   input         cfg_dout6017,
   input         cfg_dout6018,
   input         cfg_dout6019,
   input         cfg_dout6020,
   input         cfg_dout6021,
   input         cfg_dout6022,
   input         cfg_dout6023,
   input         cfg_dout6024,
   input         cfg_dout6025,
   input         cfg_dout6026,
   input         cfg_dout6027,
   input         cfg_dout6028,
   input         cfg_dout6029,
   input         cfg_dout6030,
   input         cfg_dout6031,
   input         cfg_dout6032,
   input         cfg_dout6033,
   input         cfg_dout6034,
   input         cfg_dout6035,
   input         cfg_dout6036,
   input         cfg_dout6037,
   input         cfg_dout6038,
   input         cfg_dout6039,
   input         cfg_dout6040,
   input         cfg_dout6041,
   input         cfg_dout6042,
   input         cfg_dout6043,
   input         cfg_dout6044,
   input         cfg_dout6045,
   input         cfg_dout6046,
   input         cfg_dout6047,
   input         cfg_dout6048,
   input         cfg_dout6049,
   input         cfg_dout6050,
   input         cfg_dout6051,
   input         cfg_dout6052,
   input         cfg_dout6053,
   input         cfg_dout6054,
   input         cfg_dout6055,
   input         cfg_dout6056,
   input         cfg_dout6057,
   input         cfg_dout6058,
   input         cfg_dout6059,
   input         cfg_dout6060,
   input         cfg_dout6061,
   input         cfg_dout6062,
   input         cfg_dout6063,
   input         cfg_dout6064,
   input         cfg_dout6065,
   input         cfg_dout6066,
   input         cfg_dout6067,
   input         cfg_dout6068,
   input         cfg_dout6069,
   input         cfg_dout6070,
   input         cfg_dout6071,
   input         cfg_dout6072,
   input         cfg_dout6073,
   input         cfg_dout6074,
   input         cfg_dout6075,
   input         cfg_dout6076,
   input         cfg_dout6077,
   input         cfg_dout6078,
   input         cfg_dout6079,
   input         cfg_dout6080,
   input         cfg_dout6081,
   input         cfg_dout6082,
   input         cfg_dout6083,
   input         cfg_dout6084,
   input         cfg_dout6085,
   input         cfg_dout6086,
   input         cfg_dout6087,
   input         cfg_dout6088,
   input         cfg_dout6089,
   input         cfg_dout6090,
   input         cfg_dout6091,
   input         cfg_dout6092,
   input         cfg_dout6093,
   input         cfg_dout6094,
   input         cfg_dout6095,
   input         cfg_dout6096,
   input         cfg_dout6097,
   input         cfg_dout6098,
   input         cfg_dout6099,
   input         cfg_dout6100,
   input         cfg_dout6101,
   input         cfg_dout6102,
   input         cfg_dout6103,
   input         cfg_dout6104,
   input         cfg_dout6105,
   input         cfg_dout6106,
   input         cfg_dout6107,
   input         cfg_dout6108,
   input         cfg_dout6109,
   input         cfg_dout6110,
   input         cfg_dout6111,
   input         cfg_dout6112,
   input         cfg_dout6113,
   input         cfg_dout6114,
   input         cfg_dout6115,
   input         cfg_dout6116,
   input         cfg_dout6117,
   input         cfg_dout6118,
   input         cfg_dout6119,
   input         cfg_dout6120,
   input         cfg_dout6121,
   input         cfg_dout6122,
   input         cfg_dout6123,
   input         cfg_dout6124,
   input         cfg_dout6125,
   input         cfg_dout6126,
   input         cfg_dout6127,
   input         cfg_dout6128,
   input         cfg_dout6129,
   input         cfg_dout6130,
   input         cfg_dout6131,
   input         cfg_dout6132,
   input         cfg_dout6133,
   input         cfg_dout6134,
   input         cfg_dout6135,
   input         cfg_dout6136,
   input         cfg_dout6137,
   input         cfg_dout6138,
   input         cfg_dout6139,
   input         cfg_dout6140,
   input         cfg_dout6141,
   input         cfg_dout6142,
   input         cfg_dout6143,
   input         cfg_dout6144,
   input         cfg_dout6145,
   input         cfg_dout6146,
   input         cfg_dout6147,
   input         cfg_dout6148,
   input         cfg_dout6149,
   input         cfg_dout6150,
   input         cfg_dout6151,
   input         cfg_dout6152,
   input         cfg_dout6153,
   input         cfg_dout6154,
   input         cfg_dout6155,
   input         cfg_dout6156,
   input         cfg_dout6157,
   input         cfg_dout6158,
   input         cfg_dout6159,
   input         cfg_dout6160,
   input         cfg_dout6161,
   input         cfg_dout6162,
   input         cfg_dout6163,
   input         cfg_dout6164,
   input         cfg_dout6165,
   input         cfg_dout6166,
   input         cfg_dout6167,
   input         cfg_dout6168,
   input         cfg_dout6169,
   input         cfg_dout6170,
   input         cfg_dout6171,
   input         cfg_dout6172,
   input         cfg_dout6173,
   input         cfg_dout6174,
   input         cfg_dout6175,
   input         cfg_dout6176,
   input         cfg_dout6177,
   input         cfg_dout6178,
   input         cfg_dout6179,
   input         cfg_dout6180,
   input         cfg_dout6181,
   input         cfg_dout6182,
   input         cfg_dout6183,
   input         cfg_dout6184,
   input         cfg_dout6185,
   input         cfg_dout6186,
   input         cfg_dout6187,
   input         cfg_dout6188,
   input         cfg_dout6189,
   input         cfg_dout6190,
   input         cfg_dout6191,
   input         cfg_dout6192,
   input         cfg_dout6193,
   input         cfg_dout6194,
   input         cfg_dout6195,
   input         cfg_dout6196,
   input         cfg_dout6197,
   input         cfg_dout6198,
   input         cfg_dout6199,
   input         cfg_dout6200,
   input         cfg_dout6201,
   input         cfg_dout6202,
   input         cfg_dout6203,
   input         cfg_dout6204,
   input         cfg_dout6205,
   input         cfg_dout6206,
   input         cfg_dout6207,
   input         cfg_dout6208,
   input         cfg_dout6209,
   input         cfg_dout6210,
   input         cfg_dout6211,
   input         cfg_dout6212,
   input         cfg_dout6213,
   input         cfg_dout6214,
   input         cfg_dout6215,
   input         cfg_dout6216,
   input         cfg_dout6217,
   input         cfg_dout6218,
   input         cfg_dout6219,
   input         cfg_dout6220,
   input         cfg_dout6221,
   input         cfg_dout6222,
   input         cfg_dout6223,
   input         cfg_dout6224,
   input         cfg_dout6225,
   input         cfg_dout6226,
   input         cfg_dout6227,
   input         cfg_dout6228,
   input         cfg_dout6229,
   input         cfg_dout6230,
   input         cfg_dout6231,
   input         cfg_dout6232,
   input         cfg_dout6233,
   input         cfg_dout6234,
   input         cfg_dout6235,
   input         cfg_dout6236,
   input         cfg_dout6237,
   input         cfg_dout6238,
   input         cfg_dout6239,
   input         cfg_dout6240,
   input         cfg_dout6241,
   input         cfg_dout6242,
   input         cfg_dout6243,
   input         cfg_dout6244,
   input         cfg_dout6245,
   input         cfg_dout6246,
   input         cfg_dout6247,
   input         cfg_dout6248,
   input         cfg_dout6249,
   input         cfg_dout6250,
   input         cfg_dout6251,
   input         cfg_dout6252,
   input         cfg_dout6253,
   input         cfg_dout6254,
   input         cfg_dout6255,
   input         cfg_dout6256,
   input         cfg_dout6257,
   input         cfg_dout6258,
   input         cfg_dout6259,
   input         cfg_dout6260,
   input         cfg_dout6261,
   input         cfg_dout6262,
   input         cfg_dout6263,
   input         cfg_dout6264,
   input         cfg_dout6265,
   input         cfg_dout6266,
   input         cfg_dout6267,
   input         cfg_dout6268,
   input         cfg_dout6269,
   input         cfg_dout6270,
   input         cfg_dout6271,
   input         cfg_dout6272,
   input         cfg_dout6273,
   input         cfg_dout6274,
   input         cfg_dout6275,
   input         cfg_dout6276,
   input         cfg_dout6277,
   input         cfg_dout6278,
   input         cfg_dout6279,
   input         cfg_dout6280,
   input         cfg_dout6281,
   input         cfg_dout6282,
   input         cfg_dout6283,
   input         cfg_dout6284,
   input         cfg_dout6285,
   input         cfg_dout6286,
   input         cfg_dout6287,
   input         cfg_dout6288,
   input         cfg_dout6289,
   input         cfg_dout6290,
   input         cfg_dout6291,
   input         cfg_dout6292,
   input         cfg_dout6293,
   input         cfg_dout6294,
   input         cfg_dout6295,
   input         cfg_dout6296,
   input         cfg_dout6297,
   input         cfg_dout6298,
   input         cfg_dout6299,
   input         cfg_dout6300,
   input         cfg_dout6301,
   input         cfg_dout6302,
   input         cfg_dout6303,
   input         cfg_dout6304,
   input         cfg_dout6305,
   input         cfg_dout6306,
   input         cfg_dout6307,
   input         cfg_dout6308,
   input         cfg_dout6309,
   input         cfg_dout6310,
   input         cfg_dout6311,
   input         cfg_dout6312,
   input         cfg_dout6313,
   input         cfg_dout6314,
   input         cfg_dout6315,
   input         cfg_dout6316,
   input         cfg_dout6317,
   input         cfg_dout6318,
   input         cfg_dout6319,
   input         cfg_dout6320,
   input         cfg_dout6321,
   input         cfg_dout6322,
   input         cfg_dout6323,
   input         cfg_dout6324,
   input         cfg_dout6325,
   input         cfg_dout6326,
   input         cfg_dout6327,
   input         cfg_dout6328,
   input         cfg_dout6329,
   input         cfg_dout6330,
   input         cfg_dout6331,
   input         cfg_dout6332,
   input         cfg_dout6333,
   input         cfg_dout6334,
   input         cfg_dout6335,
   input         cfg_dout6336,
   input         cfg_dout6337,
   input         cfg_dout6338,
   input         cfg_dout6339,
   input         cfg_dout6340,
   input         cfg_dout6341,
   input         cfg_dout6342,
   input         cfg_dout6343,
   input         cfg_dout6344,
   input         cfg_dout6345,
   input         cfg_dout6346,
   input         cfg_dout6347,
   input         cfg_dout6348,
   input         cfg_dout6349,
   input         cfg_dout6350,
   input         cfg_dout6351,
   input         cfg_dout6352,
   input         cfg_dout6353,
   input         cfg_dout6354,
   input         cfg_dout6355,
   input         cfg_dout6356,
   input         cfg_dout6357,
   input         cfg_dout6358,
   input         cfg_dout6359,
   input         cfg_dout6360,
   input         cfg_dout6361,
   input         cfg_dout6362,
   input         cfg_dout6363,
   input         cfg_dout6364,
   input         cfg_dout6365,
   input         cfg_dout6366,
   input         cfg_dout6367,
   input         cfg_dout6368,
   input         cfg_dout6369,
   input         cfg_dout6370,
   input         cfg_dout6371,
   input         cfg_dout6372,
   input         cfg_dout6373,
   input         cfg_dout6374,
   input         cfg_dout6375,
   input         cfg_dout6376,
   input         cfg_dout6377,
   input         cfg_dout6378,
   input         cfg_dout6379,
   input         cfg_dout6380,
   input         cfg_dout6381,
   input         cfg_dout6382,
   input         cfg_dout6383,
   input         cfg_dout6384,
   input         cfg_dout6385,
   input         cfg_dout6386,
   input         cfg_dout6387,
   input         cfg_dout6388,
   input         cfg_dout6389,
   input         cfg_dout6390,
   input         cfg_dout6391,
   input         cfg_dout6392,
   input         cfg_dout6393,
   input         cfg_dout6394,
   input         cfg_dout6395,
   input         cfg_dout6396,
   input         cfg_dout6397,
   input         cfg_dout6398,
   input         cfg_dout6399,
   input         cfg_dout6400,
   input         cfg_dout6401,
   input         cfg_dout6402,
   input         cfg_dout6403,
   input         cfg_dout6404,
   input         cfg_dout6405,
   input         cfg_dout6406,
   input         cfg_dout6407,
   input         cfg_dout6408,
   input         cfg_dout6409,
   input         cfg_dout6410,
   input         cfg_dout6411,
   input         cfg_dout6412,
   input         cfg_dout6413,
   input         cfg_dout6414,
   input         cfg_dout6415,
   input         cfg_dout6416,
   input         cfg_dout6417,
   input         cfg_dout6418,
   input         cfg_dout6419,
   input         cfg_dout6420,
   input         cfg_dout6421,
   input         cfg_dout6422,
   input         cfg_dout6423,
   input         cfg_dout6424,
   input         cfg_dout6425,
   input         cfg_dout6426,
   input         cfg_dout6427,
   input         cfg_dout6428,
   input         cfg_dout6429,
   input         cfg_dout6430,
   input         cfg_dout6431,
   input         cfg_dout6432,
   input         cfg_dout6433,
   input         cfg_dout6434,
   input         cfg_dout6435,
   input         cfg_dout6436,
   input         cfg_dout6437,
   input         cfg_dout6438,
   input         cfg_dout6439,
   input         cfg_dout6440,
   input         cfg_dout6441,
   input         cfg_dout6442,
   input         cfg_dout6443,
   input         cfg_dout6444,
   input         cfg_dout6445,
   input         cfg_dout6446,
   input         cfg_dout6447,
   input         cfg_dout6448,
   input         cfg_dout6449,
   input         cfg_dout6450,
   input         cfg_dout6451,
   input         cfg_dout6452,
   input         cfg_dout6453,
   input         cfg_dout6454,
   input         cfg_dout6455,
   input         cfg_dout6456,
   input         cfg_dout6457,
   input         cfg_dout6458,
   input         cfg_dout6459,
   input         cfg_dout6460,
   input         cfg_dout6461,
   input         cfg_dout6462,
   input         cfg_dout6463,
   input         cfg_dout6464,
   input         cfg_dout6465,
   input         cfg_dout6466,
   input         cfg_dout6467,
   input         cfg_dout6468,
   input         cfg_dout6469,
   input         cfg_dout6470,
   input         cfg_dout6471,
   input         cfg_dout6472,
   input         cfg_dout6473,
   input         cfg_dout6474,
   input         cfg_dout6475,
   input         cfg_dout6476,
   input         cfg_dout6477,
   input         cfg_dout6478,
   input         cfg_dout6479,
   input         cfg_dout6480,
   input         cfg_dout6481,
   input         cfg_dout6482,
   input         cfg_dout6483,
   input         cfg_dout6484,
   input         cfg_dout6485,
   input         cfg_dout6486,
   input         cfg_dout6487,
   input         cfg_dout6488,
   input         cfg_dout6489,
   input         cfg_dout6490,
   input         cfg_dout6491,
   input         cfg_dout6492,
   input         cfg_dout6493,
   input         cfg_dout6494,
   input         cfg_dout6495,
   input         cfg_dout6496,
   input         cfg_dout6497,
   input         cfg_dout6498,
   input         cfg_dout6499,
   input         cfg_dout6500,
   input         cfg_dout6501,
   input         cfg_dout6502,
   input         cfg_dout6503,
   input         cfg_dout6504,
   input         cfg_dout6505,
   input         cfg_dout6506,
   input         cfg_dout6507,
   input         cfg_dout6508,
   input         cfg_dout6509,
   input         cfg_dout6510,
   input         cfg_dout6511,
   input         cfg_dout6512,
   input         cfg_dout6513,
   input         cfg_dout6514,
   input         cfg_dout6515,
   input         cfg_dout6516,
   input         cfg_dout6517,
   input         cfg_dout6518,
   input         cfg_dout6519,
   input         cfg_dout6520,
   input         cfg_dout6521,
   input         cfg_dout6522,
   input         cfg_dout6523,
   input         cfg_dout6524,
   input         cfg_dout6525,
   input         cfg_dout6526,
   input         cfg_dout6527,
   input         cfg_dout6528,
   input         cfg_dout6529,
   input         cfg_dout6530,
   input         cfg_dout6531,
   input         cfg_dout6532,
   input         cfg_dout6533,
   input         cfg_dout6534,
   input         cfg_dout6535,
   input         cfg_dout6536,
   input         cfg_dout6537,
   input         cfg_dout6538,
   input         cfg_dout6539,
   input         cfg_dout6540,
   input         cfg_dout6541,
   input         cfg_dout6542,
   input         cfg_dout6543,
   input         cfg_dout6544,
   input         cfg_dout6545,
   input         cfg_dout6546,
   input         cfg_dout6547,
   input         cfg_dout6548,
   input         cfg_dout6549,
   input         cfg_dout6550,
   input         cfg_dout6551,
   input         cfg_dout6552,
   input         cfg_dout6553,
   input         cfg_dout6554,
   input         cfg_dout6555,
   input         cfg_dout6556,
   input         cfg_dout6557,
   input         cfg_dout6558,
   input         cfg_dout6559,
   input         cfg_dout6560,
   input         cfg_dout6561,
   input         cfg_dout6562,
   input         cfg_dout6563,
   input         cfg_dout6564,
   input         cfg_dout6565,
   input         cfg_dout6566,
   input         cfg_dout6567,
   input         cfg_dout6568,
   input         cfg_dout6569,
   input         cfg_dout6570,
   input         cfg_dout6571,
   input         cfg_dout6572,
   input         cfg_dout6573,
   input         cfg_dout6574,
   input         cfg_dout6575,
   input         cfg_dout6576,
   input         cfg_dout6577,
   input         cfg_dout6578,
   input         cfg_dout6579,
   input         cfg_dout6580,
   input         cfg_dout6581,
   input         cfg_dout6582,
   input         cfg_dout6583,
   input         cfg_dout6584,
   input         cfg_dout6585,
   input         cfg_dout6586,
   input         cfg_dout6587,
   input         cfg_dout6588,
   input         cfg_dout6589,
   input         cfg_dout6590,
   input         cfg_dout6591,
   input         cfg_dout6592,
   input         cfg_dout6593,
   input         cfg_dout6594,
   input         cfg_dout6595,
   input         cfg_dout6596,
   input         cfg_dout6597,
   input         cfg_dout6598,
   input         cfg_dout6599,
   input         cfg_dout6600,
   input         cfg_dout6601,
   input         cfg_dout6602,
   input         cfg_dout6603,
   input         cfg_dout6604,
   input         cfg_dout6605,
   input         cfg_dout6606,
   input         cfg_dout6607,
   input         cfg_dout6608,
   input         cfg_dout6609,
   input         cfg_dout6610,
   input         cfg_dout6611,
   input         cfg_dout6612,
   input         cfg_dout6613,
   input         cfg_dout6614,
   input         cfg_dout6615,
   input         cfg_dout6616,
   input         cfg_dout6617,
   input         cfg_dout6618,
   input         cfg_dout6619,
   input         cfg_dout6620,
   input         cfg_dout6621,
   input         cfg_dout6622,
   input         cfg_dout6623,
   input         cfg_dout6624,
   input         cfg_dout6625,
   input         cfg_dout6626,
   input         cfg_dout6627,
   input         cfg_dout6628,
   input         cfg_dout6629,
   input         cfg_dout6630,
   input         cfg_dout6631,
   input         cfg_dout6632,
   input         cfg_dout6633,
   input         cfg_dout6634,
   input         cfg_dout6635,
   input         cfg_dout6636,
   input         cfg_dout6637,
   input         cfg_dout6638,
   input         cfg_dout6639,
   input         cfg_dout6640,
   input         cfg_dout6641,
   input         cfg_dout6642,
   input         cfg_dout6643,
   input         cfg_dout6644,
   input         cfg_dout6645,
   input         cfg_dout6646,
   input         cfg_dout6647,
   input         cfg_dout6648,
   input         cfg_dout6649,
   input         cfg_dout6650,
   input         cfg_dout6651,
   input         cfg_dout6652,
   input         cfg_dout6653,
   input         cfg_dout6654,
   input         cfg_dout6655,
   input         cfg_dout6656,
   input         cfg_dout6657,
   input         cfg_dout6658,
   input         cfg_dout6659,
   input         cfg_dout6660,
   input         cfg_dout6661,
   input         cfg_dout6662,
   input         cfg_dout6663,
   input         cfg_dout6664,
   input         cfg_dout6665,
   input         cfg_dout6666,
   input         cfg_dout6667,
   input         cfg_dout6668,
   input         cfg_dout6669,
   input         cfg_dout6670,
   input         cfg_dout6671,
   input         cfg_dout6672,
   input         cfg_dout6673,
   input         cfg_dout6674,
   input         cfg_dout6675,
   input         cfg_dout6676,
   input         cfg_dout6677,
   input         cfg_dout6678,
   input         cfg_dout6679,
   input         cfg_dout6680,
   input         cfg_dout6681,
   input         cfg_dout6682,
   input         cfg_dout6683,
   input         cfg_dout6684,
   input         cfg_dout6685,
   input         cfg_dout6686,
   input         cfg_dout6687,
   input         cfg_dout6688,
   input         cfg_dout6689,
   input         cfg_dout6690,
   input         cfg_dout6691,
   input         cfg_dout6692,
   input         cfg_dout6693,
   input         cfg_dout6694,
   input         cfg_dout6695,
   input         cfg_dout6696,
   input         cfg_dout6697,
   input         cfg_dout6698,
   input         cfg_dout6699,
   input         cfg_dout6700,
   input         cfg_dout6701,
   input         cfg_dout6702,
   input         cfg_dout6703,
   input         cfg_dout6704,
   input         cfg_dout6705,
   input         cfg_dout6706,
   input         cfg_dout6707,
   input         cfg_dout6708,
   input         cfg_dout6709,
   input         cfg_dout6710,
   input         cfg_dout6711,
   input         cfg_dout6712,
   input         cfg_dout6713,
   input         cfg_dout6714,
   input         cfg_dout6715,
   input         cfg_dout6716,
   input         cfg_dout6717,
   input         cfg_dout6718,
   input         cfg_dout6719,
   input         cfg_dout6720,
   input         cfg_dout6721,
   input         cfg_dout6722,
   input         cfg_dout6723,
   input         cfg_dout6724,
   input         cfg_dout6725,
   input         cfg_dout6726,
   input         cfg_dout6727,
   input         cfg_dout6728,
   input         cfg_dout6729,
   input         cfg_dout6730,
   input         cfg_dout6731,
   input         cfg_dout6732,
   input         cfg_dout6733,
   input         cfg_dout6734,
   input         cfg_dout6735,
   input         cfg_dout6736,
   input         cfg_dout6737,
   input         cfg_dout6738,
   input         cfg_dout6739,
   input         cfg_dout6740,
   input         cfg_dout6741,
   input         cfg_dout6742,
   input         cfg_dout6743,
   input         cfg_dout6744,
   input         cfg_dout6745,
   input         cfg_dout6746,
   input         cfg_dout6747,
   input         cfg_dout6748,
   input         cfg_dout6749,
   input         cfg_dout6750,
   input         cfg_dout6751,
   input         cfg_dout6752,
   input         cfg_dout6753,
   input         cfg_dout6754,
   input         cfg_dout6755,
   input         cfg_dout6756,
   input         cfg_dout6757,
   input         cfg_dout6758,
   input         cfg_dout6759,
   input         cfg_dout6760,
   input         cfg_dout6761,
   input         cfg_dout6762,
   input         cfg_dout6763,
   input         cfg_dout6764,
   input         cfg_dout6765,
   input         cfg_dout6766,
   input         cfg_dout6767,
   input         cfg_dout6768,
   input         cfg_dout6769,
   input         cfg_dout6770,
   input         cfg_dout6771,
   input         cfg_dout6772,
   input         cfg_dout6773,
   input         cfg_dout6774,
   input         cfg_dout6775,
   input         cfg_dout6776,
   input         cfg_dout6777,
   input         cfg_dout6778,
   input         cfg_dout6779,
   input         cfg_dout6780,
   input         cfg_dout6781,
   input         cfg_dout6782,
   input         cfg_dout6783,
   input         cfg_dout6784,
   input         cfg_dout6785,
   input         cfg_dout6786,
   input         cfg_dout6787,
   input         cfg_dout6788,
   input         cfg_dout6789,
   input         cfg_dout6790,
   input         cfg_dout6791,
   input         cfg_dout6792,
   input         cfg_dout6793,
   input         cfg_dout6794,
   input         cfg_dout6795,
   input         cfg_dout6796,
   input         cfg_dout6797,
   input         cfg_dout6798,
   input         cfg_dout6799,
   input         cfg_dout6800,
   input         cfg_dout6801,
   input         cfg_dout6802,
   input         cfg_dout6803,
   input         cfg_dout6804,
   input         cfg_dout6805,
   input         cfg_dout6806,
   input         cfg_dout6807,
   input         cfg_dout6808,
   input         cfg_dout6809,
   input         cfg_dout6810,
   input         cfg_dout6811,
   input         cfg_dout6812,
   input         cfg_dout6813,
   input         cfg_dout6814,
   input         cfg_dout6815,
   input         cfg_dout6816,
   input         cfg_dout6817,
   input         cfg_dout6818,
   input         cfg_dout6819,
   input         cfg_dout6820,
   input         cfg_dout6821,
   input         cfg_dout6822,
   input         cfg_dout6823,
   input         cfg_dout6824,
   input         cfg_dout6825,
   input         cfg_dout6826,
   input         cfg_dout6827,
   input         cfg_dout6828,
   input         cfg_dout6829,
   input         cfg_dout6830,
   input         cfg_dout6831,
   input         cfg_dout6832,
   input         cfg_dout6833,
   input         cfg_dout6834,
   input         cfg_dout6835,
   input         cfg_dout6836,
   input         cfg_dout6837,
   input         cfg_dout6838,
   input         cfg_dout6839,
   input         cfg_dout6840,
   input         cfg_dout6841,
   input         cfg_dout6842,
   input         cfg_dout6843,
   input         cfg_dout6844,
   input         cfg_dout6845,
   input         cfg_dout6846,
   input         cfg_dout6847,
   input         cfg_dout6848,
   input         cfg_dout6849,
   input         cfg_dout6850,
   input         cfg_dout6851,
   input         cfg_dout6852,
   input         cfg_dout6853,
   input         cfg_dout6854,
   input         cfg_dout6855,
   input         cfg_dout6856,
   input         cfg_dout6857,
   input         cfg_dout6858,
   input         cfg_dout6859,
   input         cfg_dout6860,
   input         cfg_dout6861,
   input         cfg_dout6862,
   input         cfg_dout6863,
   input         cfg_dout6864,
   input         cfg_dout6865,
   input         cfg_dout6866,
   input         cfg_dout6867,
   input         cfg_dout6868,
   input         cfg_dout6869,
   input         cfg_dout6870,
   input         cfg_dout6871,
   input         cfg_dout6872,
   input         cfg_dout6873,
   input         cfg_dout6874,
   input         cfg_dout6875,
   input         cfg_dout6876,
   input         cfg_dout6877,
   input         cfg_dout6878,
   input         cfg_dout6879,
   input         cfg_dout6880,
   input         cfg_dout6881,
   input         cfg_dout6882,
   input         cfg_dout6883,
   input         cfg_dout6884,
   input         cfg_dout6885,
   input         cfg_dout6886,
   input         cfg_dout6887,
   input         cfg_dout6888,
   input         cfg_dout6889,
   input         cfg_dout6890,
   input         cfg_dout6891,
   input         cfg_dout6892,
   input         cfg_dout6893,
   input         cfg_dout6894,
   input         cfg_dout6895,
   input         cfg_dout6896,
   input         cfg_dout6897,
   input         cfg_dout6898,
   input         cfg_dout6899,
   input         cfg_dout6900,
   input         cfg_dout6901,
   input         cfg_dout6902,
   input         cfg_dout6903,
   input         cfg_dout6904,
   input         cfg_dout6905,
   input         cfg_dout6906,
   input         cfg_dout6907,
   input         cfg_dout6908,
   input         cfg_dout6909,
   input         cfg_dout6910,
   input         cfg_dout6911,
   input         cfg_dout6912,
   input         cfg_dout6913,
   input         cfg_dout6914,
   input         cfg_dout6915,
   input         cfg_dout6916,
   input         cfg_dout6917,
   input         cfg_dout6918,
   input         cfg_dout6919,
   input         cfg_dout6920,
   input         cfg_dout6921,
   input         cfg_dout6922,
   input         cfg_dout6923,
   input         cfg_dout6924,
   input         cfg_dout6925,
   input         cfg_dout6926,
   input         cfg_dout6927,
   input         cfg_dout6928,
   input         cfg_dout6929,
   input         cfg_dout6930,
   input         cfg_dout6931,
   input         cfg_dout6932,
   input         cfg_dout6933,
   input         cfg_dout6934,
   input         cfg_dout6935,
   input         cfg_dout6936,
   input         cfg_dout6937,
   input         cfg_dout6938,
   input         cfg_dout6939,
   input         cfg_dout6940,
   input         cfg_dout6941,
   input         cfg_dout6942,
   input         cfg_dout6943,
   input         cfg_dout6944,
   input         cfg_dout6945,
   input         cfg_dout6946,
   input         cfg_dout6947,
   input         cfg_dout6948,
   input         cfg_dout6949,
   input         cfg_dout6950,
   input         cfg_dout6951,
   input         cfg_dout6952,
   input         cfg_dout6953,
   input         cfg_dout6954,
   input         cfg_dout6955,
   input         cfg_dout6956,
   input         cfg_dout6957,
   input         cfg_dout6958,
   input         cfg_dout6959,
   input         cfg_dout6960,
   input         cfg_dout6961,
   input         cfg_dout6962,
   input         cfg_dout6963,
   input         cfg_dout6964,
   input         cfg_dout6965,
   input         cfg_dout6966,
   input         cfg_dout6967,
   input         cfg_dout6968,
   input         cfg_dout6969,
   input         cfg_dout6970,
   input         cfg_dout6971,
   input         cfg_dout6972,
   input         cfg_dout6973,
   input         cfg_dout6974,
   input         cfg_dout6975,
   input         cfg_dout6976,
   input         cfg_dout6977,
   input         cfg_dout6978,
   input         cfg_dout6979,
   input         cfg_dout6980,
   input         cfg_dout6981,
   input         cfg_dout6982,
   input         cfg_dout6983,
   input         cfg_dout6984,
   input         cfg_dout6985,
   input         cfg_dout6986,
   input         cfg_dout6987,
   input         cfg_dout6988,
   input         cfg_dout6989,
   input         cfg_dout6990,
   input         cfg_dout6991,
   input         cfg_dout6992,
   input         cfg_dout6993,
   input         cfg_dout6994,
   input         cfg_dout6995,
   input         cfg_dout6996,
   input         cfg_dout6997,
   input         cfg_dout6998,
   input         cfg_dout6999,
   input         cfg_dout7000,
   input         cfg_dout7001,
   input         cfg_dout7002,
   input         cfg_dout7003,
   input         cfg_dout7004,
   input         cfg_dout7005,
   input         cfg_dout7006,
   input         cfg_dout7007,
   input         cfg_dout7008,
   input         cfg_dout7009,
   input         cfg_dout7010,
   input         cfg_dout7011,
   input         cfg_dout7012,
   input         cfg_dout7013,
   input         cfg_dout7014,
   input         cfg_dout7015,
   input         cfg_dout7016,
   input         cfg_dout7017,
   input         cfg_dout7018,
   input         cfg_dout7019,
   input         cfg_dout7020,
   input         cfg_dout7021,
   input         cfg_dout7022,
   input         cfg_dout7023,
   input         cfg_dout7024,
   input         cfg_dout7025,
   input         cfg_dout7026,
   input         cfg_dout7027,
   input         cfg_dout7028,
   input         cfg_dout7029,
   input         cfg_dout7030,
   input         cfg_dout7031,
   input         cfg_dout7032,
   input         cfg_dout7033,
   input         cfg_dout7034,
   input         cfg_dout7035,
   input         cfg_dout7036,
   input         cfg_dout7037,
   input         cfg_dout7038,
   input         cfg_dout7039,
   input         cfg_dout7040,
   input         cfg_dout7041,
   input         cfg_dout7042,
   input         cfg_dout7043,
   input         cfg_dout7044,
   input         cfg_dout7045,
   input         cfg_dout7046,
   input         cfg_dout7047,
   input         cfg_dout7048,
   input         cfg_dout7049,
   input         cfg_dout7050,
   input         cfg_dout7051,
   input         cfg_dout7052,
   input         cfg_dout7053,
   input         cfg_dout7054,
   input         cfg_dout7055,
   input         cfg_dout7056,
   input         cfg_dout7057,
   input         cfg_dout7058,
   input         cfg_dout7059,
   input         cfg_dout7060,
   input         cfg_dout7061,
   input         cfg_dout7062,
   input         cfg_dout7063,
   input         cfg_dout7064,
   input         cfg_dout7065,
   input         cfg_dout7066,
   input         cfg_dout7067,
   input         cfg_dout7068,
   input         cfg_dout7069,
   input         cfg_dout7070,
   input         cfg_dout7071,
   input         cfg_dout7072,
   input         cfg_dout7073,
   input         cfg_dout7074,
   input         cfg_dout7075,
   input         cfg_dout7076,
   input         cfg_dout7077,
   input         cfg_dout7078,
   input         cfg_dout7079,
   input         cfg_dout7080,
   input         cfg_dout7081,
   input         cfg_dout7082,
   input         cfg_dout7083,
   input         cfg_dout7084,
   input         cfg_dout7085,
   input         cfg_dout7086,
   input         cfg_dout7087,
   input         cfg_dout7088,
   input         cfg_dout7089,
   input         cfg_dout7090,
   input         cfg_dout7091,
   input         cfg_dout7092,
   input         cfg_dout7093,
   input         cfg_dout7094,
   input         cfg_dout7095,
   input         cfg_dout7096,
   input         cfg_dout7097,
   input         cfg_dout7098,
   input         cfg_dout7099,
   input         cfg_dout7100,
   input         cfg_dout7101,
   input         cfg_dout7102,
   input         cfg_dout7103,
   input         cfg_dout7104,
   input         cfg_dout7105,
   input         cfg_dout7106,
   input         cfg_dout7107,
   input         cfg_dout7108,
   input         cfg_dout7109,
   input         cfg_dout7110,
   input         cfg_dout7111,
   input         cfg_dout7112,
   input         cfg_dout7113,
   input         cfg_dout7114,
   input         cfg_dout7115,
   input         cfg_dout7116,
   input         cfg_dout7117,
   input         cfg_dout7118,
   input         cfg_dout7119,
   input         cfg_dout7120,
   input         cfg_dout7121,
   input         cfg_dout7122,
   input         cfg_dout7123,
   input         cfg_dout7124,
   input         cfg_dout7125,
   input         cfg_dout7126,
   input         cfg_dout7127,
   input         cfg_dout7128,
   input         cfg_dout7129,
   input         cfg_dout7130,
   input         cfg_dout7131,
   input         cfg_dout7132,
   input         cfg_dout7133,
   input         cfg_dout7134,
   input         cfg_dout7135,
   input         cfg_dout7136,
   input         cfg_dout7137,
   input         cfg_dout7138,
   input         cfg_dout7139,
   input         cfg_dout7140,
   input         cfg_dout7141,
   input         cfg_dout7142,
   input         cfg_dout7143,
   input         cfg_dout7144,
   input         cfg_dout7145,
   input         cfg_dout7146,
   input         cfg_dout7147,
   input         cfg_dout7148,
   input         cfg_dout7149,
   input         cfg_dout7150,
   input         cfg_dout7151,
   input         cfg_dout7152,
   input         cfg_dout7153,
   input         cfg_dout7154,
   input         cfg_dout7155,
   input         cfg_dout7156,
   input         cfg_dout7157,
   input         cfg_dout7158,
   input         cfg_dout7159,
   input         cfg_dout7160,
   input         cfg_dout7161,
   input         cfg_dout7162,
   input         cfg_dout7163,
   input         cfg_dout7164,
   input         cfg_dout7165,
   input         cfg_dout7166,
   input         cfg_dout7167,
   input         cfg_dout7168,
   input         cfg_dout7169,
   input         cfg_dout7170,
   input         cfg_dout7171,
   input         cfg_dout7172,
   input         cfg_dout7173,
   input         cfg_dout7174,
   input         cfg_dout7175,
   input         cfg_dout7176,
   input         cfg_dout7177,
   input         cfg_dout7178,
   input         cfg_dout7179,
   input         cfg_dout7180,
   input         cfg_dout7181,
   input         cfg_dout7182,
   input         cfg_dout7183,
   input         cfg_dout7184,
   input         cfg_dout7185,
   input         cfg_dout7186,
   input         cfg_dout7187,
   input         cfg_dout7188,
   input         cfg_dout7189,
   input         cfg_dout7190,
   input         cfg_dout7191,
   input         cfg_dout7192,
   input         cfg_dout7193,
   input         cfg_dout7194,
   input         cfg_dout7195,
   input         cfg_dout7196,
   input         cfg_dout7197,
   input         cfg_dout7198,
   input         cfg_dout7199,
   input         cfg_dout7200,
   input         cfg_dout7201,
   input         cfg_dout7202,
   input         cfg_dout7203,
   input         cfg_dout7204,
   input         cfg_dout7205,
   input         cfg_dout7206,
   input         cfg_dout7207,
   input         cfg_dout7208,
   input         cfg_dout7209,
   input         cfg_dout7210,
   input         cfg_dout7211,
   input         cfg_dout7212,
   input         cfg_dout7213,
   input         cfg_dout7214,
   input         cfg_dout7215,
   input         cfg_dout7216,
   input         cfg_dout7217,
   input         cfg_dout7218,
   input         cfg_dout7219,
   input         cfg_dout7220,
   input         cfg_dout7221,
   input         cfg_dout7222,
   input         cfg_dout7223,
   input         cfg_dout7224,
   input         cfg_dout7225,
   input         cfg_dout7226,
   input         cfg_dout7227,
   input         cfg_dout7228,
   input         cfg_dout7229,
   input         cfg_dout7230,
   input         cfg_dout7231,
   input         cfg_dout7232,
   input         cfg_dout7233,
   input         cfg_dout7234,
   input         cfg_dout7235,
   input         cfg_dout7236,
   input         cfg_dout7237,
   input         cfg_dout7238,
   input         cfg_dout7239,
   input         cfg_dout7240,
   input         cfg_dout7241,
   input         cfg_dout7242,
   input         cfg_dout7243,
   input         cfg_dout7244,
   input         cfg_dout7245,
   input         cfg_dout7246,
   input         cfg_dout7247,
   input         cfg_dout7248,
   input         cfg_dout7249,
   input         cfg_dout7250,
   input         cfg_dout7251,
   input         cfg_dout7252,
   input         cfg_dout7253,
   input         cfg_dout7254,
   input         cfg_dout7255,
   input         cfg_dout7256,
   input         cfg_dout7257,
   input         cfg_dout7258,
   input         cfg_dout7259,
   input         cfg_dout7260,
   input         cfg_dout7261,
   input         cfg_dout7262,
   input         cfg_dout7263,
   input         cfg_dout7264,
   input         cfg_dout7265,
   input         cfg_dout7266,
   input         cfg_dout7267,
   input         cfg_dout7268,
   input         cfg_dout7269,
   input         cfg_dout7270,
   input         cfg_dout7271,
   input         cfg_dout7272,
   input         cfg_dout7273,
   input         cfg_dout7274,
   input         cfg_dout7275,
   input         cfg_dout7276,
   input         cfg_dout7277,
   input         cfg_dout7278,
   input         cfg_dout7279,
   input         cfg_dout7280,
   input         cfg_dout7281,
   input         cfg_dout7282,
   input         cfg_dout7283,
   input         cfg_dout7284,
   input         cfg_dout7285,
   input         cfg_dout7286,
   input         cfg_dout7287,
   input         cfg_dout7288,
   input         cfg_dout7289,
   input         cfg_dout7290,
   input         cfg_dout7291,
   input         cfg_dout7292,
   input         cfg_dout7293,
   input         cfg_dout7294,
   input         cfg_dout7295,
   input         cfg_dout7296,
   input         cfg_dout7297,
   input         cfg_dout7298,
   input         cfg_dout7299,
   input         cfg_dout7300,
   input         cfg_dout7301,
   input         cfg_dout7302,
   input         cfg_dout7303,
   input         cfg_dout7304,
   input         cfg_dout7305,
   input         cfg_dout7306,
   input         cfg_dout7307,
   input         cfg_dout7308,
   input         cfg_dout7309,
   input         cfg_dout7310,
   input         cfg_dout7311,
   input         cfg_dout7312,
   input         cfg_dout7313,
   input         cfg_dout7314,
   input         cfg_dout7315,
   input         cfg_dout7316,
   input         cfg_dout7317,
   input         cfg_dout7318,
   input         cfg_dout7319,
   input         cfg_dout7320,
   input         cfg_dout7321,
   input         cfg_dout7322,
   input         cfg_dout7323,
   input         cfg_dout7324,
   input         cfg_dout7325,
   input         cfg_dout7326,
   input         cfg_dout7327,
   input         cfg_dout7328,
   input         cfg_dout7329,
   input         cfg_dout7330,
   input         cfg_dout7331,
   input         cfg_dout7332,
   input         cfg_dout7333,
   input         cfg_dout7334,
   input         cfg_dout7335,
   input         cfg_dout7336,
   input         cfg_dout7337,
   input         cfg_dout7338,
   input         cfg_dout7339,
   input         cfg_dout7340,
   input         cfg_dout7341,
   input         cfg_dout7342,
   input         cfg_dout7343,
   input         cfg_dout7344,
   input         cfg_dout7345,
   input         cfg_dout7346,
   input         cfg_dout7347,
   input         cfg_dout7348,
   input         cfg_dout7349,
   input         cfg_dout7350,
   input         cfg_dout7351,
   input         cfg_dout7352,
   input         cfg_dout7353,
   input         cfg_dout7354,
   input         cfg_dout7355,
   input         cfg_dout7356,
   input         cfg_dout7357,
   input         cfg_dout7358,
   input         cfg_dout7359,
   input         cfg_dout7360,
   input         cfg_dout7361,
   input         cfg_dout7362,
   input         cfg_dout7363,
   input         cfg_dout7364,
   input         cfg_dout7365,
   input         cfg_dout7366,
   input         cfg_dout7367,
   input         cfg_dout7368,
   input         cfg_dout7369,
   input         cfg_dout7370,
   input         cfg_dout7371,
   input         cfg_dout7372,
   input         cfg_dout7373,
   input         cfg_dout7374,
   input         cfg_dout7375,
   input         cfg_dout7376,
   input         cfg_dout7377,
   input         cfg_dout7378,
   input         cfg_dout7379,
   input         cfg_dout7380,
   input         cfg_dout7381,
   input         cfg_dout7382,
   input         cfg_dout7383,
   input         cfg_dout7384,
   input         cfg_dout7385,
   input         cfg_dout7386,
   input         cfg_dout7387,
   input         cfg_dout7388,
   input         cfg_dout7389,
   input         cfg_dout7390,
   input         cfg_dout7391,
   input         cfg_dout7392,
   input         cfg_dout7393,
   input         cfg_dout7394,
   input         cfg_dout7395,
   input         cfg_dout7396,
   input         cfg_dout7397,
   input         cfg_dout7398,
   input         cfg_dout7399,
   input         cfg_dout7400,
   input         cfg_dout7401,
   input         cfg_dout7402,
   input         cfg_dout7403,
   input         cfg_dout7404,
   input         cfg_dout7405,
   input         cfg_dout7406,
   input         cfg_dout7407,
   input         cfg_dout7408,
   input         cfg_dout7409,
   input         cfg_dout7410,
   input         cfg_dout7411,
   input         cfg_dout7412,
   input         cfg_dout7413,
   input         cfg_dout7414,
   input         cfg_dout7415,
   input         cfg_dout7416,
   input         cfg_dout7417,
   input         cfg_dout7418,
   input         cfg_dout7419,
   input         cfg_dout7420,
   input         cfg_dout7421,
   input         cfg_dout7422,
   input         cfg_dout7423,
   input         cfg_dout7424,
   input         cfg_dout7425,
   input         cfg_dout7426,
   input         cfg_dout7427,
   input         cfg_dout7428,
   input         cfg_dout7429,
   input         cfg_dout7430,
   input         cfg_dout7431,
   input         cfg_dout7432,
   input         cfg_dout7433,
   input         cfg_dout7434,
   input         cfg_dout7435,
   input         cfg_dout7436,
   input         cfg_dout7437,
   input         cfg_dout7438,
   input         cfg_dout7439,
   input         cfg_dout7440,
   input         cfg_dout7441,
   input         cfg_dout7442,
   input         cfg_dout7443,
   input         cfg_dout7444,
   input         cfg_dout7445,
   input         cfg_dout7446,
   input         cfg_dout7447,
   input         cfg_dout7448,
   input         cfg_dout7449,
   input         cfg_dout7450,
   input         cfg_dout7451,
   input         cfg_dout7452,
   input         cfg_dout7453,
   input         cfg_dout7454,
   input         cfg_dout7455,
   input         cfg_dout7456,
   input         cfg_dout7457,
   input         cfg_dout7458,
   input         cfg_dout7459,
   input         cfg_dout7460,
   input         cfg_dout7461,
   input         cfg_dout7462,
   input         cfg_dout7463,
   input         cfg_dout7464,
   input         cfg_dout7465,
   input         cfg_dout7466,
   input         cfg_dout7467,
   input         cfg_dout7468,
   input         cfg_dout7469,
   input         cfg_dout7470,
   input         cfg_dout7471,
   input         cfg_dout7472,
   input         cfg_dout7473,
   input         cfg_dout7474,
   input         cfg_dout7475,
   input         cfg_dout7476,
   input         cfg_dout7477,
   input         cfg_dout7478,
   input         cfg_dout7479,
   input         cfg_dout7480,
   input         cfg_dout7481,
   input         cfg_dout7482,
   input         cfg_dout7483,
   input         cfg_dout7484,
   input         cfg_dout7485,
   input         cfg_dout7486,
   input         cfg_dout7487,
   input         cfg_dout7488,
   input         cfg_dout7489,
   input         cfg_dout7490,
   input         cfg_dout7491,
   input         cfg_dout7492,
   input         cfg_dout7493,
   input         cfg_dout7494,
   input         cfg_dout7495,
   input         cfg_dout7496,
   input         cfg_dout7497,
   input         cfg_dout7498,
   input         cfg_dout7499,
   input         cfg_dout7500,
   input         cfg_dout7501,
   input         cfg_dout7502,
   input         cfg_dout7503,
   input         cfg_dout7504,
   input         cfg_dout7505,
   input         cfg_dout7506,
   input         cfg_dout7507,
   input         cfg_dout7508,
   input         cfg_dout7509,
   input         cfg_dout7510,
   input         cfg_dout7511,
   input         cfg_dout7512,
   input         cfg_dout7513,
   input         cfg_dout7514,
   input         cfg_dout7515,
   input         cfg_dout7516,
   input         cfg_dout7517,
   input         cfg_dout7518,
   input         cfg_dout7519,
   input         cfg_dout7520,
   input         cfg_dout7521,
   input         cfg_dout7522,
   input         cfg_dout7523,
   input         cfg_dout7524,
   input         cfg_dout7525,
   input         cfg_dout7526,
   input         cfg_dout7527,
   input         cfg_dout7528,
   input         cfg_dout7529,
   input         cfg_dout7530,
   input         cfg_dout7531,
   input         cfg_dout7532,
   input         cfg_dout7533,
   input         cfg_dout7534,
   input         cfg_dout7535,
   input         cfg_dout7536,
   input         cfg_dout7537,
   input         cfg_dout7538,
   input         cfg_dout7539,
   input         cfg_dout7540,
   input         cfg_dout7541,
   input         cfg_dout7542,
   input         cfg_dout7543,
   input         cfg_dout7544,
   input         cfg_dout7545,
   input         cfg_dout7546,
   input         cfg_dout7547,
   input         cfg_dout7548,
   input         cfg_dout7549,
   input         cfg_dout7550,
   input         cfg_dout7551,
   input         cfg_dout7552,
   input         cfg_dout7553,
   input         cfg_dout7554,
   input         cfg_dout7555,
   input         cfg_dout7556,
   input         cfg_dout7557,
   input         cfg_dout7558,
   input         cfg_dout7559,
   input         cfg_dout7560,
   input         cfg_dout7561,
   input         cfg_dout7562,
   input         cfg_dout7563,
   input         cfg_dout7564,
   input         cfg_dout7565,
   input         cfg_dout7566,
   input         cfg_dout7567,
   input         cfg_dout7568,
   input         cfg_dout7569,
   input         cfg_dout7570,
   input         cfg_dout7571,
   input         cfg_dout7572,
   input         cfg_dout7573,
   input         cfg_dout7574,
   input         cfg_dout7575,
   input         cfg_dout7576,
   input         cfg_dout7577,
   input         cfg_dout7578,
   input         cfg_dout7579,
   input         cfg_dout7580,
   input         cfg_dout7581,
   input         cfg_dout7582,
   input         cfg_dout7583,
   input         cfg_dout7584,
   input         cfg_dout7585,
   input         cfg_dout7586,
   input         cfg_dout7587,
   input         cfg_dout7588,
   input         cfg_dout7589,
   input         cfg_dout7590,
   input         cfg_dout7591,
   input         cfg_dout7592,
   input         cfg_dout7593,
   input         cfg_dout7594,
   input         cfg_dout7595,
   input         cfg_dout7596,
   input         cfg_dout7597,
   input         cfg_dout7598,
   input         cfg_dout7599,
   input         cfg_dout7600,
   input         cfg_dout7601,
   input         cfg_dout7602,
   input         cfg_dout7603,
   input         cfg_dout7604,
   input         cfg_dout7605,
   input         cfg_dout7606,
   input         cfg_dout7607,
   input         cfg_dout7608,
   input         cfg_dout7609,
   input         cfg_dout7610,
   input         cfg_dout7611,
   input         cfg_dout7612,
   input         cfg_dout7613,
   input         cfg_dout7614,
   input         cfg_dout7615,
   input         cfg_dout7616,
   input         cfg_dout7617,
   input         cfg_dout7618,
   input         cfg_dout7619,
   input         cfg_dout7620,
   input         cfg_dout7621,
   input         cfg_dout7622,
   input         cfg_dout7623,
   input         cfg_dout7624,
   input         cfg_dout7625,
   input         cfg_dout7626,
   input         cfg_dout7627,
   input         cfg_dout7628,
   input         cfg_dout7629,
   input         cfg_dout7630,
   input         cfg_dout7631,
   input         cfg_dout7632,
   input         cfg_dout7633,
   input         cfg_dout7634,
   input         cfg_dout7635,
   input         cfg_dout7636,
   input         cfg_dout7637,
   input         cfg_dout7638,
   input         cfg_dout7639,
   input         cfg_dout7640,
   input         cfg_dout7641,
   input         cfg_dout7642,
   input         cfg_dout7643,
   input         cfg_dout7644,
   input         cfg_dout7645,
   input         cfg_dout7646,
   input         cfg_dout7647,
   input         cfg_dout7648,
   input         cfg_dout7649,
   input         cfg_dout7650,
   input         cfg_dout7651,
   input         cfg_dout7652,
   input         cfg_dout7653,
   input         cfg_dout7654,
   input         cfg_dout7655,
   input         cfg_dout7656,
   input         cfg_dout7657,
   input         cfg_dout7658,
   input         cfg_dout7659,
   input         cfg_dout7660,
   input         cfg_dout7661,
   input         cfg_dout7662,
   input         cfg_dout7663,
   input         cfg_dout7664,
   input         cfg_dout7665,
   input         cfg_dout7666,
   input         cfg_dout7667,
   input         cfg_dout7668,
   input         cfg_dout7669,
   input         cfg_dout7670,
   input         cfg_dout7671,
   input         cfg_dout7672,
   input         cfg_dout7673,
   input         cfg_dout7674,
   input         cfg_dout7675,
   input         cfg_dout7676,
   input         cfg_dout7677,
   input         cfg_dout7678,
   input         cfg_dout7679,
   input         cfg_dout7680,
   input         cfg_dout7681,
   input         cfg_dout7682,
   input         cfg_dout7683,
   input         cfg_dout7684,
   input         cfg_dout7685,
   input         cfg_dout7686,
   input         cfg_dout7687,
   input         cfg_dout7688,
   input         cfg_dout7689,
   input         cfg_dout7690,
   input         cfg_dout7691,
   input         cfg_dout7692,
   input         cfg_dout7693,
   input         cfg_dout7694,
   input         cfg_dout7695,
   input         cfg_dout7696,
   input         cfg_dout7697,
   input         cfg_dout7698,
   input         cfg_dout7699,
   input         cfg_dout7700,
   input         cfg_dout7701,
   input         cfg_dout7702,
   input         cfg_dout7703,
   input         cfg_dout7704,
   input         cfg_dout7705,
   input         cfg_dout7706,
   input         cfg_dout7707,
   input         cfg_dout7708,
   input         cfg_dout7709,
   input         cfg_dout7710,
   input         cfg_dout7711,
   input         cfg_dout7712,
   input         cfg_dout7713,
   input         cfg_dout7714,
   input         cfg_dout7715,
   input         cfg_dout7716,
   input         cfg_dout7717,
   input         cfg_dout7718,
   input         cfg_dout7719,
   input         cfg_dout7720,
   input         cfg_dout7721,
   input         cfg_dout7722,
   input         cfg_dout7723,
   input         cfg_dout7724,
   input         cfg_dout7725,
   input         cfg_dout7726,
   input         cfg_dout7727,
   input         cfg_dout7728,
   input         cfg_dout7729,
   input         cfg_dout7730,
   input         cfg_dout7731,
   input         cfg_dout7732,
   input         cfg_dout7733,
   input         cfg_dout7734,
   input         cfg_dout7735,
   input         cfg_dout7736,
   input         cfg_dout7737,
   input         cfg_dout7738,
   input         cfg_dout7739,
   input         cfg_dout7740,
   input         cfg_dout7741,
   input         cfg_dout7742,
   input         cfg_dout7743,
   input         cfg_dout7744,
   input         cfg_dout7745,
   input         cfg_dout7746,
   input         cfg_dout7747,
   input         cfg_dout7748,
   input         cfg_dout7749,
   input         cfg_dout7750,
   input         cfg_dout7751,
   input         cfg_dout7752,
   input         cfg_dout7753,
   input         cfg_dout7754,
   input         cfg_dout7755,
   input         cfg_dout7756,
   input         cfg_dout7757,
   input         cfg_dout7758,
   input         cfg_dout7759,
   input         cfg_dout7760,
   input         cfg_dout7761,
   input         cfg_dout7762,
   input         cfg_dout7763,
   input         cfg_dout7764,
   input         cfg_dout7765,
   input         cfg_dout7766,
   input         cfg_dout7767,
   input         cfg_dout7768,
   input         cfg_dout7769,
   input         cfg_dout7770,
   input         cfg_dout7771,
   input         cfg_dout7772,
   input         cfg_dout7773,
   input         cfg_dout7774,
   input         cfg_dout7775,
   input         cfg_dout7776,
   input         cfg_dout7777,
   input         cfg_dout7778,
   input         cfg_dout7779,
   input         cfg_dout7780,
   input         cfg_dout7781,
   input         cfg_dout7782,
   input         cfg_dout7783,
   input         cfg_dout7784,
   input         cfg_dout7785,
   input         cfg_dout7786,
   input         cfg_dout7787,
   input         cfg_dout7788,
   input         cfg_dout7789,
   input         cfg_dout7790,
   input         cfg_dout7791,
   input         cfg_dout7792,
   input         cfg_dout7793,
   input         cfg_dout7794,
   input         cfg_dout7795,
   input         cfg_dout7796,
   input         cfg_dout7797,
   input         cfg_dout7798,
   input         cfg_dout7799,
   input         cfg_dout7800,
   input         cfg_dout7801,
   input         cfg_dout7802,
   input         cfg_dout7803,
   input         cfg_dout7804,
   input         cfg_dout7805,
   input         cfg_dout7806,
   input         cfg_dout7807,
   input         cfg_dout7808,
   input         cfg_dout7809,
   input         cfg_dout7810,
   input         cfg_dout7811,
   input         cfg_dout7812,
   input         cfg_dout7813,
   input         cfg_dout7814,
   input         cfg_dout7815,
   input         cfg_dout7816,
   input         cfg_dout7817,
   input         cfg_dout7818,
   input         cfg_dout7819,
   input         cfg_dout7820,
   input         cfg_dout7821,
   input         cfg_dout7822,
   input         cfg_dout7823,
   input         cfg_dout7824,
   input         cfg_dout7825,
   input         cfg_dout7826,
   input         cfg_dout7827,
   input         cfg_dout7828,
   input         cfg_dout7829,
   input         cfg_dout7830,
   input         cfg_dout7831,
   input         cfg_dout7832,
   input         cfg_dout7833,
   input         cfg_dout7834,
   input         cfg_dout7835,
   input         cfg_dout7836,
   input         cfg_dout7837,
   input         cfg_dout7838,
   input         cfg_dout7839,
   input         cfg_dout7840,
   input         cfg_dout7841,
   input         cfg_dout7842,
   input         cfg_dout7843,
   input         cfg_dout7844,
   input         cfg_dout7845,
   input         cfg_dout7846,
   input         cfg_dout7847,
   input         cfg_dout7848,
   input         cfg_dout7849,
   input         cfg_dout7850,
   input         cfg_dout7851,
   input         cfg_dout7852,
   input         cfg_dout7853,
   input         cfg_dout7854,
   input         cfg_dout7855,
   input         cfg_dout7856,
   input         cfg_dout7857,
   input         cfg_dout7858,
   input         cfg_dout7859,
   input         cfg_dout7860,
   input         cfg_dout7861,
   input         cfg_dout7862,
   input         cfg_dout7863,
   input         cfg_dout7864,
   input         cfg_dout7865,
   input         cfg_dout7866,
   input         cfg_dout7867,
   input         cfg_dout7868,
   input         cfg_dout7869,
   input         cfg_dout7870,
   input         cfg_dout7871,
   input         cfg_dout7872,
   input         cfg_dout7873,
   input         cfg_dout7874,
   input         cfg_dout7875,
   input         cfg_dout7876,
   input         cfg_dout7877,
   input         cfg_dout7878,
   input         cfg_dout7879,
   input         cfg_dout7880,
   input         cfg_dout7881,
   input         cfg_dout7882,
   input         cfg_dout7883,
   input         cfg_dout7884,
   input         cfg_dout7885,
   input         cfg_dout7886,
   input         cfg_dout7887,
   input         cfg_dout7888,
   input         cfg_dout7889,
   input         cfg_dout7890,
   input         cfg_dout7891,
   input         cfg_dout7892,
   input         cfg_dout7893,
   input         cfg_dout7894,
   input         cfg_dout7895,
   input         cfg_dout7896,
   input         cfg_dout7897,
   input         cfg_dout7898,
   input         cfg_dout7899,
   input         cfg_dout7900,
   input         cfg_dout7901,
   input         cfg_dout7902,
   input         cfg_dout7903,
   input         cfg_dout7904,
   input         cfg_dout7905,
   input         cfg_dout7906,
   input         cfg_dout7907,
   input         cfg_dout7908,
   input         cfg_dout7909,
   input         cfg_dout7910,
   input         cfg_dout7911,
   input         cfg_dout7912,
   input         cfg_dout7913,
   input         cfg_dout7914,
   input         cfg_dout7915,
   input         cfg_dout7916,
   input         cfg_dout7917,
   input         cfg_dout7918,
   input         cfg_dout7919,
   input         cfg_dout7920,
   input         cfg_dout7921,
   input         cfg_dout7922,
   input         cfg_dout7923,
   input         cfg_dout7924,
   input         cfg_dout7925,
   input         cfg_dout7926,
   input         cfg_dout7927,
   input         cfg_dout7928,
   input         cfg_dout7929,
   input         cfg_dout7930,
   input         cfg_dout7931,
   input         cfg_dout7932,
   input         cfg_dout7933,
   input         cfg_dout7934,
   input         cfg_dout7935,
   input         cfg_dout7936,
   input         cfg_dout7937,
   input         cfg_dout7938,
   input         cfg_dout7939,
   input         cfg_dout7940,
   input         cfg_dout7941,
   input         cfg_dout7942,
   input         cfg_dout7943,
   input         cfg_dout7944,
   input         cfg_dout7945,
   input         cfg_dout7946,
   input         cfg_dout7947,
   input         cfg_dout7948,
   input         cfg_dout7949,
   input         cfg_dout7950,
   input         cfg_dout7951,
   input         cfg_dout7952,
   input         cfg_dout7953,
   input         cfg_dout7954,
   input         cfg_dout7955,
   input         cfg_dout7956,
   input         cfg_dout7957,
   input         cfg_dout7958,
   input         cfg_dout7959,
   input         cfg_dout7960,
   input         cfg_dout7961,
   input         cfg_dout7962,
   input         cfg_dout7963,
   input         cfg_dout7964,
   input         cfg_dout7965,
   input         cfg_dout7966,
   input         cfg_dout7967,
   input         cfg_dout7968,
   input         cfg_dout7969,
   input         cfg_dout7970,
   input         cfg_dout7971,
   input         cfg_dout7972,
   input         cfg_dout7973,
   input         cfg_dout7974,
   input         cfg_dout7975,
   input         cfg_dout7976,
   input         cfg_dout7977,
   input         cfg_dout7978,
   input         cfg_dout7979,
   input         cfg_dout7980,
   input         cfg_dout7981,
   input         cfg_dout7982,
   input         cfg_dout7983,
   input         cfg_dout7984,
   input         cfg_dout7985,
   input         cfg_dout7986,
   input         cfg_dout7987,
   input         cfg_dout7988,
   input         cfg_dout7989,
   input         cfg_dout7990,
   input         cfg_dout7991,
   input         cfg_dout7992,
   input         cfg_dout7993,
   input         cfg_dout7994,
   input         cfg_dout7995,
   input         cfg_dout7996,
   input         cfg_dout7997,
   input         cfg_dout7998,
   input         cfg_dout7999,
   input         cfg_dout8000,
   input         cfg_dout8001,
   input         cfg_dout8002,
   input         cfg_dout8003,
   input         cfg_dout8004,
   input         cfg_dout8005,
   input         cfg_dout8006,
   input         cfg_dout8007,
   input         cfg_dout8008,
   input         cfg_dout8009,
   input         cfg_dout8010,
   input         cfg_dout8011,
   input         cfg_dout8012,
   input         cfg_dout8013,
   input         cfg_dout8014,
   input         cfg_dout8015,
   input         cfg_dout8016,
   input         cfg_dout8017,
   input         cfg_dout8018,
   input         cfg_dout8019,
   input         cfg_dout8020,
   input         cfg_dout8021,
   input         cfg_dout8022,
   input         cfg_dout8023,
   input         cfg_dout8024,
   input         cfg_dout8025,
   input         cfg_dout8026,
   input         cfg_dout8027,
   input         cfg_dout8028,
   input         cfg_dout8029,
   input         cfg_dout8030,
   input         cfg_dout8031,
   input         cfg_dout8032,
   input         cfg_dout8033,
   input         cfg_dout8034,
   input         cfg_dout8035,
   input         cfg_dout8036,
   input         cfg_dout8037,
   input         cfg_dout8038,
   input         cfg_dout8039,
   input         cfg_dout8040,
   input         cfg_dout8041,
   input         cfg_dout8042,
   input         cfg_dout8043,
   input         cfg_dout8044,
   input         cfg_dout8045,
   input         cfg_dout8046,
   input         cfg_dout8047,
   input         cfg_dout8048,
   input         cfg_dout8049,
   input         cfg_dout8050,
   input         cfg_dout8051,
   input         cfg_dout8052,
   input         cfg_dout8053,
   input         cfg_dout8054,
   input         cfg_dout8055,
   input         cfg_dout8056,
   input         cfg_dout8057,
   input         cfg_dout8058,
   input         cfg_dout8059,
   input         cfg_dout8060,
   input         cfg_dout8061,
   input         cfg_dout8062,
   input         cfg_dout8063,
   input         cfg_dout8064,
   input         cfg_dout8065,
   input         cfg_dout8066,
   input         cfg_dout8067,
   input         cfg_dout8068,
   input         cfg_dout8069,
   input         cfg_dout8070,
   input         cfg_dout8071,
   input         cfg_dout8072,
   input         cfg_dout8073,
   input         cfg_dout8074,
   input         cfg_dout8075,
   input         cfg_dout8076,
   input         cfg_dout8077,
   input         cfg_dout8078,
   input         cfg_dout8079,
   input         cfg_dout8080,
   input         cfg_dout8081,
   input         cfg_dout8082,
   input         cfg_dout8083,
   input         cfg_dout8084,
   input         cfg_dout8085,
   input         cfg_dout8086,
   input         cfg_dout8087,
   input         cfg_dout8088,
   input         cfg_dout8089,
   input         cfg_dout8090,
   input         cfg_dout8091,
   input         cfg_dout8092,
   input         cfg_dout8093,
   input         cfg_dout8094,
   input         cfg_dout8095,
   input         cfg_dout8096,
   input         cfg_dout8097,
   input         cfg_dout8098,
   input         cfg_dout8099,
   input         cfg_dout8100,
   input         cfg_dout8101,
   input         cfg_dout8102,
   input         cfg_dout8103,
   input         cfg_dout8104,
   input         cfg_dout8105,
   input         cfg_dout8106,
   input         cfg_dout8107,
   input         cfg_dout8108,
   input         cfg_dout8109,
   input         cfg_dout8110,
   input         cfg_dout8111,
   input         cfg_dout8112,
   input         cfg_dout8113,
   input         cfg_dout8114,
   input         cfg_dout8115,
   input         cfg_dout8116,
   input         cfg_dout8117,
   input         cfg_dout8118,
   input         cfg_dout8119,
   input         cfg_dout8120,
   input         cfg_dout8121,
   input         cfg_dout8122,
   input         cfg_dout8123,
   input         cfg_dout8124,
   input         cfg_dout8125,
   input         cfg_dout8126,
   input         cfg_dout8127,
   input         cfg_dout8128,
   input         cfg_dout8129,
   input         cfg_dout8130,
   input         cfg_dout8131,
   input         cfg_dout8132,
   input         cfg_dout8133,
   input         cfg_dout8134,
   input         cfg_dout8135,
   input         cfg_dout8136,
   input         cfg_dout8137,
   input         cfg_dout8138,
   input         cfg_dout8139,
   input         cfg_dout8140,
   input         cfg_dout8141,
   input         cfg_dout8142,
   input         cfg_dout8143,
   input         cfg_dout8144,
   input         cfg_dout8145,
   input         cfg_dout8146,
   input         cfg_dout8147,
   input         cfg_dout8148,
   input         cfg_dout8149,
   input         cfg_dout8150,
   input         cfg_dout8151,
   input         cfg_dout8152,
   input         cfg_dout8153,
   input         cfg_dout8154,
   input         cfg_dout8155,
   input         cfg_dout8156,
   input         cfg_dout8157,
   input         cfg_dout8158,
   input         cfg_dout8159,
   input         cfg_dout8160,
   input         cfg_dout8161,
   input         cfg_dout8162,
   input         cfg_dout8163,
   input         cfg_dout8164,
   input         cfg_dout8165,
   input         cfg_dout8166,
   input         cfg_dout8167,
   input         cfg_dout8168,
   input         cfg_dout8169,
   input         cfg_dout8170,
   input         cfg_dout8171,
   input         cfg_dout8172,
   input         cfg_dout8173,
   input         cfg_dout8174,
   input         cfg_dout8175,
   input         cfg_dout8176,
   input         cfg_dout8177,
   input         cfg_dout8178,
   input         cfg_dout8179,
   input         cfg_dout8180,
   input         cfg_dout8181,
   input         cfg_dout8182,
   input         cfg_dout8183,
   input         cfg_dout8184,
   input         cfg_dout8185,
   input         cfg_dout8186,
   input         cfg_dout8187,
   input         cfg_dout8188,
   input         cfg_dout8189,
   input         cfg_dout8190,
   input         cfg_dout8191,
   input         tc_cfg_dout,
   input         cc_cfg_dout0,
   input         cc_cfg_dout1,
   input         cc_cfg_dout2,
   input         cc_cfg_dout3,
   input         match_out0,
   input         match_out1,
   input         match_out2,
   input         match_out3,
   input         match_out4,
   input         match_out5,
   input         match_out6,
   input         match_out7,
   input         match_out8,
   input         match_out9,
   input         match_out10,
   input         match_out11,
   input         match_out12,
   input         match_out13,
   input         match_out14,
   input         match_out15,
   input         match_out16,
   input         match_out17,
   input         match_out18,
   input         match_out19,
   input         match_out20,
   input         match_out21,
   input         match_out22,
   input         match_out23,
   input         match_out24,
   input         match_out25,
   input         match_out26,
   input         match_out27,
   input         match_out28,
   input         match_out29,
   input         match_out30,
   input         match_out31,
   input         match_out32,
   input         match_out33,
   input         match_out34,
   input         match_out35,
   input         match_out36,
   input         match_out37,
   input         match_out38,
   input         match_out39,
   input         match_out40,
   input         match_out41,
   input         match_out42,
   input         match_out43,
   input         match_out44,
   input         match_out45,
   input         match_out46,
   input         match_out47,
   input         match_out48,
   input         match_out49,
   input         match_out50,
   input         match_out51,
   input         match_out52,
   input         match_out53,
   input         match_out54,
   input         match_out55,
   input         match_out56,
   input         match_out57,
   input         match_out58,
   input         match_out59,
   input         match_out60,
   input         match_out61,
   input         match_out62,
   input         match_out63,
   input         match_out64,
   input         match_out65,
   input         match_out66,
   input         match_out67,
   input         match_out68,
   input         match_out69,
   input         match_out70,
   input         match_out71,
   input         match_out72,
   input         match_out73,
   input         match_out74,
   input         match_out75,
   input         match_out76,
   input         match_out77,
   input         match_out78,
   input         match_out79,
   input         match_out80,
   input         match_out81,
   input         match_out82,
   input         match_out83,
   input         match_out84,
   input         match_out85,
   input         match_out86,
   input         match_out87,
   input         match_out88,
   input         match_out89,
   input         match_out90,
   input         match_out91,
   input         match_out92,
   input         match_out93,
   input         match_out94,
   input         match_out95,
   input         match_out96,
   input         match_out97,
   input         match_out98,
   input         match_out99,
   input         match_out100,
   input         match_out101,
   input         match_out102,
   input         match_out103,
   input         match_out104,
   input         match_out105,
   input         match_out106,
   input         match_out107,
   input         match_out108,
   input         match_out109,
   input         match_out110,
   input         match_out111,
   input         match_out112,
   input         match_out113,
   input         match_out114,
   input         match_out115,
   input         match_out116,
   input         match_out117,
   input         match_out118,
   input         match_out119,
   input         match_out120,
   input         match_out121,
   input         match_out122,
   input         match_out123,
   input         match_out124,
   input         match_out125,
   input         match_out126,
   input         match_out127,
   input         match_out128,
   input         match_out129,
   input         match_out130,
   input         match_out131,
   input         match_out132,
   input         match_out133,
   input         match_out134,
   input         match_out135,
   input         match_out136,
   input         match_out137,
   input         match_out138,
   input         match_out139,
   input         match_out140,
   input         match_out141,
   input         match_out142,
   input         match_out143,
   input         match_out144,
   input         match_out145,
   input         match_out146,
   input         match_out147,
   input         match_out148,
   input         match_out149,
   input         match_out150,
   input         match_out151,
   input         match_out152,
   input         match_out153,
   input         match_out154,
   input         match_out155,
   input         match_out156,
   input         match_out157,
   input         match_out158,
   input         match_out159,
   input         match_out160,
   input         match_out161,
   input         match_out162,
   input         match_out163,
   input         match_out164,
   input         match_out165,
   input         match_out166,
   input         match_out167,
   input         match_out168,
   input         match_out169,
   input         match_out170,
   input         match_out171,
   input         match_out172,
   input         match_out173,
   input         match_out174,
   input         match_out175,
   input         match_out176,
   input         match_out177,
   input         match_out178,
   input         match_out179,
   input         match_out180,
   input         match_out181,
   input         match_out182,
   input         match_out183,
   input         match_out184,
   input         match_out185,
   input         match_out186,
   input         match_out187,
   input         match_out188,
   input         match_out189,
   input         match_out190,
   input         match_out191,
   input         match_out192,
   input         match_out193,
   input         match_out194,
   input         match_out195,
   input         match_out196,
   input         match_out197,
   input         match_out198,
   input         match_out199,
   input         match_out200,
   input         match_out201,
   input         match_out202,
   input         match_out203,
   input         match_out204,
   input         match_out205,
   input         match_out206,
   input         match_out207,
   input         match_out208,
   input         match_out209,
   input         match_out210,
   input         match_out211,
   input         match_out212,
   input         match_out213,
   input         match_out214,
   input         match_out215,
   input         match_out216,
   input         match_out217,
   input         match_out218,
   input         match_out219,
   input         match_out220,
   input         match_out221,
   input         match_out222,
   input         match_out223,
   input         match_out224,
   input         match_out225,
   input         match_out226,
   input         match_out227,
   input         match_out228,
   input         match_out229,
   input         match_out230,
   input         match_out231,
   input         match_out232,
   input         match_out233,
   input         match_out234,
   input         match_out235,
   input         match_out236,
   input         match_out237,
   input         match_out238,
   input         match_out239,
   input         match_out240,
   input         match_out241,
   input         match_out242,
   input         match_out243,
   input         match_out244,
   input         match_out245,
   input         match_out246,
   input         match_out247,
   input         match_out248,
   input         match_out249,
   input         match_out250,
   input         match_out251,
   input         match_out252,
   input         match_out253,
   input         match_out254,
   input         match_out255,
   input         match_out256,
   input         match_out257,
   input         match_out258,
   input         match_out259,
   input         match_out260,
   input         match_out261,
   input         match_out262,
   input         match_out263,
   input         match_out264,
   input         match_out265,
   input         match_out266,
   input         match_out267,
   input         match_out268,
   input         match_out269,
   input         match_out270,
   input         match_out271,
   input         match_out272,
   input         match_out273,
   input         match_out274,
   input         match_out275,
   input         match_out276,
   input         match_out277,
   input         match_out278,
   input         match_out279,
   input         match_out280,
   input         match_out281,
   input         match_out282,
   input         match_out283,
   input         match_out284,
   input         match_out285,
   input         match_out286,
   input         match_out287,
   input         match_out288,
   input         match_out289,
   input         match_out290,
   input         match_out291,
   input         match_out292,
   input         match_out293,
   input         match_out294,
   input         match_out295,
   input         match_out296,
   input         match_out297,
   input         match_out298,
   input         match_out299,
   input         match_out300,
   input         match_out301,
   input         match_out302,
   input         match_out303,
   input         match_out304,
   input         match_out305,
   input         match_out306,
   input         match_out307,
   input         match_out308,
   input         match_out309,
   input         match_out310,
   input         match_out311,
   input         match_out312,
   input         match_out313,
   input         match_out314,
   input         match_out315,
   input         match_out316,
   input         match_out317,
   input         match_out318,
   input         match_out319,
   input         match_out320,
   input         match_out321,
   input         match_out322,
   input         match_out323,
   input         match_out324,
   input         match_out325,
   input         match_out326,
   input         match_out327,
   input         match_out328,
   input         match_out329,
   input         match_out330,
   input         match_out331,
   input         match_out332,
   input         match_out333,
   input         match_out334,
   input         match_out335,
   input         match_out336,
   input         match_out337,
   input         match_out338,
   input         match_out339,
   input         match_out340,
   input         match_out341,
   input         match_out342,
   input         match_out343,
   input         match_out344,
   input         match_out345,
   input         match_out346,
   input         match_out347,
   input         match_out348,
   input         match_out349,
   input         match_out350,
   input         match_out351,
   input         match_out352,
   input         match_out353,
   input         match_out354,
   input         match_out355,
   input         match_out356,
   input         match_out357,
   input         match_out358,
   input         match_out359,
   input         match_out360,
   input         match_out361,
   input         match_out362,
   input         match_out363,
   input         match_out364,
   input         match_out365,
   input         match_out366,
   input         match_out367,
   input         match_out368,
   input         match_out369,
   input         match_out370,
   input         match_out371,
   input         match_out372,
   input         match_out373,
   input         match_out374,
   input         match_out375,
   input         match_out376,
   input         match_out377,
   input         match_out378,
   input         match_out379,
   input         match_out380,
   input         match_out381,
   input         match_out382,
   input         match_out383,
   input         match_out384,
   input         match_out385,
   input         match_out386,
   input         match_out387,
   input         match_out388,
   input         match_out389,
   input         match_out390,
   input         match_out391,
   input         match_out392,
   input         match_out393,
   input         match_out394,
   input         match_out395,
   input         match_out396,
   input         match_out397,
   input         match_out398,
   input         match_out399,
   input         match_out400,
   input         match_out401,
   input         match_out402,
   input         match_out403,
   input         match_out404,
   input         match_out405,
   input         match_out406,
   input         match_out407,
   input         match_out408,
   input         match_out409,
   input         match_out410,
   input         match_out411,
   input         match_out412,
   input         match_out413,
   input         match_out414,
   input         match_out415,
   input         match_out416,
   input         match_out417,
   input         match_out418,
   input         match_out419,
   input         match_out420,
   input         match_out421,
   input         match_out422,
   input         match_out423,
   input         match_out424,
   input         match_out425,
   input         match_out426,
   input         match_out427,
   input         match_out428,
   input         match_out429,
   input         match_out430,
   input         match_out431,
   input         match_out432,
   input         match_out433,
   input         match_out434,
   input         match_out435,
   input         match_out436,
   input         match_out437,
   input         match_out438,
   input         match_out439,
   input         match_out440,
   input         match_out441,
   input         match_out442,
   input         match_out443,
   input         match_out444,
   input         match_out445,
   input         match_out446,
   input         match_out447,
   input         match_out448,
   input         match_out449,
   input         match_out450,
   input         match_out451,
   input         match_out452,
   input         match_out453,
   input         match_out454,
   input         match_out455,
   input         match_out456,
   input         match_out457,
   input         match_out458,
   input         match_out459,
   input         match_out460,
   input         match_out461,
   input         match_out462,
   input         match_out463,
   input         match_out464,
   input         match_out465,
   input         match_out466,
   input         match_out467,
   input         match_out468,
   input         match_out469,
   input         match_out470,
   input         match_out471,
   input         match_out472,
   input         match_out473,
   input         match_out474,
   input         match_out475,
   input         match_out476,
   input         match_out477,
   input         match_out478,
   input         match_out479,
   input         match_out480,
   input         match_out481,
   input         match_out482,
   input         match_out483,
   input         match_out484,
   input         match_out485,
   input         match_out486,
   input         match_out487,
   input         match_out488,
   input         match_out489,
   input         match_out490,
   input         match_out491,
   input         match_out492,
   input         match_out493,
   input         match_out494,
   input         match_out495,
   input         match_out496,
   input         match_out497,
   input         match_out498,
   input         match_out499,
   input         match_out500,
   input         match_out501,
   input         match_out502,
   input         match_out503,
   input         match_out504,
   input         match_out505,
   input         match_out506,
   input         match_out507,
   input         match_out508,
   input         match_out509,
   input         match_out510,
   input         match_out511,
   input         match_out512,
   input         match_out513,
   input         match_out514,
   input         match_out515,
   input         match_out516,
   input         match_out517,
   input         match_out518,
   input         match_out519,
   input         match_out520,
   input         match_out521,
   input         match_out522,
   input         match_out523,
   input         match_out524,
   input         match_out525,
   input         match_out526,
   input         match_out527,
   input         match_out528,
   input         match_out529,
   input         match_out530,
   input         match_out531,
   input         match_out532,
   input         match_out533,
   input         match_out534,
   input         match_out535,
   input         match_out536,
   input         match_out537,
   input         match_out538,
   input         match_out539,
   input         match_out540,
   input         match_out541,
   input         match_out542,
   input         match_out543,
   input         match_out544,
   input         match_out545,
   input         match_out546,
   input         match_out547,
   input         match_out548,
   input         match_out549,
   input         match_out550,
   input         match_out551,
   input         match_out552,
   input         match_out553,
   input         match_out554,
   input         match_out555,
   input         match_out556,
   input         match_out557,
   input         match_out558,
   input         match_out559,
   input         match_out560,
   input         match_out561,
   input         match_out562,
   input         match_out563,
   input         match_out564,
   input         match_out565,
   input         match_out566,
   input         match_out567,
   input         match_out568,
   input         match_out569,
   input         match_out570,
   input         match_out571,
   input         match_out572,
   input         match_out573,
   input         match_out574,
   input         match_out575,
   input         match_out576,
   input         match_out577,
   input         match_out578,
   input         match_out579,
   input         match_out580,
   input         match_out581,
   input         match_out582,
   input         match_out583,
   input         match_out584,
   input         match_out585,
   input         match_out586,
   input         match_out587,
   input         match_out588,
   input         match_out589,
   input         match_out590,
   input         match_out591,
   input         match_out592,
   input         match_out593,
   input         match_out594,
   input         match_out595,
   input         match_out596,
   input         match_out597,
   input         match_out598,
   input         match_out599,
   input         match_out600,
   input         match_out601,
   input         match_out602,
   input         match_out603,
   input         match_out604,
   input         match_out605,
   input         match_out606,
   input         match_out607,
   input         match_out608,
   input         match_out609,
   input         match_out610,
   input         match_out611,
   input         match_out612,
   input         match_out613,
   input         match_out614,
   input         match_out615,
   input         match_out616,
   input         match_out617,
   input         match_out618,
   input         match_out619,
   input         match_out620,
   input         match_out621,
   input         match_out622,
   input         match_out623,
   input         match_out624,
   input         match_out625,
   input         match_out626,
   input         match_out627,
   input         match_out628,
   input         match_out629,
   input         match_out630,
   input         match_out631,
   input         match_out632,
   input         match_out633,
   input         match_out634,
   input         match_out635,
   input         match_out636,
   input         match_out637,
   input         match_out638,
   input         match_out639,
   input         match_out640,
   input         match_out641,
   input         match_out642,
   input         match_out643,
   input         match_out644,
   input         match_out645,
   input         match_out646,
   input         match_out647,
   input         match_out648,
   input         match_out649,
   input         match_out650,
   input         match_out651,
   input         match_out652,
   input         match_out653,
   input         match_out654,
   input         match_out655,
   input         match_out656,
   input         match_out657,
   input         match_out658,
   input         match_out659,
   input         match_out660,
   input         match_out661,
   input         match_out662,
   input         match_out663,
   input         match_out664,
   input         match_out665,
   input         match_out666,
   input         match_out667,
   input         match_out668,
   input         match_out669,
   input         match_out670,
   input         match_out671,
   input         match_out672,
   input         match_out673,
   input         match_out674,
   input         match_out675,
   input         match_out676,
   input         match_out677,
   input         match_out678,
   input         match_out679,
   input         match_out680,
   input         match_out681,
   input         match_out682,
   input         match_out683,
   input         match_out684,
   input         match_out685,
   input         match_out686,
   input         match_out687,
   input         match_out688,
   input         match_out689,
   input         match_out690,
   input         match_out691,
   input         match_out692,
   input         match_out693,
   input         match_out694,
   input         match_out695,
   input         match_out696,
   input         match_out697,
   input         match_out698,
   input         match_out699,
   input         match_out700,
   input         match_out701,
   input         match_out702,
   input         match_out703,
   input         match_out704,
   input         match_out705,
   input         match_out706,
   input         match_out707,
   input         match_out708,
   input         match_out709,
   input         match_out710,
   input         match_out711,
   input         match_out712,
   input         match_out713,
   input         match_out714,
   input         match_out715,
   input         match_out716,
   input         match_out717,
   input         match_out718,
   input         match_out719,
   input         match_out720,
   input         match_out721,
   input         match_out722,
   input         match_out723,
   input         match_out724,
   input         match_out725,
   input         match_out726,
   input         match_out727,
   input         match_out728,
   input         match_out729,
   input         match_out730,
   input         match_out731,
   input         match_out732,
   input         match_out733,
   input         match_out734,
   input         match_out735,
   input         match_out736,
   input         match_out737,
   input         match_out738,
   input         match_out739,
   input         match_out740,
   input         match_out741,
   input         match_out742,
   input         match_out743,
   input         match_out744,
   input         match_out745,
   input         match_out746,
   input         match_out747,
   input         match_out748,
   input         match_out749,
   input         match_out750,
   input         match_out751,
   input         match_out752,
   input         match_out753,
   input         match_out754,
   input         match_out755,
   input         match_out756,
   input         match_out757,
   input         match_out758,
   input         match_out759,
   input         match_out760,
   input         match_out761,
   input         match_out762,
   input         match_out763,
   input         match_out764,
   input         match_out765,
   input         match_out766,
   input         match_out767,
   input         match_out768,
   input         match_out769,
   input         match_out770,
   input         match_out771,
   input         match_out772,
   input         match_out773,
   input         match_out774,
   input         match_out775,
   input         match_out776,
   input         match_out777,
   input         match_out778,
   input         match_out779,
   input         match_out780,
   input         match_out781,
   input         match_out782,
   input         match_out783,
   input         match_out784,
   input         match_out785,
   input         match_out786,
   input         match_out787,
   input         match_out788,
   input         match_out789,
   input         match_out790,
   input         match_out791,
   input         match_out792,
   input         match_out793,
   input         match_out794,
   input         match_out795,
   input         match_out796,
   input         match_out797,
   input         match_out798,
   input         match_out799,
   input         match_out800,
   input         match_out801,
   input         match_out802,
   input         match_out803,
   input         match_out804,
   input         match_out805,
   input         match_out806,
   input         match_out807,
   input         match_out808,
   input         match_out809,
   input         match_out810,
   input         match_out811,
   input         match_out812,
   input         match_out813,
   input         match_out814,
   input         match_out815,
   input         match_out816,
   input         match_out817,
   input         match_out818,
   input         match_out819,
   input         match_out820,
   input         match_out821,
   input         match_out822,
   input         match_out823,
   input         match_out824,
   input         match_out825,
   input         match_out826,
   input         match_out827,
   input         match_out828,
   input         match_out829,
   input         match_out830,
   input         match_out831,
   input         match_out832,
   input         match_out833,
   input         match_out834,
   input         match_out835,
   input         match_out836,
   input         match_out837,
   input         match_out838,
   input         match_out839,
   input         match_out840,
   input         match_out841,
   input         match_out842,
   input         match_out843,
   input         match_out844,
   input         match_out845,
   input         match_out846,
   input         match_out847,
   input         match_out848,
   input         match_out849,
   input         match_out850,
   input         match_out851,
   input         match_out852,
   input         match_out853,
   input         match_out854,
   input         match_out855,
   input         match_out856,
   input         match_out857,
   input         match_out858,
   input         match_out859,
   input         match_out860,
   input         match_out861,
   input         match_out862,
   input         match_out863,
   input         match_out864,
   input         match_out865,
   input         match_out866,
   input         match_out867,
   input         match_out868,
   input         match_out869,
   input         match_out870,
   input         match_out871,
   input         match_out872,
   input         match_out873,
   input         match_out874,
   input         match_out875,
   input         match_out876,
   input         match_out877,
   input         match_out878,
   input         match_out879,
   input         match_out880,
   input         match_out881,
   input         match_out882,
   input         match_out883,
   input         match_out884,
   input         match_out885,
   input         match_out886,
   input         match_out887,
   input         match_out888,
   input         match_out889,
   input         match_out890,
   input         match_out891,
   input         match_out892,
   input         match_out893,
   input         match_out894,
   input         match_out895,
   input         match_out896,
   input         match_out897,
   input         match_out898,
   input         match_out899,
   input         match_out900,
   input         match_out901,
   input         match_out902,
   input         match_out903,
   input         match_out904,
   input         match_out905,
   input         match_out906,
   input         match_out907,
   input         match_out908,
   input         match_out909,
   input         match_out910,
   input         match_out911,
   input         match_out912,
   input         match_out913,
   input         match_out914,
   input         match_out915,
   input         match_out916,
   input         match_out917,
   input         match_out918,
   input         match_out919,
   input         match_out920,
   input         match_out921,
   input         match_out922,
   input         match_out923,
   input         match_out924,
   input         match_out925,
   input         match_out926,
   input         match_out927,
   input         match_out928,
   input         match_out929,
   input         match_out930,
   input         match_out931,
   input         match_out932,
   input         match_out933,
   input         match_out934,
   input         match_out935,
   input         match_out936,
   input         match_out937,
   input         match_out938,
   input         match_out939,
   input         match_out940,
   input         match_out941,
   input         match_out942,
   input         match_out943,
   input         match_out944,
   input         match_out945,
   input         match_out946,
   input         match_out947,
   input         match_out948,
   input         match_out949,
   input         match_out950,
   input         match_out951,
   input         match_out952,
   input         match_out953,
   input         match_out954,
   input         match_out955,
   input         match_out956,
   input         match_out957,
   input         match_out958,
   input         match_out959,
   input         match_out960,
   input         match_out961,
   input         match_out962,
   input         match_out963,
   input         match_out964,
   input         match_out965,
   input         match_out966,
   input         match_out967,
   input         match_out968,
   input         match_out969,
   input         match_out970,
   input         match_out971,
   input         match_out972,
   input         match_out973,
   input         match_out974,
   input         match_out975,
   input         match_out976,
   input         match_out977,
   input         match_out978,
   input         match_out979,
   input         match_out980,
   input         match_out981,
   input         match_out982,
   input         match_out983,
   input         match_out984,
   input         match_out985,
   input         match_out986,
   input         match_out987,
   input         match_out988,
   input         match_out989,
   input         match_out990,
   input         match_out991,
   input         match_out992,
   input         match_out993,
   input         match_out994,
   input         match_out995,
   input         match_out996,
   input         match_out997,
   input         match_out998,
   input         match_out999,
   input         match_out1000,
   input         match_out1001,
   input         match_out1002,
   input         match_out1003,
   input         match_out1004,
   input         match_out1005,
   input         match_out1006,
   input         match_out1007,
   input         match_out1008,
   input         match_out1009,
   input         match_out1010,
   input         match_out1011,
   input         match_out1012,
   input         match_out1013,
   input         match_out1014,
   input         match_out1015,
   input         match_out1016,
   input         match_out1017,
   input         match_out1018,
   input         match_out1019,
   input         match_out1020,
   input         match_out1021,
   input         match_out1022,
   input         match_out1023,
   input         match_out1024,
   input         match_out1025,
   input         match_out1026,
   input         match_out1027,
   input         match_out1028,
   input         match_out1029,
   input         match_out1030,
   input         match_out1031,
   input         match_out1032,
   input         match_out1033,
   input         match_out1034,
   input         match_out1035,
   input         match_out1036,
   input         match_out1037,
   input         match_out1038,
   input         match_out1039,
   input         match_out1040,
   input         match_out1041,
   input         match_out1042,
   input         match_out1043,
   input         match_out1044,
   input         match_out1045,
   input         match_out1046,
   input         match_out1047,
   input         match_out1048,
   input         match_out1049,
   input         match_out1050,
   input         match_out1051,
   input         match_out1052,
   input         match_out1053,
   input         match_out1054,
   input         match_out1055,
   input         match_out1056,
   input         match_out1057,
   input         match_out1058,
   input         match_out1059,
   input         match_out1060,
   input         match_out1061,
   input         match_out1062,
   input         match_out1063,
   input         match_out1064,
   input         match_out1065,
   input         match_out1066,
   input         match_out1067,
   input         match_out1068,
   input         match_out1069,
   input         match_out1070,
   input         match_out1071,
   input         match_out1072,
   input         match_out1073,
   input         match_out1074,
   input         match_out1075,
   input         match_out1076,
   input         match_out1077,
   input         match_out1078,
   input         match_out1079,
   input         match_out1080,
   input         match_out1081,
   input         match_out1082,
   input         match_out1083,
   input         match_out1084,
   input         match_out1085,
   input         match_out1086,
   input         match_out1087,
   input         match_out1088,
   input         match_out1089,
   input         match_out1090,
   input         match_out1091,
   input         match_out1092,
   input         match_out1093,
   input         match_out1094,
   input         match_out1095,
   input         match_out1096,
   input         match_out1097,
   input         match_out1098,
   input         match_out1099,
   input         match_out1100,
   input         match_out1101,
   input         match_out1102,
   input         match_out1103,
   input         match_out1104,
   input         match_out1105,
   input         match_out1106,
   input         match_out1107,
   input         match_out1108,
   input         match_out1109,
   input         match_out1110,
   input         match_out1111,
   input         match_out1112,
   input         match_out1113,
   input         match_out1114,
   input         match_out1115,
   input         match_out1116,
   input         match_out1117,
   input         match_out1118,
   input         match_out1119,
   input         match_out1120,
   input         match_out1121,
   input         match_out1122,
   input         match_out1123,
   input         match_out1124,
   input         match_out1125,
   input         match_out1126,
   input         match_out1127,
   input         match_out1128,
   input         match_out1129,
   input         match_out1130,
   input         match_out1131,
   input         match_out1132,
   input         match_out1133,
   input         match_out1134,
   input         match_out1135,
   input         match_out1136,
   input         match_out1137,
   input         match_out1138,
   input         match_out1139,
   input         match_out1140,
   input         match_out1141,
   input         match_out1142,
   input         match_out1143,
   input         match_out1144,
   input         match_out1145,
   input         match_out1146,
   input         match_out1147,
   input         match_out1148,
   input         match_out1149,
   input         match_out1150,
   input         match_out1151,
   input         match_out1152,
   input         match_out1153,
   input         match_out1154,
   input         match_out1155,
   input         match_out1156,
   input         match_out1157,
   input         match_out1158,
   input         match_out1159,
   input         match_out1160,
   input         match_out1161,
   input         match_out1162,
   input         match_out1163,
   input         match_out1164,
   input         match_out1165,
   input         match_out1166,
   input         match_out1167,
   input         match_out1168,
   input         match_out1169,
   input         match_out1170,
   input         match_out1171,
   input         match_out1172,
   input         match_out1173,
   input         match_out1174,
   input         match_out1175,
   input         match_out1176,
   input         match_out1177,
   input         match_out1178,
   input         match_out1179,
   input         match_out1180,
   input         match_out1181,
   input         match_out1182,
   input         match_out1183,
   input         match_out1184,
   input         match_out1185,
   input         match_out1186,
   input         match_out1187,
   input         match_out1188,
   input         match_out1189,
   input         match_out1190,
   input         match_out1191,
   input         match_out1192,
   input         match_out1193,
   input         match_out1194,
   input         match_out1195,
   input         match_out1196,
   input         match_out1197,
   input         match_out1198,
   input         match_out1199,
   input         match_out1200,
   input         match_out1201,
   input         match_out1202,
   input         match_out1203,
   input         match_out1204,
   input         match_out1205,
   input         match_out1206,
   input         match_out1207,
   input         match_out1208,
   input         match_out1209,
   input         match_out1210,
   input         match_out1211,
   input         match_out1212,
   input         match_out1213,
   input         match_out1214,
   input         match_out1215,
   input         match_out1216,
   input         match_out1217,
   input         match_out1218,
   input         match_out1219,
   input         match_out1220,
   input         match_out1221,
   input         match_out1222,
   input         match_out1223,
   input         match_out1224,
   input         match_out1225,
   input         match_out1226,
   input         match_out1227,
   input         match_out1228,
   input         match_out1229,
   input         match_out1230,
   input         match_out1231,
   input         match_out1232,
   input         match_out1233,
   input         match_out1234,
   input         match_out1235,
   input         match_out1236,
   input         match_out1237,
   input         match_out1238,
   input         match_out1239,
   input         match_out1240,
   input         match_out1241,
   input         match_out1242,
   input         match_out1243,
   input         match_out1244,
   input         match_out1245,
   input         match_out1246,
   input         match_out1247,
   input         match_out1248,
   input         match_out1249,
   input         match_out1250,
   input         match_out1251,
   input         match_out1252,
   input         match_out1253,
   input         match_out1254,
   input         match_out1255,
   input         match_out1256,
   input         match_out1257,
   input         match_out1258,
   input         match_out1259,
   input         match_out1260,
   input         match_out1261,
   input         match_out1262,
   input         match_out1263,
   input         match_out1264,
   input         match_out1265,
   input         match_out1266,
   input         match_out1267,
   input         match_out1268,
   input         match_out1269,
   input         match_out1270,
   input         match_out1271,
   input         match_out1272,
   input         match_out1273,
   input         match_out1274,
   input         match_out1275,
   input         match_out1276,
   input         match_out1277,
   input         match_out1278,
   input         match_out1279,
   input         match_out1280,
   input         match_out1281,
   input         match_out1282,
   input         match_out1283,
   input         match_out1284,
   input         match_out1285,
   input         match_out1286,
   input         match_out1287,
   input         match_out1288,
   input         match_out1289,
   input         match_out1290,
   input         match_out1291,
   input         match_out1292,
   input         match_out1293,
   input         match_out1294,
   input         match_out1295,
   input         match_out1296,
   input         match_out1297,
   input         match_out1298,
   input         match_out1299,
   input         match_out1300,
   input         match_out1301,
   input         match_out1302,
   input         match_out1303,
   input         match_out1304,
   input         match_out1305,
   input         match_out1306,
   input         match_out1307,
   input         match_out1308,
   input         match_out1309,
   input         match_out1310,
   input         match_out1311,
   input         match_out1312,
   input         match_out1313,
   input         match_out1314,
   input         match_out1315,
   input         match_out1316,
   input         match_out1317,
   input         match_out1318,
   input         match_out1319,
   input         match_out1320,
   input         match_out1321,
   input         match_out1322,
   input         match_out1323,
   input         match_out1324,
   input         match_out1325,
   input         match_out1326,
   input         match_out1327,
   input         match_out1328,
   input         match_out1329,
   input         match_out1330,
   input         match_out1331,
   input         match_out1332,
   input         match_out1333,
   input         match_out1334,
   input         match_out1335,
   input         match_out1336,
   input         match_out1337,
   input         match_out1338,
   input         match_out1339,
   input         match_out1340,
   input         match_out1341,
   input         match_out1342,
   input         match_out1343,
   input         match_out1344,
   input         match_out1345,
   input         match_out1346,
   input         match_out1347,
   input         match_out1348,
   input         match_out1349,
   input         match_out1350,
   input         match_out1351,
   input         match_out1352,
   input         match_out1353,
   input         match_out1354,
   input         match_out1355,
   input         match_out1356,
   input         match_out1357,
   input         match_out1358,
   input         match_out1359,
   input         match_out1360,
   input         match_out1361,
   input         match_out1362,
   input         match_out1363,
   input         match_out1364,
   input         match_out1365,
   input         match_out1366,
   input         match_out1367,
   input         match_out1368,
   input         match_out1369,
   input         match_out1370,
   input         match_out1371,
   input         match_out1372,
   input         match_out1373,
   input         match_out1374,
   input         match_out1375,
   input         match_out1376,
   input         match_out1377,
   input         match_out1378,
   input         match_out1379,
   input         match_out1380,
   input         match_out1381,
   input         match_out1382,
   input         match_out1383,
   input         match_out1384,
   input         match_out1385,
   input         match_out1386,
   input         match_out1387,
   input         match_out1388,
   input         match_out1389,
   input         match_out1390,
   input         match_out1391,
   input         match_out1392,
   input         match_out1393,
   input         match_out1394,
   input         match_out1395,
   input         match_out1396,
   input         match_out1397,
   input         match_out1398,
   input         match_out1399,
   input         match_out1400,
   input         match_out1401,
   input         match_out1402,
   input         match_out1403,
   input         match_out1404,
   input         match_out1405,
   input         match_out1406,
   input         match_out1407,
   input         match_out1408,
   input         match_out1409,
   input         match_out1410,
   input         match_out1411,
   input         match_out1412,
   input         match_out1413,
   input         match_out1414,
   input         match_out1415,
   input         match_out1416,
   input         match_out1417,
   input         match_out1418,
   input         match_out1419,
   input         match_out1420,
   input         match_out1421,
   input         match_out1422,
   input         match_out1423,
   input         match_out1424,
   input         match_out1425,
   input         match_out1426,
   input         match_out1427,
   input         match_out1428,
   input         match_out1429,
   input         match_out1430,
   input         match_out1431,
   input         match_out1432,
   input         match_out1433,
   input         match_out1434,
   input         match_out1435,
   input         match_out1436,
   input         match_out1437,
   input         match_out1438,
   input         match_out1439,
   input         match_out1440,
   input         match_out1441,
   input         match_out1442,
   input         match_out1443,
   input         match_out1444,
   input         match_out1445,
   input         match_out1446,
   input         match_out1447,
   input         match_out1448,
   input         match_out1449,
   input         match_out1450,
   input         match_out1451,
   input         match_out1452,
   input         match_out1453,
   input         match_out1454,
   input         match_out1455,
   input         match_out1456,
   input         match_out1457,
   input         match_out1458,
   input         match_out1459,
   input         match_out1460,
   input         match_out1461,
   input         match_out1462,
   input         match_out1463,
   input         match_out1464,
   input         match_out1465,
   input         match_out1466,
   input         match_out1467,
   input         match_out1468,
   input         match_out1469,
   input         match_out1470,
   input         match_out1471,
   input         match_out1472,
   input         match_out1473,
   input         match_out1474,
   input         match_out1475,
   input         match_out1476,
   input         match_out1477,
   input         match_out1478,
   input         match_out1479,
   input         match_out1480,
   input         match_out1481,
   input         match_out1482,
   input         match_out1483,
   input         match_out1484,
   input         match_out1485,
   input         match_out1486,
   input         match_out1487,
   input         match_out1488,
   input         match_out1489,
   input         match_out1490,
   input         match_out1491,
   input         match_out1492,
   input         match_out1493,
   input         match_out1494,
   input         match_out1495,
   input         match_out1496,
   input         match_out1497,
   input         match_out1498,
   input         match_out1499,
   input         match_out1500,
   input         match_out1501,
   input         match_out1502,
   input         match_out1503,
   input         match_out1504,
   input         match_out1505,
   input         match_out1506,
   input         match_out1507,
   input         match_out1508,
   input         match_out1509,
   input         match_out1510,
   input         match_out1511,
   input         match_out1512,
   input         match_out1513,
   input         match_out1514,
   input         match_out1515,
   input         match_out1516,
   input         match_out1517,
   input         match_out1518,
   input         match_out1519,
   input         match_out1520,
   input         match_out1521,
   input         match_out1522,
   input         match_out1523,
   input         match_out1524,
   input         match_out1525,
   input         match_out1526,
   input         match_out1527,
   input         match_out1528,
   input         match_out1529,
   input         match_out1530,
   input         match_out1531,
   input         match_out1532,
   input         match_out1533,
   input         match_out1534,
   input         match_out1535,
   input         match_out1536,
   input         match_out1537,
   input         match_out1538,
   input         match_out1539,
   input         match_out1540,
   input         match_out1541,
   input         match_out1542,
   input         match_out1543,
   input         match_out1544,
   input         match_out1545,
   input         match_out1546,
   input         match_out1547,
   input         match_out1548,
   input         match_out1549,
   input         match_out1550,
   input         match_out1551,
   input         match_out1552,
   input         match_out1553,
   input         match_out1554,
   input         match_out1555,
   input         match_out1556,
   input         match_out1557,
   input         match_out1558,
   input         match_out1559,
   input         match_out1560,
   input         match_out1561,
   input         match_out1562,
   input         match_out1563,
   input         match_out1564,
   input         match_out1565,
   input         match_out1566,
   input         match_out1567,
   input         match_out1568,
   input         match_out1569,
   input         match_out1570,
   input         match_out1571,
   input         match_out1572,
   input         match_out1573,
   input         match_out1574,
   input         match_out1575,
   input         match_out1576,
   input         match_out1577,
   input         match_out1578,
   input         match_out1579,
   input         match_out1580,
   input         match_out1581,
   input         match_out1582,
   input         match_out1583,
   input         match_out1584,
   input         match_out1585,
   input         match_out1586,
   input         match_out1587,
   input         match_out1588,
   input         match_out1589,
   input         match_out1590,
   input         match_out1591,
   input         match_out1592,
   input         match_out1593,
   input         match_out1594,
   input         match_out1595,
   input         match_out1596,
   input         match_out1597,
   input         match_out1598,
   input         match_out1599,
   input         match_out1600,
   input         match_out1601,
   input         match_out1602,
   input         match_out1603,
   input         match_out1604,
   input         match_out1605,
   input         match_out1606,
   input         match_out1607,
   input         match_out1608,
   input         match_out1609,
   input         match_out1610,
   input         match_out1611,
   input         match_out1612,
   input         match_out1613,
   input         match_out1614,
   input         match_out1615,
   input         match_out1616,
   input         match_out1617,
   input         match_out1618,
   input         match_out1619,
   input         match_out1620,
   input         match_out1621,
   input         match_out1622,
   input         match_out1623,
   input         match_out1624,
   input         match_out1625,
   input         match_out1626,
   input         match_out1627,
   input         match_out1628,
   input         match_out1629,
   input         match_out1630,
   input         match_out1631,
   input         match_out1632,
   input         match_out1633,
   input         match_out1634,
   input         match_out1635,
   input         match_out1636,
   input         match_out1637,
   input         match_out1638,
   input         match_out1639,
   input         match_out1640,
   input         match_out1641,
   input         match_out1642,
   input         match_out1643,
   input         match_out1644,
   input         match_out1645,
   input         match_out1646,
   input         match_out1647,
   input         match_out1648,
   input         match_out1649,
   input         match_out1650,
   input         match_out1651,
   input         match_out1652,
   input         match_out1653,
   input         match_out1654,
   input         match_out1655,
   input         match_out1656,
   input         match_out1657,
   input         match_out1658,
   input         match_out1659,
   input         match_out1660,
   input         match_out1661,
   input         match_out1662,
   input         match_out1663,
   input         match_out1664,
   input         match_out1665,
   input         match_out1666,
   input         match_out1667,
   input         match_out1668,
   input         match_out1669,
   input         match_out1670,
   input         match_out1671,
   input         match_out1672,
   input         match_out1673,
   input         match_out1674,
   input         match_out1675,
   input         match_out1676,
   input         match_out1677,
   input         match_out1678,
   input         match_out1679,
   input         match_out1680,
   input         match_out1681,
   input         match_out1682,
   input         match_out1683,
   input         match_out1684,
   input         match_out1685,
   input         match_out1686,
   input         match_out1687,
   input         match_out1688,
   input         match_out1689,
   input         match_out1690,
   input         match_out1691,
   input         match_out1692,
   input         match_out1693,
   input         match_out1694,
   input         match_out1695,
   input         match_out1696,
   input         match_out1697,
   input         match_out1698,
   input         match_out1699,
   input         match_out1700,
   input         match_out1701,
   input         match_out1702,
   input         match_out1703,
   input         match_out1704,
   input         match_out1705,
   input         match_out1706,
   input         match_out1707,
   input         match_out1708,
   input         match_out1709,
   input         match_out1710,
   input         match_out1711,
   input         match_out1712,
   input         match_out1713,
   input         match_out1714,
   input         match_out1715,
   input         match_out1716,
   input         match_out1717,
   input         match_out1718,
   input         match_out1719,
   input         match_out1720,
   input         match_out1721,
   input         match_out1722,
   input         match_out1723,
   input         match_out1724,
   input         match_out1725,
   input         match_out1726,
   input         match_out1727,
   input         match_out1728,
   input         match_out1729,
   input         match_out1730,
   input         match_out1731,
   input         match_out1732,
   input         match_out1733,
   input         match_out1734,
   input         match_out1735,
   input         match_out1736,
   input         match_out1737,
   input         match_out1738,
   input         match_out1739,
   input         match_out1740,
   input         match_out1741,
   input         match_out1742,
   input         match_out1743,
   input         match_out1744,
   input         match_out1745,
   input         match_out1746,
   input         match_out1747,
   input         match_out1748,
   input         match_out1749,
   input         match_out1750,
   input         match_out1751,
   input         match_out1752,
   input         match_out1753,
   input         match_out1754,
   input         match_out1755,
   input         match_out1756,
   input         match_out1757,
   input         match_out1758,
   input         match_out1759,
   input         match_out1760,
   input         match_out1761,
   input         match_out1762,
   input         match_out1763,
   input         match_out1764,
   input         match_out1765,
   input         match_out1766,
   input         match_out1767,
   input         match_out1768,
   input         match_out1769,
   input         match_out1770,
   input         match_out1771,
   input         match_out1772,
   input         match_out1773,
   input         match_out1774,
   input         match_out1775,
   input         match_out1776,
   input         match_out1777,
   input         match_out1778,
   input         match_out1779,
   input         match_out1780,
   input         match_out1781,
   input         match_out1782,
   input         match_out1783,
   input         match_out1784,
   input         match_out1785,
   input         match_out1786,
   input         match_out1787,
   input         match_out1788,
   input         match_out1789,
   input         match_out1790,
   input         match_out1791,
   input         match_out1792,
   input         match_out1793,
   input         match_out1794,
   input         match_out1795,
   input         match_out1796,
   input         match_out1797,
   input         match_out1798,
   input         match_out1799,
   input         match_out1800,
   input         match_out1801,
   input         match_out1802,
   input         match_out1803,
   input         match_out1804,
   input         match_out1805,
   input         match_out1806,
   input         match_out1807,
   input         match_out1808,
   input         match_out1809,
   input         match_out1810,
   input         match_out1811,
   input         match_out1812,
   input         match_out1813,
   input         match_out1814,
   input         match_out1815,
   input         match_out1816,
   input         match_out1817,
   input         match_out1818,
   input         match_out1819,
   input         match_out1820,
   input         match_out1821,
   input         match_out1822,
   input         match_out1823,
   input         match_out1824,
   input         match_out1825,
   input         match_out1826,
   input         match_out1827,
   input         match_out1828,
   input         match_out1829,
   input         match_out1830,
   input         match_out1831,
   input         match_out1832,
   input         match_out1833,
   input         match_out1834,
   input         match_out1835,
   input         match_out1836,
   input         match_out1837,
   input         match_out1838,
   input         match_out1839,
   input         match_out1840,
   input         match_out1841,
   input         match_out1842,
   input         match_out1843,
   input         match_out1844,
   input         match_out1845,
   input         match_out1846,
   input         match_out1847,
   input         match_out1848,
   input         match_out1849,
   input         match_out1850,
   input         match_out1851,
   input         match_out1852,
   input         match_out1853,
   input         match_out1854,
   input         match_out1855,
   input         match_out1856,
   input         match_out1857,
   input         match_out1858,
   input         match_out1859,
   input         match_out1860,
   input         match_out1861,
   input         match_out1862,
   input         match_out1863,
   input         match_out1864,
   input         match_out1865,
   input         match_out1866,
   input         match_out1867,
   input         match_out1868,
   input         match_out1869,
   input         match_out1870,
   input         match_out1871,
   input         match_out1872,
   input         match_out1873,
   input         match_out1874,
   input         match_out1875,
   input         match_out1876,
   input         match_out1877,
   input         match_out1878,
   input         match_out1879,
   input         match_out1880,
   input         match_out1881,
   input         match_out1882,
   input         match_out1883,
   input         match_out1884,
   input         match_out1885,
   input         match_out1886,
   input         match_out1887,
   input         match_out1888,
   input         match_out1889,
   input         match_out1890,
   input         match_out1891,
   input         match_out1892,
   input         match_out1893,
   input         match_out1894,
   input         match_out1895,
   input         match_out1896,
   input         match_out1897,
   input         match_out1898,
   input         match_out1899,
   input         match_out1900,
   input         match_out1901,
   input         match_out1902,
   input         match_out1903,
   input         match_out1904,
   input         match_out1905,
   input         match_out1906,
   input         match_out1907,
   input         match_out1908,
   input         match_out1909,
   input         match_out1910,
   input         match_out1911,
   input         match_out1912,
   input         match_out1913,
   input         match_out1914,
   input         match_out1915,
   input         match_out1916,
   input         match_out1917,
   input         match_out1918,
   input         match_out1919,
   input         match_out1920,
   input         match_out1921,
   input         match_out1922,
   input         match_out1923,
   input         match_out1924,
   input         match_out1925,
   input         match_out1926,
   input         match_out1927,
   input         match_out1928,
   input         match_out1929,
   input         match_out1930,
   input         match_out1931,
   input         match_out1932,
   input         match_out1933,
   input         match_out1934,
   input         match_out1935,
   input         match_out1936,
   input         match_out1937,
   input         match_out1938,
   input         match_out1939,
   input         match_out1940,
   input         match_out1941,
   input         match_out1942,
   input         match_out1943,
   input         match_out1944,
   input         match_out1945,
   input         match_out1946,
   input         match_out1947,
   input         match_out1948,
   input         match_out1949,
   input         match_out1950,
   input         match_out1951,
   input         match_out1952,
   input         match_out1953,
   input         match_out1954,
   input         match_out1955,
   input         match_out1956,
   input         match_out1957,
   input         match_out1958,
   input         match_out1959,
   input         match_out1960,
   input         match_out1961,
   input         match_out1962,
   input         match_out1963,
   input         match_out1964,
   input         match_out1965,
   input         match_out1966,
   input         match_out1967,
   input         match_out1968,
   input         match_out1969,
   input         match_out1970,
   input         match_out1971,
   input         match_out1972,
   input         match_out1973,
   input         match_out1974,
   input         match_out1975,
   input         match_out1976,
   input         match_out1977,
   input         match_out1978,
   input         match_out1979,
   input         match_out1980,
   input         match_out1981,
   input         match_out1982,
   input         match_out1983,
   input         match_out1984,
   input         match_out1985,
   input         match_out1986,
   input         match_out1987,
   input         match_out1988,
   input         match_out1989,
   input         match_out1990,
   input         match_out1991,
   input         match_out1992,
   input         match_out1993,
   input         match_out1994,
   input         match_out1995,
   input         match_out1996,
   input         match_out1997,
   input         match_out1998,
   input         match_out1999,
   input         match_out2000,
   input         match_out2001,
   input         match_out2002,
   input         match_out2003,
   input         match_out2004,
   input         match_out2005,
   input         match_out2006,
   input         match_out2007,
   input         match_out2008,
   input         match_out2009,
   input         match_out2010,
   input         match_out2011,
   input         match_out2012,
   input         match_out2013,
   input         match_out2014,
   input         match_out2015,
   input         match_out2016,
   input         match_out2017,
   input         match_out2018,
   input         match_out2019,
   input         match_out2020,
   input         match_out2021,
   input         match_out2022,
   input         match_out2023,
   input         match_out2024,
   input         match_out2025,
   input         match_out2026,
   input         match_out2027,
   input         match_out2028,
   input         match_out2029,
   input         match_out2030,
   input         match_out2031,
   input         match_out2032,
   input         match_out2033,
   input         match_out2034,
   input         match_out2035,
   input         match_out2036,
   input         match_out2037,
   input         match_out2038,
   input         match_out2039,
   input         match_out2040,
   input         match_out2041,
   input         match_out2042,
   input         match_out2043,
   input         match_out2044,
   input         match_out2045,
   input         match_out2046,
   input         match_out2047,
   input         match_out2048,
   input         match_out2049,
   input         match_out2050,
   input         match_out2051,
   input         match_out2052,
   input         match_out2053,
   input         match_out2054,
   input         match_out2055,
   input         match_out2056,
   input         match_out2057,
   input         match_out2058,
   input         match_out2059,
   input         match_out2060,
   input         match_out2061,
   input         match_out2062,
   input         match_out2063,
   input         match_out2064,
   input         match_out2065,
   input         match_out2066,
   input         match_out2067,
   input         match_out2068,
   input         match_out2069,
   input         match_out2070,
   input         match_out2071,
   input         match_out2072,
   input         match_out2073,
   input         match_out2074,
   input         match_out2075,
   input         match_out2076,
   input         match_out2077,
   input         match_out2078,
   input         match_out2079,
   input         match_out2080,
   input         match_out2081,
   input         match_out2082,
   input         match_out2083,
   input         match_out2084,
   input         match_out2085,
   input         match_out2086,
   input         match_out2087,
   input         match_out2088,
   input         match_out2089,
   input         match_out2090,
   input         match_out2091,
   input         match_out2092,
   input         match_out2093,
   input         match_out2094,
   input         match_out2095,
   input         match_out2096,
   input         match_out2097,
   input         match_out2098,
   input         match_out2099,
   input         match_out2100,
   input         match_out2101,
   input         match_out2102,
   input         match_out2103,
   input         match_out2104,
   input         match_out2105,
   input         match_out2106,
   input         match_out2107,
   input         match_out2108,
   input         match_out2109,
   input         match_out2110,
   input         match_out2111,
   input         match_out2112,
   input         match_out2113,
   input         match_out2114,
   input         match_out2115,
   input         match_out2116,
   input         match_out2117,
   input         match_out2118,
   input         match_out2119,
   input         match_out2120,
   input         match_out2121,
   input         match_out2122,
   input         match_out2123,
   input         match_out2124,
   input         match_out2125,
   input         match_out2126,
   input         match_out2127,
   input         match_out2128,
   input         match_out2129,
   input         match_out2130,
   input         match_out2131,
   input         match_out2132,
   input         match_out2133,
   input         match_out2134,
   input         match_out2135,
   input         match_out2136,
   input         match_out2137,
   input         match_out2138,
   input         match_out2139,
   input         match_out2140,
   input         match_out2141,
   input         match_out2142,
   input         match_out2143,
   input         match_out2144,
   input         match_out2145,
   input         match_out2146,
   input         match_out2147,
   input         match_out2148,
   input         match_out2149,
   input         match_out2150,
   input         match_out2151,
   input         match_out2152,
   input         match_out2153,
   input         match_out2154,
   input         match_out2155,
   input         match_out2156,
   input         match_out2157,
   input         match_out2158,
   input         match_out2159,
   input         match_out2160,
   input         match_out2161,
   input         match_out2162,
   input         match_out2163,
   input         match_out2164,
   input         match_out2165,
   input         match_out2166,
   input         match_out2167,
   input         match_out2168,
   input         match_out2169,
   input         match_out2170,
   input         match_out2171,
   input         match_out2172,
   input         match_out2173,
   input         match_out2174,
   input         match_out2175,
   input         match_out2176,
   input         match_out2177,
   input         match_out2178,
   input         match_out2179,
   input         match_out2180,
   input         match_out2181,
   input         match_out2182,
   input         match_out2183,
   input         match_out2184,
   input         match_out2185,
   input         match_out2186,
   input         match_out2187,
   input         match_out2188,
   input         match_out2189,
   input         match_out2190,
   input         match_out2191,
   input         match_out2192,
   input         match_out2193,
   input         match_out2194,
   input         match_out2195,
   input         match_out2196,
   input         match_out2197,
   input         match_out2198,
   input         match_out2199,
   input         match_out2200,
   input         match_out2201,
   input         match_out2202,
   input         match_out2203,
   input         match_out2204,
   input         match_out2205,
   input         match_out2206,
   input         match_out2207,
   input         match_out2208,
   input         match_out2209,
   input         match_out2210,
   input         match_out2211,
   input         match_out2212,
   input         match_out2213,
   input         match_out2214,
   input         match_out2215,
   input         match_out2216,
   input         match_out2217,
   input         match_out2218,
   input         match_out2219,
   input         match_out2220,
   input         match_out2221,
   input         match_out2222,
   input         match_out2223,
   input         match_out2224,
   input         match_out2225,
   input         match_out2226,
   input         match_out2227,
   input         match_out2228,
   input         match_out2229,
   input         match_out2230,
   input         match_out2231,
   input         match_out2232,
   input         match_out2233,
   input         match_out2234,
   input         match_out2235,
   input         match_out2236,
   input         match_out2237,
   input         match_out2238,
   input         match_out2239,
   input         match_out2240,
   input         match_out2241,
   input         match_out2242,
   input         match_out2243,
   input         match_out2244,
   input         match_out2245,
   input         match_out2246,
   input         match_out2247,
   input         match_out2248,
   input         match_out2249,
   input         match_out2250,
   input         match_out2251,
   input         match_out2252,
   input         match_out2253,
   input         match_out2254,
   input         match_out2255,
   input         match_out2256,
   input         match_out2257,
   input         match_out2258,
   input         match_out2259,
   input         match_out2260,
   input         match_out2261,
   input         match_out2262,
   input         match_out2263,
   input         match_out2264,
   input         match_out2265,
   input         match_out2266,
   input         match_out2267,
   input         match_out2268,
   input         match_out2269,
   input         match_out2270,
   input         match_out2271,
   input         match_out2272,
   input         match_out2273,
   input         match_out2274,
   input         match_out2275,
   input         match_out2276,
   input         match_out2277,
   input         match_out2278,
   input         match_out2279,
   input         match_out2280,
   input         match_out2281,
   input         match_out2282,
   input         match_out2283,
   input         match_out2284,
   input         match_out2285,
   input         match_out2286,
   input         match_out2287,
   input         match_out2288,
   input         match_out2289,
   input         match_out2290,
   input         match_out2291,
   input         match_out2292,
   input         match_out2293,
   input         match_out2294,
   input         match_out2295,
   input         match_out2296,
   input         match_out2297,
   input         match_out2298,
   input         match_out2299,
   input         match_out2300,
   input         match_out2301,
   input         match_out2302,
   input         match_out2303,
   input         match_out2304,
   input         match_out2305,
   input         match_out2306,
   input         match_out2307,
   input         match_out2308,
   input         match_out2309,
   input         match_out2310,
   input         match_out2311,
   input         match_out2312,
   input         match_out2313,
   input         match_out2314,
   input         match_out2315,
   input         match_out2316,
   input         match_out2317,
   input         match_out2318,
   input         match_out2319,
   input         match_out2320,
   input         match_out2321,
   input         match_out2322,
   input         match_out2323,
   input         match_out2324,
   input         match_out2325,
   input         match_out2326,
   input         match_out2327,
   input         match_out2328,
   input         match_out2329,
   input         match_out2330,
   input         match_out2331,
   input         match_out2332,
   input         match_out2333,
   input         match_out2334,
   input         match_out2335,
   input         match_out2336,
   input         match_out2337,
   input         match_out2338,
   input         match_out2339,
   input         match_out2340,
   input         match_out2341,
   input         match_out2342,
   input         match_out2343,
   input         match_out2344,
   input         match_out2345,
   input         match_out2346,
   input         match_out2347,
   input         match_out2348,
   input         match_out2349,
   input         match_out2350,
   input         match_out2351,
   input         match_out2352,
   input         match_out2353,
   input         match_out2354,
   input         match_out2355,
   input         match_out2356,
   input         match_out2357,
   input         match_out2358,
   input         match_out2359,
   input         match_out2360,
   input         match_out2361,
   input         match_out2362,
   input         match_out2363,
   input         match_out2364,
   input         match_out2365,
   input         match_out2366,
   input         match_out2367,
   input         match_out2368,
   input         match_out2369,
   input         match_out2370,
   input         match_out2371,
   input         match_out2372,
   input         match_out2373,
   input         match_out2374,
   input         match_out2375,
   input         match_out2376,
   input         match_out2377,
   input         match_out2378,
   input         match_out2379,
   input         match_out2380,
   input         match_out2381,
   input         match_out2382,
   input         match_out2383,
   input         match_out2384,
   input         match_out2385,
   input         match_out2386,
   input         match_out2387,
   input         match_out2388,
   input         match_out2389,
   input         match_out2390,
   input         match_out2391,
   input         match_out2392,
   input         match_out2393,
   input         match_out2394,
   input         match_out2395,
   input         match_out2396,
   input         match_out2397,
   input         match_out2398,
   input         match_out2399,
   input         match_out2400,
   input         match_out2401,
   input         match_out2402,
   input         match_out2403,
   input         match_out2404,
   input         match_out2405,
   input         match_out2406,
   input         match_out2407,
   input         match_out2408,
   input         match_out2409,
   input         match_out2410,
   input         match_out2411,
   input         match_out2412,
   input         match_out2413,
   input         match_out2414,
   input         match_out2415,
   input         match_out2416,
   input         match_out2417,
   input         match_out2418,
   input         match_out2419,
   input         match_out2420,
   input         match_out2421,
   input         match_out2422,
   input         match_out2423,
   input         match_out2424,
   input         match_out2425,
   input         match_out2426,
   input         match_out2427,
   input         match_out2428,
   input         match_out2429,
   input         match_out2430,
   input         match_out2431,
   input         match_out2432,
   input         match_out2433,
   input         match_out2434,
   input         match_out2435,
   input         match_out2436,
   input         match_out2437,
   input         match_out2438,
   input         match_out2439,
   input         match_out2440,
   input         match_out2441,
   input         match_out2442,
   input         match_out2443,
   input         match_out2444,
   input         match_out2445,
   input         match_out2446,
   input         match_out2447,
   input         match_out2448,
   input         match_out2449,
   input         match_out2450,
   input         match_out2451,
   input         match_out2452,
   input         match_out2453,
   input         match_out2454,
   input         match_out2455,
   input         match_out2456,
   input         match_out2457,
   input         match_out2458,
   input         match_out2459,
   input         match_out2460,
   input         match_out2461,
   input         match_out2462,
   input         match_out2463,
   input         match_out2464,
   input         match_out2465,
   input         match_out2466,
   input         match_out2467,
   input         match_out2468,
   input         match_out2469,
   input         match_out2470,
   input         match_out2471,
   input         match_out2472,
   input         match_out2473,
   input         match_out2474,
   input         match_out2475,
   input         match_out2476,
   input         match_out2477,
   input         match_out2478,
   input         match_out2479,
   input         match_out2480,
   input         match_out2481,
   input         match_out2482,
   input         match_out2483,
   input         match_out2484,
   input         match_out2485,
   input         match_out2486,
   input         match_out2487,
   input         match_out2488,
   input         match_out2489,
   input         match_out2490,
   input         match_out2491,
   input         match_out2492,
   input         match_out2493,
   input         match_out2494,
   input         match_out2495,
   input         match_out2496,
   input         match_out2497,
   input         match_out2498,
   input         match_out2499,
   input         match_out2500,
   input         match_out2501,
   input         match_out2502,
   input         match_out2503,
   input         match_out2504,
   input         match_out2505,
   input         match_out2506,
   input         match_out2507,
   input         match_out2508,
   input         match_out2509,
   input         match_out2510,
   input         match_out2511,
   input         match_out2512,
   input         match_out2513,
   input         match_out2514,
   input         match_out2515,
   input         match_out2516,
   input         match_out2517,
   input         match_out2518,
   input         match_out2519,
   input         match_out2520,
   input         match_out2521,
   input         match_out2522,
   input         match_out2523,
   input         match_out2524,
   input         match_out2525,
   input         match_out2526,
   input         match_out2527,
   input         match_out2528,
   input         match_out2529,
   input         match_out2530,
   input         match_out2531,
   input         match_out2532,
   input         match_out2533,
   input         match_out2534,
   input         match_out2535,
   input         match_out2536,
   input         match_out2537,
   input         match_out2538,
   input         match_out2539,
   input         match_out2540,
   input         match_out2541,
   input         match_out2542,
   input         match_out2543,
   input         match_out2544,
   input         match_out2545,
   input         match_out2546,
   input         match_out2547,
   input         match_out2548,
   input         match_out2549,
   input         match_out2550,
   input         match_out2551,
   input         match_out2552,
   input         match_out2553,
   input         match_out2554,
   input         match_out2555,
   input         match_out2556,
   input         match_out2557,
   input         match_out2558,
   input         match_out2559,
   input         match_out2560,
   input         match_out2561,
   input         match_out2562,
   input         match_out2563,
   input         match_out2564,
   input         match_out2565,
   input         match_out2566,
   input         match_out2567,
   input         match_out2568,
   input         match_out2569,
   input         match_out2570,
   input         match_out2571,
   input         match_out2572,
   input         match_out2573,
   input         match_out2574,
   input         match_out2575,
   input         match_out2576,
   input         match_out2577,
   input         match_out2578,
   input         match_out2579,
   input         match_out2580,
   input         match_out2581,
   input         match_out2582,
   input         match_out2583,
   input         match_out2584,
   input         match_out2585,
   input         match_out2586,
   input         match_out2587,
   input         match_out2588,
   input         match_out2589,
   input         match_out2590,
   input         match_out2591,
   input         match_out2592,
   input         match_out2593,
   input         match_out2594,
   input         match_out2595,
   input         match_out2596,
   input         match_out2597,
   input         match_out2598,
   input         match_out2599,
   input         match_out2600,
   input         match_out2601,
   input         match_out2602,
   input         match_out2603,
   input         match_out2604,
   input         match_out2605,
   input         match_out2606,
   input         match_out2607,
   input         match_out2608,
   input         match_out2609,
   input         match_out2610,
   input         match_out2611,
   input         match_out2612,
   input         match_out2613,
   input         match_out2614,
   input         match_out2615,
   input         match_out2616,
   input         match_out2617,
   input         match_out2618,
   input         match_out2619,
   input         match_out2620,
   input         match_out2621,
   input         match_out2622,
   input         match_out2623,
   input         match_out2624,
   input         match_out2625,
   input         match_out2626,
   input         match_out2627,
   input         match_out2628,
   input         match_out2629,
   input         match_out2630,
   input         match_out2631,
   input         match_out2632,
   input         match_out2633,
   input         match_out2634,
   input         match_out2635,
   input         match_out2636,
   input         match_out2637,
   input         match_out2638,
   input         match_out2639,
   input         match_out2640,
   input         match_out2641,
   input         match_out2642,
   input         match_out2643,
   input         match_out2644,
   input         match_out2645,
   input         match_out2646,
   input         match_out2647,
   input         match_out2648,
   input         match_out2649,
   input         match_out2650,
   input         match_out2651,
   input         match_out2652,
   input         match_out2653,
   input         match_out2654,
   input         match_out2655,
   input         match_out2656,
   input         match_out2657,
   input         match_out2658,
   input         match_out2659,
   input         match_out2660,
   input         match_out2661,
   input         match_out2662,
   input         match_out2663,
   input         match_out2664,
   input         match_out2665,
   input         match_out2666,
   input         match_out2667,
   input         match_out2668,
   input         match_out2669,
   input         match_out2670,
   input         match_out2671,
   input         match_out2672,
   input         match_out2673,
   input         match_out2674,
   input         match_out2675,
   input         match_out2676,
   input         match_out2677,
   input         match_out2678,
   input         match_out2679,
   input         match_out2680,
   input         match_out2681,
   input         match_out2682,
   input         match_out2683,
   input         match_out2684,
   input         match_out2685,
   input         match_out2686,
   input         match_out2687,
   input         match_out2688,
   input         match_out2689,
   input         match_out2690,
   input         match_out2691,
   input         match_out2692,
   input         match_out2693,
   input         match_out2694,
   input         match_out2695,
   input         match_out2696,
   input         match_out2697,
   input         match_out2698,
   input         match_out2699,
   input         match_out2700,
   input         match_out2701,
   input         match_out2702,
   input         match_out2703,
   input         match_out2704,
   input         match_out2705,
   input         match_out2706,
   input         match_out2707,
   input         match_out2708,
   input         match_out2709,
   input         match_out2710,
   input         match_out2711,
   input         match_out2712,
   input         match_out2713,
   input         match_out2714,
   input         match_out2715,
   input         match_out2716,
   input         match_out2717,
   input         match_out2718,
   input         match_out2719,
   input         match_out2720,
   input         match_out2721,
   input         match_out2722,
   input         match_out2723,
   input         match_out2724,
   input         match_out2725,
   input         match_out2726,
   input         match_out2727,
   input         match_out2728,
   input         match_out2729,
   input         match_out2730,
   input         match_out2731,
   input         match_out2732,
   input         match_out2733,
   input         match_out2734,
   input         match_out2735,
   input         match_out2736,
   input         match_out2737,
   input         match_out2738,
   input         match_out2739,
   input         match_out2740,
   input         match_out2741,
   input         match_out2742,
   input         match_out2743,
   input         match_out2744,
   input         match_out2745,
   input         match_out2746,
   input         match_out2747,
   input         match_out2748,
   input         match_out2749,
   input         match_out2750,
   input         match_out2751,
   input         match_out2752,
   input         match_out2753,
   input         match_out2754,
   input         match_out2755,
   input         match_out2756,
   input         match_out2757,
   input         match_out2758,
   input         match_out2759,
   input         match_out2760,
   input         match_out2761,
   input         match_out2762,
   input         match_out2763,
   input         match_out2764,
   input         match_out2765,
   input         match_out2766,
   input         match_out2767,
   input         match_out2768,
   input         match_out2769,
   input         match_out2770,
   input         match_out2771,
   input         match_out2772,
   input         match_out2773,
   input         match_out2774,
   input         match_out2775,
   input         match_out2776,
   input         match_out2777,
   input         match_out2778,
   input         match_out2779,
   input         match_out2780,
   input         match_out2781,
   input         match_out2782,
   input         match_out2783,
   input         match_out2784,
   input         match_out2785,
   input         match_out2786,
   input         match_out2787,
   input         match_out2788,
   input         match_out2789,
   input         match_out2790,
   input         match_out2791,
   input         match_out2792,
   input         match_out2793,
   input         match_out2794,
   input         match_out2795,
   input         match_out2796,
   input         match_out2797,
   input         match_out2798,
   input         match_out2799,
   input         match_out2800,
   input         match_out2801,
   input         match_out2802,
   input         match_out2803,
   input         match_out2804,
   input         match_out2805,
   input         match_out2806,
   input         match_out2807,
   input         match_out2808,
   input         match_out2809,
   input         match_out2810,
   input         match_out2811,
   input         match_out2812,
   input         match_out2813,
   input         match_out2814,
   input         match_out2815,
   input         match_out2816,
   input         match_out2817,
   input         match_out2818,
   input         match_out2819,
   input         match_out2820,
   input         match_out2821,
   input         match_out2822,
   input         match_out2823,
   input         match_out2824,
   input         match_out2825,
   input         match_out2826,
   input         match_out2827,
   input         match_out2828,
   input         match_out2829,
   input         match_out2830,
   input         match_out2831,
   input         match_out2832,
   input         match_out2833,
   input         match_out2834,
   input         match_out2835,
   input         match_out2836,
   input         match_out2837,
   input         match_out2838,
   input         match_out2839,
   input         match_out2840,
   input         match_out2841,
   input         match_out2842,
   input         match_out2843,
   input         match_out2844,
   input         match_out2845,
   input         match_out2846,
   input         match_out2847,
   input         match_out2848,
   input         match_out2849,
   input         match_out2850,
   input         match_out2851,
   input         match_out2852,
   input         match_out2853,
   input         match_out2854,
   input         match_out2855,
   input         match_out2856,
   input         match_out2857,
   input         match_out2858,
   input         match_out2859,
   input         match_out2860,
   input         match_out2861,
   input         match_out2862,
   input         match_out2863,
   input         match_out2864,
   input         match_out2865,
   input         match_out2866,
   input         match_out2867,
   input         match_out2868,
   input         match_out2869,
   input         match_out2870,
   input         match_out2871,
   input         match_out2872,
   input         match_out2873,
   input         match_out2874,
   input         match_out2875,
   input         match_out2876,
   input         match_out2877,
   input         match_out2878,
   input         match_out2879,
   input         match_out2880,
   input         match_out2881,
   input         match_out2882,
   input         match_out2883,
   input         match_out2884,
   input         match_out2885,
   input         match_out2886,
   input         match_out2887,
   input         match_out2888,
   input         match_out2889,
   input         match_out2890,
   input         match_out2891,
   input         match_out2892,
   input         match_out2893,
   input         match_out2894,
   input         match_out2895,
   input         match_out2896,
   input         match_out2897,
   input         match_out2898,
   input         match_out2899,
   input         match_out2900,
   input         match_out2901,
   input         match_out2902,
   input         match_out2903,
   input         match_out2904,
   input         match_out2905,
   input         match_out2906,
   input         match_out2907,
   input         match_out2908,
   input         match_out2909,
   input         match_out2910,
   input         match_out2911,
   input         match_out2912,
   input         match_out2913,
   input         match_out2914,
   input         match_out2915,
   input         match_out2916,
   input         match_out2917,
   input         match_out2918,
   input         match_out2919,
   input         match_out2920,
   input         match_out2921,
   input         match_out2922,
   input         match_out2923,
   input         match_out2924,
   input         match_out2925,
   input         match_out2926,
   input         match_out2927,
   input         match_out2928,
   input         match_out2929,
   input         match_out2930,
   input         match_out2931,
   input         match_out2932,
   input         match_out2933,
   input         match_out2934,
   input         match_out2935,
   input         match_out2936,
   input         match_out2937,
   input         match_out2938,
   input         match_out2939,
   input         match_out2940,
   input         match_out2941,
   input         match_out2942,
   input         match_out2943,
   input         match_out2944,
   input         match_out2945,
   input         match_out2946,
   input         match_out2947,
   input         match_out2948,
   input         match_out2949,
   input         match_out2950,
   input         match_out2951,
   input         match_out2952,
   input         match_out2953,
   input         match_out2954,
   input         match_out2955,
   input         match_out2956,
   input         match_out2957,
   input         match_out2958,
   input         match_out2959,
   input         match_out2960,
   input         match_out2961,
   input         match_out2962,
   input         match_out2963,
   input         match_out2964,
   input         match_out2965,
   input         match_out2966,
   input         match_out2967,
   input         match_out2968,
   input         match_out2969,
   input         match_out2970,
   input         match_out2971,
   input         match_out2972,
   input         match_out2973,
   input         match_out2974,
   input         match_out2975,
   input         match_out2976,
   input         match_out2977,
   input         match_out2978,
   input         match_out2979,
   input         match_out2980,
   input         match_out2981,
   input         match_out2982,
   input         match_out2983,
   input         match_out2984,
   input         match_out2985,
   input         match_out2986,
   input         match_out2987,
   input         match_out2988,
   input         match_out2989,
   input         match_out2990,
   input         match_out2991,
   input         match_out2992,
   input         match_out2993,
   input         match_out2994,
   input         match_out2995,
   input         match_out2996,
   input         match_out2997,
   input         match_out2998,
   input         match_out2999,
   input         match_out3000,
   input         match_out3001,
   input         match_out3002,
   input         match_out3003,
   input         match_out3004,
   input         match_out3005,
   input         match_out3006,
   input         match_out3007,
   input         match_out3008,
   input         match_out3009,
   input         match_out3010,
   input         match_out3011,
   input         match_out3012,
   input         match_out3013,
   input         match_out3014,
   input         match_out3015,
   input         match_out3016,
   input         match_out3017,
   input         match_out3018,
   input         match_out3019,
   input         match_out3020,
   input         match_out3021,
   input         match_out3022,
   input         match_out3023,
   input         match_out3024,
   input         match_out3025,
   input         match_out3026,
   input         match_out3027,
   input         match_out3028,
   input         match_out3029,
   input         match_out3030,
   input         match_out3031,
   input         match_out3032,
   input         match_out3033,
   input         match_out3034,
   input         match_out3035,
   input         match_out3036,
   input         match_out3037,
   input         match_out3038,
   input         match_out3039,
   input         match_out3040,
   input         match_out3041,
   input         match_out3042,
   input         match_out3043,
   input         match_out3044,
   input         match_out3045,
   input         match_out3046,
   input         match_out3047,
   input         match_out3048,
   input         match_out3049,
   input         match_out3050,
   input         match_out3051,
   input         match_out3052,
   input         match_out3053,
   input         match_out3054,
   input         match_out3055,
   input         match_out3056,
   input         match_out3057,
   input         match_out3058,
   input         match_out3059,
   input         match_out3060,
   input         match_out3061,
   input         match_out3062,
   input         match_out3063,
   input         match_out3064,
   input         match_out3065,
   input         match_out3066,
   input         match_out3067,
   input         match_out3068,
   input         match_out3069,
   input         match_out3070,
   input         match_out3071,
   input         match_out3072,
   input         match_out3073,
   input         match_out3074,
   input         match_out3075,
   input         match_out3076,
   input         match_out3077,
   input         match_out3078,
   input         match_out3079,
   input         match_out3080,
   input         match_out3081,
   input         match_out3082,
   input         match_out3083,
   input         match_out3084,
   input         match_out3085,
   input         match_out3086,
   input         match_out3087,
   input         match_out3088,
   input         match_out3089,
   input         match_out3090,
   input         match_out3091,
   input         match_out3092,
   input         match_out3093,
   input         match_out3094,
   input         match_out3095,
   input         match_out3096,
   input         match_out3097,
   input         match_out3098,
   input         match_out3099,
   input         match_out3100,
   input         match_out3101,
   input         match_out3102,
   input         match_out3103,
   input         match_out3104,
   input         match_out3105,
   input         match_out3106,
   input         match_out3107,
   input         match_out3108,
   input         match_out3109,
   input         match_out3110,
   input         match_out3111,
   input         match_out3112,
   input         match_out3113,
   input         match_out3114,
   input         match_out3115,
   input         match_out3116,
   input         match_out3117,
   input         match_out3118,
   input         match_out3119,
   input         match_out3120,
   input         match_out3121,
   input         match_out3122,
   input         match_out3123,
   input         match_out3124,
   input         match_out3125,
   input         match_out3126,
   input         match_out3127,
   input         match_out3128,
   input         match_out3129,
   input         match_out3130,
   input         match_out3131,
   input         match_out3132,
   input         match_out3133,
   input         match_out3134,
   input         match_out3135,
   input         match_out3136,
   input         match_out3137,
   input         match_out3138,
   input         match_out3139,
   input         match_out3140,
   input         match_out3141,
   input         match_out3142,
   input         match_out3143,
   input         match_out3144,
   input         match_out3145,
   input         match_out3146,
   input         match_out3147,
   input         match_out3148,
   input         match_out3149,
   input         match_out3150,
   input         match_out3151,
   input         match_out3152,
   input         match_out3153,
   input         match_out3154,
   input         match_out3155,
   input         match_out3156,
   input         match_out3157,
   input         match_out3158,
   input         match_out3159,
   input         match_out3160,
   input         match_out3161,
   input         match_out3162,
   input         match_out3163,
   input         match_out3164,
   input         match_out3165,
   input         match_out3166,
   input         match_out3167,
   input         match_out3168,
   input         match_out3169,
   input         match_out3170,
   input         match_out3171,
   input         match_out3172,
   input         match_out3173,
   input         match_out3174,
   input         match_out3175,
   input         match_out3176,
   input         match_out3177,
   input         match_out3178,
   input         match_out3179,
   input         match_out3180,
   input         match_out3181,
   input         match_out3182,
   input         match_out3183,
   input         match_out3184,
   input         match_out3185,
   input         match_out3186,
   input         match_out3187,
   input         match_out3188,
   input         match_out3189,
   input         match_out3190,
   input         match_out3191,
   input         match_out3192,
   input         match_out3193,
   input         match_out3194,
   input         match_out3195,
   input         match_out3196,
   input         match_out3197,
   input         match_out3198,
   input         match_out3199,
   input         match_out3200,
   input         match_out3201,
   input         match_out3202,
   input         match_out3203,
   input         match_out3204,
   input         match_out3205,
   input         match_out3206,
   input         match_out3207,
   input         match_out3208,
   input         match_out3209,
   input         match_out3210,
   input         match_out3211,
   input         match_out3212,
   input         match_out3213,
   input         match_out3214,
   input         match_out3215,
   input         match_out3216,
   input         match_out3217,
   input         match_out3218,
   input         match_out3219,
   input         match_out3220,
   input         match_out3221,
   input         match_out3222,
   input         match_out3223,
   input         match_out3224,
   input         match_out3225,
   input         match_out3226,
   input         match_out3227,
   input         match_out3228,
   input         match_out3229,
   input         match_out3230,
   input         match_out3231,
   input         match_out3232,
   input         match_out3233,
   input         match_out3234,
   input         match_out3235,
   input         match_out3236,
   input         match_out3237,
   input         match_out3238,
   input         match_out3239,
   input         match_out3240,
   input         match_out3241,
   input         match_out3242,
   input         match_out3243,
   input         match_out3244,
   input         match_out3245,
   input         match_out3246,
   input         match_out3247,
   input         match_out3248,
   input         match_out3249,
   input         match_out3250,
   input         match_out3251,
   input         match_out3252,
   input         match_out3253,
   input         match_out3254,
   input         match_out3255,
   input         match_out3256,
   input         match_out3257,
   input         match_out3258,
   input         match_out3259,
   input         match_out3260,
   input         match_out3261,
   input         match_out3262,
   input         match_out3263,
   input         match_out3264,
   input         match_out3265,
   input         match_out3266,
   input         match_out3267,
   input         match_out3268,
   input         match_out3269,
   input         match_out3270,
   input         match_out3271,
   input         match_out3272,
   input         match_out3273,
   input         match_out3274,
   input         match_out3275,
   input         match_out3276,
   input         match_out3277,
   input         match_out3278,
   input         match_out3279,
   input         match_out3280,
   input         match_out3281,
   input         match_out3282,
   input         match_out3283,
   input         match_out3284,
   input         match_out3285,
   input         match_out3286,
   input         match_out3287,
   input         match_out3288,
   input         match_out3289,
   input         match_out3290,
   input         match_out3291,
   input         match_out3292,
   input         match_out3293,
   input         match_out3294,
   input         match_out3295,
   input         match_out3296,
   input         match_out3297,
   input         match_out3298,
   input         match_out3299,
   input         match_out3300,
   input         match_out3301,
   input         match_out3302,
   input         match_out3303,
   input         match_out3304,
   input         match_out3305,
   input         match_out3306,
   input         match_out3307,
   input         match_out3308,
   input         match_out3309,
   input         match_out3310,
   input         match_out3311,
   input         match_out3312,
   input         match_out3313,
   input         match_out3314,
   input         match_out3315,
   input         match_out3316,
   input         match_out3317,
   input         match_out3318,
   input         match_out3319,
   input         match_out3320,
   input         match_out3321,
   input         match_out3322,
   input         match_out3323,
   input         match_out3324,
   input         match_out3325,
   input         match_out3326,
   input         match_out3327,
   input         match_out3328,
   input         match_out3329,
   input         match_out3330,
   input         match_out3331,
   input         match_out3332,
   input         match_out3333,
   input         match_out3334,
   input         match_out3335,
   input         match_out3336,
   input         match_out3337,
   input         match_out3338,
   input         match_out3339,
   input         match_out3340,
   input         match_out3341,
   input         match_out3342,
   input         match_out3343,
   input         match_out3344,
   input         match_out3345,
   input         match_out3346,
   input         match_out3347,
   input         match_out3348,
   input         match_out3349,
   input         match_out3350,
   input         match_out3351,
   input         match_out3352,
   input         match_out3353,
   input         match_out3354,
   input         match_out3355,
   input         match_out3356,
   input         match_out3357,
   input         match_out3358,
   input         match_out3359,
   input         match_out3360,
   input         match_out3361,
   input         match_out3362,
   input         match_out3363,
   input         match_out3364,
   input         match_out3365,
   input         match_out3366,
   input         match_out3367,
   input         match_out3368,
   input         match_out3369,
   input         match_out3370,
   input         match_out3371,
   input         match_out3372,
   input         match_out3373,
   input         match_out3374,
   input         match_out3375,
   input         match_out3376,
   input         match_out3377,
   input         match_out3378,
   input         match_out3379,
   input         match_out3380,
   input         match_out3381,
   input         match_out3382,
   input         match_out3383,
   input         match_out3384,
   input         match_out3385,
   input         match_out3386,
   input         match_out3387,
   input         match_out3388,
   input         match_out3389,
   input         match_out3390,
   input         match_out3391,
   input         match_out3392,
   input         match_out3393,
   input         match_out3394,
   input         match_out3395,
   input         match_out3396,
   input         match_out3397,
   input         match_out3398,
   input         match_out3399,
   input         match_out3400,
   input         match_out3401,
   input         match_out3402,
   input         match_out3403,
   input         match_out3404,
   input         match_out3405,
   input         match_out3406,
   input         match_out3407,
   input         match_out3408,
   input         match_out3409,
   input         match_out3410,
   input         match_out3411,
   input         match_out3412,
   input         match_out3413,
   input         match_out3414,
   input         match_out3415,
   input         match_out3416,
   input         match_out3417,
   input         match_out3418,
   input         match_out3419,
   input         match_out3420,
   input         match_out3421,
   input         match_out3422,
   input         match_out3423,
   input         match_out3424,
   input         match_out3425,
   input         match_out3426,
   input         match_out3427,
   input         match_out3428,
   input         match_out3429,
   input         match_out3430,
   input         match_out3431,
   input         match_out3432,
   input         match_out3433,
   input         match_out3434,
   input         match_out3435,
   input         match_out3436,
   input         match_out3437,
   input         match_out3438,
   input         match_out3439,
   input         match_out3440,
   input         match_out3441,
   input         match_out3442,
   input         match_out3443,
   input         match_out3444,
   input         match_out3445,
   input         match_out3446,
   input         match_out3447,
   input         match_out3448,
   input         match_out3449,
   input         match_out3450,
   input         match_out3451,
   input         match_out3452,
   input         match_out3453,
   input         match_out3454,
   input         match_out3455,
   input         match_out3456,
   input         match_out3457,
   input         match_out3458,
   input         match_out3459,
   input         match_out3460,
   input         match_out3461,
   input         match_out3462,
   input         match_out3463,
   input         match_out3464,
   input         match_out3465,
   input         match_out3466,
   input         match_out3467,
   input         match_out3468,
   input         match_out3469,
   input         match_out3470,
   input         match_out3471,
   input         match_out3472,
   input         match_out3473,
   input         match_out3474,
   input         match_out3475,
   input         match_out3476,
   input         match_out3477,
   input         match_out3478,
   input         match_out3479,
   input         match_out3480,
   input         match_out3481,
   input         match_out3482,
   input         match_out3483,
   input         match_out3484,
   input         match_out3485,
   input         match_out3486,
   input         match_out3487,
   input         match_out3488,
   input         match_out3489,
   input         match_out3490,
   input         match_out3491,
   input         match_out3492,
   input         match_out3493,
   input         match_out3494,
   input         match_out3495,
   input         match_out3496,
   input         match_out3497,
   input         match_out3498,
   input         match_out3499,
   input         match_out3500,
   input         match_out3501,
   input         match_out3502,
   input         match_out3503,
   input         match_out3504,
   input         match_out3505,
   input         match_out3506,
   input         match_out3507,
   input         match_out3508,
   input         match_out3509,
   input         match_out3510,
   input         match_out3511,
   input         match_out3512,
   input         match_out3513,
   input         match_out3514,
   input         match_out3515,
   input         match_out3516,
   input         match_out3517,
   input         match_out3518,
   input         match_out3519,
   input         match_out3520,
   input         match_out3521,
   input         match_out3522,
   input         match_out3523,
   input         match_out3524,
   input         match_out3525,
   input         match_out3526,
   input         match_out3527,
   input         match_out3528,
   input         match_out3529,
   input         match_out3530,
   input         match_out3531,
   input         match_out3532,
   input         match_out3533,
   input         match_out3534,
   input         match_out3535,
   input         match_out3536,
   input         match_out3537,
   input         match_out3538,
   input         match_out3539,
   input         match_out3540,
   input         match_out3541,
   input         match_out3542,
   input         match_out3543,
   input         match_out3544,
   input         match_out3545,
   input         match_out3546,
   input         match_out3547,
   input         match_out3548,
   input         match_out3549,
   input         match_out3550,
   input         match_out3551,
   input         match_out3552,
   input         match_out3553,
   input         match_out3554,
   input         match_out3555,
   input         match_out3556,
   input         match_out3557,
   input         match_out3558,
   input         match_out3559,
   input         match_out3560,
   input         match_out3561,
   input         match_out3562,
   input         match_out3563,
   input         match_out3564,
   input         match_out3565,
   input         match_out3566,
   input         match_out3567,
   input         match_out3568,
   input         match_out3569,
   input         match_out3570,
   input         match_out3571,
   input         match_out3572,
   input         match_out3573,
   input         match_out3574,
   input         match_out3575,
   input         match_out3576,
   input         match_out3577,
   input         match_out3578,
   input         match_out3579,
   input         match_out3580,
   input         match_out3581,
   input         match_out3582,
   input         match_out3583,
   input         match_out3584,
   input         match_out3585,
   input         match_out3586,
   input         match_out3587,
   input         match_out3588,
   input         match_out3589,
   input         match_out3590,
   input         match_out3591,
   input         match_out3592,
   input         match_out3593,
   input         match_out3594,
   input         match_out3595,
   input         match_out3596,
   input         match_out3597,
   input         match_out3598,
   input         match_out3599,
   input         match_out3600,
   input         match_out3601,
   input         match_out3602,
   input         match_out3603,
   input         match_out3604,
   input         match_out3605,
   input         match_out3606,
   input         match_out3607,
   input         match_out3608,
   input         match_out3609,
   input         match_out3610,
   input         match_out3611,
   input         match_out3612,
   input         match_out3613,
   input         match_out3614,
   input         match_out3615,
   input         match_out3616,
   input         match_out3617,
   input         match_out3618,
   input         match_out3619,
   input         match_out3620,
   input         match_out3621,
   input         match_out3622,
   input         match_out3623,
   input         match_out3624,
   input         match_out3625,
   input         match_out3626,
   input         match_out3627,
   input         match_out3628,
   input         match_out3629,
   input         match_out3630,
   input         match_out3631,
   input         match_out3632,
   input         match_out3633,
   input         match_out3634,
   input         match_out3635,
   input         match_out3636,
   input         match_out3637,
   input         match_out3638,
   input         match_out3639,
   input         match_out3640,
   input         match_out3641,
   input         match_out3642,
   input         match_out3643,
   input         match_out3644,
   input         match_out3645,
   input         match_out3646,
   input         match_out3647,
   input         match_out3648,
   input         match_out3649,
   input         match_out3650,
   input         match_out3651,
   input         match_out3652,
   input         match_out3653,
   input         match_out3654,
   input         match_out3655,
   input         match_out3656,
   input         match_out3657,
   input         match_out3658,
   input         match_out3659,
   input         match_out3660,
   input         match_out3661,
   input         match_out3662,
   input         match_out3663,
   input         match_out3664,
   input         match_out3665,
   input         match_out3666,
   input         match_out3667,
   input         match_out3668,
   input         match_out3669,
   input         match_out3670,
   input         match_out3671,
   input         match_out3672,
   input         match_out3673,
   input         match_out3674,
   input         match_out3675,
   input         match_out3676,
   input         match_out3677,
   input         match_out3678,
   input         match_out3679,
   input         match_out3680,
   input         match_out3681,
   input         match_out3682,
   input         match_out3683,
   input         match_out3684,
   input         match_out3685,
   input         match_out3686,
   input         match_out3687,
   input         match_out3688,
   input         match_out3689,
   input         match_out3690,
   input         match_out3691,
   input         match_out3692,
   input         match_out3693,
   input         match_out3694,
   input         match_out3695,
   input         match_out3696,
   input         match_out3697,
   input         match_out3698,
   input         match_out3699,
   input         match_out3700,
   input         match_out3701,
   input         match_out3702,
   input         match_out3703,
   input         match_out3704,
   input         match_out3705,
   input         match_out3706,
   input         match_out3707,
   input         match_out3708,
   input         match_out3709,
   input         match_out3710,
   input         match_out3711,
   input         match_out3712,
   input         match_out3713,
   input         match_out3714,
   input         match_out3715,
   input         match_out3716,
   input         match_out3717,
   input         match_out3718,
   input         match_out3719,
   input         match_out3720,
   input         match_out3721,
   input         match_out3722,
   input         match_out3723,
   input         match_out3724,
   input         match_out3725,
   input         match_out3726,
   input         match_out3727,
   input         match_out3728,
   input         match_out3729,
   input         match_out3730,
   input         match_out3731,
   input         match_out3732,
   input         match_out3733,
   input         match_out3734,
   input         match_out3735,
   input         match_out3736,
   input         match_out3737,
   input         match_out3738,
   input         match_out3739,
   input         match_out3740,
   input         match_out3741,
   input         match_out3742,
   input         match_out3743,
   input         match_out3744,
   input         match_out3745,
   input         match_out3746,
   input         match_out3747,
   input         match_out3748,
   input         match_out3749,
   input         match_out3750,
   input         match_out3751,
   input         match_out3752,
   input         match_out3753,
   input         match_out3754,
   input         match_out3755,
   input         match_out3756,
   input         match_out3757,
   input         match_out3758,
   input         match_out3759,
   input         match_out3760,
   input         match_out3761,
   input         match_out3762,
   input         match_out3763,
   input         match_out3764,
   input         match_out3765,
   input         match_out3766,
   input         match_out3767,
   input         match_out3768,
   input         match_out3769,
   input         match_out3770,
   input         match_out3771,
   input         match_out3772,
   input         match_out3773,
   input         match_out3774,
   input         match_out3775,
   input         match_out3776,
   input         match_out3777,
   input         match_out3778,
   input         match_out3779,
   input         match_out3780,
   input         match_out3781,
   input         match_out3782,
   input         match_out3783,
   input         match_out3784,
   input         match_out3785,
   input         match_out3786,
   input         match_out3787,
   input         match_out3788,
   input         match_out3789,
   input         match_out3790,
   input         match_out3791,
   input         match_out3792,
   input         match_out3793,
   input         match_out3794,
   input         match_out3795,
   input         match_out3796,
   input         match_out3797,
   input         match_out3798,
   input         match_out3799,
   input         match_out3800,
   input         match_out3801,
   input         match_out3802,
   input         match_out3803,
   input         match_out3804,
   input         match_out3805,
   input         match_out3806,
   input         match_out3807,
   input         match_out3808,
   input         match_out3809,
   input         match_out3810,
   input         match_out3811,
   input         match_out3812,
   input         match_out3813,
   input         match_out3814,
   input         match_out3815,
   input         match_out3816,
   input         match_out3817,
   input         match_out3818,
   input         match_out3819,
   input         match_out3820,
   input         match_out3821,
   input         match_out3822,
   input         match_out3823,
   input         match_out3824,
   input         match_out3825,
   input         match_out3826,
   input         match_out3827,
   input         match_out3828,
   input         match_out3829,
   input         match_out3830,
   input         match_out3831,
   input         match_out3832,
   input         match_out3833,
   input         match_out3834,
   input         match_out3835,
   input         match_out3836,
   input         match_out3837,
   input         match_out3838,
   input         match_out3839,
   input         match_out3840,
   input         match_out3841,
   input         match_out3842,
   input         match_out3843,
   input         match_out3844,
   input         match_out3845,
   input         match_out3846,
   input         match_out3847,
   input         match_out3848,
   input         match_out3849,
   input         match_out3850,
   input         match_out3851,
   input         match_out3852,
   input         match_out3853,
   input         match_out3854,
   input         match_out3855,
   input         match_out3856,
   input         match_out3857,
   input         match_out3858,
   input         match_out3859,
   input         match_out3860,
   input         match_out3861,
   input         match_out3862,
   input         match_out3863,
   input         match_out3864,
   input         match_out3865,
   input         match_out3866,
   input         match_out3867,
   input         match_out3868,
   input         match_out3869,
   input         match_out3870,
   input         match_out3871,
   input         match_out3872,
   input         match_out3873,
   input         match_out3874,
   input         match_out3875,
   input         match_out3876,
   input         match_out3877,
   input         match_out3878,
   input         match_out3879,
   input         match_out3880,
   input         match_out3881,
   input         match_out3882,
   input         match_out3883,
   input         match_out3884,
   input         match_out3885,
   input         match_out3886,
   input         match_out3887,
   input         match_out3888,
   input         match_out3889,
   input         match_out3890,
   input         match_out3891,
   input         match_out3892,
   input         match_out3893,
   input         match_out3894,
   input         match_out3895,
   input         match_out3896,
   input         match_out3897,
   input         match_out3898,
   input         match_out3899,
   input         match_out3900,
   input         match_out3901,
   input         match_out3902,
   input         match_out3903,
   input         match_out3904,
   input         match_out3905,
   input         match_out3906,
   input         match_out3907,
   input         match_out3908,
   input         match_out3909,
   input         match_out3910,
   input         match_out3911,
   input         match_out3912,
   input         match_out3913,
   input         match_out3914,
   input         match_out3915,
   input         match_out3916,
   input         match_out3917,
   input         match_out3918,
   input         match_out3919,
   input         match_out3920,
   input         match_out3921,
   input         match_out3922,
   input         match_out3923,
   input         match_out3924,
   input         match_out3925,
   input         match_out3926,
   input         match_out3927,
   input         match_out3928,
   input         match_out3929,
   input         match_out3930,
   input         match_out3931,
   input         match_out3932,
   input         match_out3933,
   input         match_out3934,
   input         match_out3935,
   input         match_out3936,
   input         match_out3937,
   input         match_out3938,
   input         match_out3939,
   input         match_out3940,
   input         match_out3941,
   input         match_out3942,
   input         match_out3943,
   input         match_out3944,
   input         match_out3945,
   input         match_out3946,
   input         match_out3947,
   input         match_out3948,
   input         match_out3949,
   input         match_out3950,
   input         match_out3951,
   input         match_out3952,
   input         match_out3953,
   input         match_out3954,
   input         match_out3955,
   input         match_out3956,
   input         match_out3957,
   input         match_out3958,
   input         match_out3959,
   input         match_out3960,
   input         match_out3961,
   input         match_out3962,
   input         match_out3963,
   input         match_out3964,
   input         match_out3965,
   input         match_out3966,
   input         match_out3967,
   input         match_out3968,
   input         match_out3969,
   input         match_out3970,
   input         match_out3971,
   input         match_out3972,
   input         match_out3973,
   input         match_out3974,
   input         match_out3975,
   input         match_out3976,
   input         match_out3977,
   input         match_out3978,
   input         match_out3979,
   input         match_out3980,
   input         match_out3981,
   input         match_out3982,
   input         match_out3983,
   input         match_out3984,
   input         match_out3985,
   input         match_out3986,
   input         match_out3987,
   input         match_out3988,
   input         match_out3989,
   input         match_out3990,
   input         match_out3991,
   input         match_out3992,
   input         match_out3993,
   input         match_out3994,
   input         match_out3995,
   input         match_out3996,
   input         match_out3997,
   input         match_out3998,
   input         match_out3999,
   input         match_out4000,
   input         match_out4001,
   input         match_out4002,
   input         match_out4003,
   input         match_out4004,
   input         match_out4005,
   input         match_out4006,
   input         match_out4007,
   input         match_out4008,
   input         match_out4009,
   input         match_out4010,
   input         match_out4011,
   input         match_out4012,
   input         match_out4013,
   input         match_out4014,
   input         match_out4015,
   input         match_out4016,
   input         match_out4017,
   input         match_out4018,
   input         match_out4019,
   input         match_out4020,
   input         match_out4021,
   input         match_out4022,
   input         match_out4023,
   input         match_out4024,
   input         match_out4025,
   input         match_out4026,
   input         match_out4027,
   input         match_out4028,
   input         match_out4029,
   input         match_out4030,
   input         match_out4031,
   input         match_out4032,
   input         match_out4033,
   input         match_out4034,
   input         match_out4035,
   input         match_out4036,
   input         match_out4037,
   input         match_out4038,
   input         match_out4039,
   input         match_out4040,
   input         match_out4041,
   input         match_out4042,
   input         match_out4043,
   input         match_out4044,
   input         match_out4045,
   input         match_out4046,
   input         match_out4047,
   input         match_out4048,
   input         match_out4049,
   input         match_out4050,
   input         match_out4051,
   input         match_out4052,
   input         match_out4053,
   input         match_out4054,
   input         match_out4055,
   input         match_out4056,
   input         match_out4057,
   input         match_out4058,
   input         match_out4059,
   input         match_out4060,
   input         match_out4061,
   input         match_out4062,
   input         match_out4063,
   input         match_out4064,
   input         match_out4065,
   input         match_out4066,
   input         match_out4067,
   input         match_out4068,
   input         match_out4069,
   input         match_out4070,
   input         match_out4071,
   input         match_out4072,
   input         match_out4073,
   input         match_out4074,
   input         match_out4075,
   input         match_out4076,
   input         match_out4077,
   input         match_out4078,
   input         match_out4079,
   input         match_out4080,
   input         match_out4081,
   input         match_out4082,
   input         match_out4083,
   input         match_out4084,
   input         match_out4085,
   input         match_out4086,
   input         match_out4087,
   input         match_out4088,
   input         match_out4089,
   input         match_out4090,
   input         match_out4091,
   input         match_out4092,
   input         match_out4093,
   input         match_out4094,
   input         match_out4095,
   input         match_out4096,
   input         match_out4097,
   input         match_out4098,
   input         match_out4099,
   input         match_out4100,
   input         match_out4101,
   input         match_out4102,
   input         match_out4103,
   input         match_out4104,
   input         match_out4105,
   input         match_out4106,
   input         match_out4107,
   input         match_out4108,
   input         match_out4109,
   input         match_out4110,
   input         match_out4111,
   input         match_out4112,
   input         match_out4113,
   input         match_out4114,
   input         match_out4115,
   input         match_out4116,
   input         match_out4117,
   input         match_out4118,
   input         match_out4119,
   input         match_out4120,
   input         match_out4121,
   input         match_out4122,
   input         match_out4123,
   input         match_out4124,
   input         match_out4125,
   input         match_out4126,
   input         match_out4127,
   input         match_out4128,
   input         match_out4129,
   input         match_out4130,
   input         match_out4131,
   input         match_out4132,
   input         match_out4133,
   input         match_out4134,
   input         match_out4135,
   input         match_out4136,
   input         match_out4137,
   input         match_out4138,
   input         match_out4139,
   input         match_out4140,
   input         match_out4141,
   input         match_out4142,
   input         match_out4143,
   input         match_out4144,
   input         match_out4145,
   input         match_out4146,
   input         match_out4147,
   input         match_out4148,
   input         match_out4149,
   input         match_out4150,
   input         match_out4151,
   input         match_out4152,
   input         match_out4153,
   input         match_out4154,
   input         match_out4155,
   input         match_out4156,
   input         match_out4157,
   input         match_out4158,
   input         match_out4159,
   input         match_out4160,
   input         match_out4161,
   input         match_out4162,
   input         match_out4163,
   input         match_out4164,
   input         match_out4165,
   input         match_out4166,
   input         match_out4167,
   input         match_out4168,
   input         match_out4169,
   input         match_out4170,
   input         match_out4171,
   input         match_out4172,
   input         match_out4173,
   input         match_out4174,
   input         match_out4175,
   input         match_out4176,
   input         match_out4177,
   input         match_out4178,
   input         match_out4179,
   input         match_out4180,
   input         match_out4181,
   input         match_out4182,
   input         match_out4183,
   input         match_out4184,
   input         match_out4185,
   input         match_out4186,
   input         match_out4187,
   input         match_out4188,
   input         match_out4189,
   input         match_out4190,
   input         match_out4191,
   input         match_out4192,
   input         match_out4193,
   input         match_out4194,
   input         match_out4195,
   input         match_out4196,
   input         match_out4197,
   input         match_out4198,
   input         match_out4199,
   input         match_out4200,
   input         match_out4201,
   input         match_out4202,
   input         match_out4203,
   input         match_out4204,
   input         match_out4205,
   input         match_out4206,
   input         match_out4207,
   input         match_out4208,
   input         match_out4209,
   input         match_out4210,
   input         match_out4211,
   input         match_out4212,
   input         match_out4213,
   input         match_out4214,
   input         match_out4215,
   input         match_out4216,
   input         match_out4217,
   input         match_out4218,
   input         match_out4219,
   input         match_out4220,
   input         match_out4221,
   input         match_out4222,
   input         match_out4223,
   input         match_out4224,
   input         match_out4225,
   input         match_out4226,
   input         match_out4227,
   input         match_out4228,
   input         match_out4229,
   input         match_out4230,
   input         match_out4231,
   input         match_out4232,
   input         match_out4233,
   input         match_out4234,
   input         match_out4235,
   input         match_out4236,
   input         match_out4237,
   input         match_out4238,
   input         match_out4239,
   input         match_out4240,
   input         match_out4241,
   input         match_out4242,
   input         match_out4243,
   input         match_out4244,
   input         match_out4245,
   input         match_out4246,
   input         match_out4247,
   input         match_out4248,
   input         match_out4249,
   input         match_out4250,
   input         match_out4251,
   input         match_out4252,
   input         match_out4253,
   input         match_out4254,
   input         match_out4255,
   input         match_out4256,
   input         match_out4257,
   input         match_out4258,
   input         match_out4259,
   input         match_out4260,
   input         match_out4261,
   input         match_out4262,
   input         match_out4263,
   input         match_out4264,
   input         match_out4265,
   input         match_out4266,
   input         match_out4267,
   input         match_out4268,
   input         match_out4269,
   input         match_out4270,
   input         match_out4271,
   input         match_out4272,
   input         match_out4273,
   input         match_out4274,
   input         match_out4275,
   input         match_out4276,
   input         match_out4277,
   input         match_out4278,
   input         match_out4279,
   input         match_out4280,
   input         match_out4281,
   input         match_out4282,
   input         match_out4283,
   input         match_out4284,
   input         match_out4285,
   input         match_out4286,
   input         match_out4287,
   input         match_out4288,
   input         match_out4289,
   input         match_out4290,
   input         match_out4291,
   input         match_out4292,
   input         match_out4293,
   input         match_out4294,
   input         match_out4295,
   input         match_out4296,
   input         match_out4297,
   input         match_out4298,
   input         match_out4299,
   input         match_out4300,
   input         match_out4301,
   input         match_out4302,
   input         match_out4303,
   input         match_out4304,
   input         match_out4305,
   input         match_out4306,
   input         match_out4307,
   input         match_out4308,
   input         match_out4309,
   input         match_out4310,
   input         match_out4311,
   input         match_out4312,
   input         match_out4313,
   input         match_out4314,
   input         match_out4315,
   input         match_out4316,
   input         match_out4317,
   input         match_out4318,
   input         match_out4319,
   input         match_out4320,
   input         match_out4321,
   input         match_out4322,
   input         match_out4323,
   input         match_out4324,
   input         match_out4325,
   input         match_out4326,
   input         match_out4327,
   input         match_out4328,
   input         match_out4329,
   input         match_out4330,
   input         match_out4331,
   input         match_out4332,
   input         match_out4333,
   input         match_out4334,
   input         match_out4335,
   input         match_out4336,
   input         match_out4337,
   input         match_out4338,
   input         match_out4339,
   input         match_out4340,
   input         match_out4341,
   input         match_out4342,
   input         match_out4343,
   input         match_out4344,
   input         match_out4345,
   input         match_out4346,
   input         match_out4347,
   input         match_out4348,
   input         match_out4349,
   input         match_out4350,
   input         match_out4351,
   input         match_out4352,
   input         match_out4353,
   input         match_out4354,
   input         match_out4355,
   input         match_out4356,
   input         match_out4357,
   input         match_out4358,
   input         match_out4359,
   input         match_out4360,
   input         match_out4361,
   input         match_out4362,
   input         match_out4363,
   input         match_out4364,
   input         match_out4365,
   input         match_out4366,
   input         match_out4367,
   input         match_out4368,
   input         match_out4369,
   input         match_out4370,
   input         match_out4371,
   input         match_out4372,
   input         match_out4373,
   input         match_out4374,
   input         match_out4375,
   input         match_out4376,
   input         match_out4377,
   input         match_out4378,
   input         match_out4379,
   input         match_out4380,
   input         match_out4381,
   input         match_out4382,
   input         match_out4383,
   input         match_out4384,
   input         match_out4385,
   input         match_out4386,
   input         match_out4387,
   input         match_out4388,
   input         match_out4389,
   input         match_out4390,
   input         match_out4391,
   input         match_out4392,
   input         match_out4393,
   input         match_out4394,
   input         match_out4395,
   input         match_out4396,
   input         match_out4397,
   input         match_out4398,
   input         match_out4399,
   input         match_out4400,
   input         match_out4401,
   input         match_out4402,
   input         match_out4403,
   input         match_out4404,
   input         match_out4405,
   input         match_out4406,
   input         match_out4407,
   input         match_out4408,
   input         match_out4409,
   input         match_out4410,
   input         match_out4411,
   input         match_out4412,
   input         match_out4413,
   input         match_out4414,
   input         match_out4415,
   input         match_out4416,
   input         match_out4417,
   input         match_out4418,
   input         match_out4419,
   input         match_out4420,
   input         match_out4421,
   input         match_out4422,
   input         match_out4423,
   input         match_out4424,
   input         match_out4425,
   input         match_out4426,
   input         match_out4427,
   input         match_out4428,
   input         match_out4429,
   input         match_out4430,
   input         match_out4431,
   input         match_out4432,
   input         match_out4433,
   input         match_out4434,
   input         match_out4435,
   input         match_out4436,
   input         match_out4437,
   input         match_out4438,
   input         match_out4439,
   input         match_out4440,
   input         match_out4441,
   input         match_out4442,
   input         match_out4443,
   input         match_out4444,
   input         match_out4445,
   input         match_out4446,
   input         match_out4447,
   input         match_out4448,
   input         match_out4449,
   input         match_out4450,
   input         match_out4451,
   input         match_out4452,
   input         match_out4453,
   input         match_out4454,
   input         match_out4455,
   input         match_out4456,
   input         match_out4457,
   input         match_out4458,
   input         match_out4459,
   input         match_out4460,
   input         match_out4461,
   input         match_out4462,
   input         match_out4463,
   input         match_out4464,
   input         match_out4465,
   input         match_out4466,
   input         match_out4467,
   input         match_out4468,
   input         match_out4469,
   input         match_out4470,
   input         match_out4471,
   input         match_out4472,
   input         match_out4473,
   input         match_out4474,
   input         match_out4475,
   input         match_out4476,
   input         match_out4477,
   input         match_out4478,
   input         match_out4479,
   input         match_out4480,
   input         match_out4481,
   input         match_out4482,
   input         match_out4483,
   input         match_out4484,
   input         match_out4485,
   input         match_out4486,
   input         match_out4487,
   input         match_out4488,
   input         match_out4489,
   input         match_out4490,
   input         match_out4491,
   input         match_out4492,
   input         match_out4493,
   input         match_out4494,
   input         match_out4495,
   input         match_out4496,
   input         match_out4497,
   input         match_out4498,
   input         match_out4499,
   input         match_out4500,
   input         match_out4501,
   input         match_out4502,
   input         match_out4503,
   input         match_out4504,
   input         match_out4505,
   input         match_out4506,
   input         match_out4507,
   input         match_out4508,
   input         match_out4509,
   input         match_out4510,
   input         match_out4511,
   input         match_out4512,
   input         match_out4513,
   input         match_out4514,
   input         match_out4515,
   input         match_out4516,
   input         match_out4517,
   input         match_out4518,
   input         match_out4519,
   input         match_out4520,
   input         match_out4521,
   input         match_out4522,
   input         match_out4523,
   input         match_out4524,
   input         match_out4525,
   input         match_out4526,
   input         match_out4527,
   input         match_out4528,
   input         match_out4529,
   input         match_out4530,
   input         match_out4531,
   input         match_out4532,
   input         match_out4533,
   input         match_out4534,
   input         match_out4535,
   input         match_out4536,
   input         match_out4537,
   input         match_out4538,
   input         match_out4539,
   input         match_out4540,
   input         match_out4541,
   input         match_out4542,
   input         match_out4543,
   input         match_out4544,
   input         match_out4545,
   input         match_out4546,
   input         match_out4547,
   input         match_out4548,
   input         match_out4549,
   input         match_out4550,
   input         match_out4551,
   input         match_out4552,
   input         match_out4553,
   input         match_out4554,
   input         match_out4555,
   input         match_out4556,
   input         match_out4557,
   input         match_out4558,
   input         match_out4559,
   input         match_out4560,
   input         match_out4561,
   input         match_out4562,
   input         match_out4563,
   input         match_out4564,
   input         match_out4565,
   input         match_out4566,
   input         match_out4567,
   input         match_out4568,
   input         match_out4569,
   input         match_out4570,
   input         match_out4571,
   input         match_out4572,
   input         match_out4573,
   input         match_out4574,
   input         match_out4575,
   input         match_out4576,
   input         match_out4577,
   input         match_out4578,
   input         match_out4579,
   input         match_out4580,
   input         match_out4581,
   input         match_out4582,
   input         match_out4583,
   input         match_out4584,
   input         match_out4585,
   input         match_out4586,
   input         match_out4587,
   input         match_out4588,
   input         match_out4589,
   input         match_out4590,
   input         match_out4591,
   input         match_out4592,
   input         match_out4593,
   input         match_out4594,
   input         match_out4595,
   input         match_out4596,
   input         match_out4597,
   input         match_out4598,
   input         match_out4599,
   input         match_out4600,
   input         match_out4601,
   input         match_out4602,
   input         match_out4603,
   input         match_out4604,
   input         match_out4605,
   input         match_out4606,
   input         match_out4607,
   input         match_out4608,
   input         match_out4609,
   input         match_out4610,
   input         match_out4611,
   input         match_out4612,
   input         match_out4613,
   input         match_out4614,
   input         match_out4615,
   input         match_out4616,
   input         match_out4617,
   input         match_out4618,
   input         match_out4619,
   input         match_out4620,
   input         match_out4621,
   input         match_out4622,
   input         match_out4623,
   input         match_out4624,
   input         match_out4625,
   input         match_out4626,
   input         match_out4627,
   input         match_out4628,
   input         match_out4629,
   input         match_out4630,
   input         match_out4631,
   input         match_out4632,
   input         match_out4633,
   input         match_out4634,
   input         match_out4635,
   input         match_out4636,
   input         match_out4637,
   input         match_out4638,
   input         match_out4639,
   input         match_out4640,
   input         match_out4641,
   input         match_out4642,
   input         match_out4643,
   input         match_out4644,
   input         match_out4645,
   input         match_out4646,
   input         match_out4647,
   input         match_out4648,
   input         match_out4649,
   input         match_out4650,
   input         match_out4651,
   input         match_out4652,
   input         match_out4653,
   input         match_out4654,
   input         match_out4655,
   input         match_out4656,
   input         match_out4657,
   input         match_out4658,
   input         match_out4659,
   input         match_out4660,
   input         match_out4661,
   input         match_out4662,
   input         match_out4663,
   input         match_out4664,
   input         match_out4665,
   input         match_out4666,
   input         match_out4667,
   input         match_out4668,
   input         match_out4669,
   input         match_out4670,
   input         match_out4671,
   input         match_out4672,
   input         match_out4673,
   input         match_out4674,
   input         match_out4675,
   input         match_out4676,
   input         match_out4677,
   input         match_out4678,
   input         match_out4679,
   input         match_out4680,
   input         match_out4681,
   input         match_out4682,
   input         match_out4683,
   input         match_out4684,
   input         match_out4685,
   input         match_out4686,
   input         match_out4687,
   input         match_out4688,
   input         match_out4689,
   input         match_out4690,
   input         match_out4691,
   input         match_out4692,
   input         match_out4693,
   input         match_out4694,
   input         match_out4695,
   input         match_out4696,
   input         match_out4697,
   input         match_out4698,
   input         match_out4699,
   input         match_out4700,
   input         match_out4701,
   input         match_out4702,
   input         match_out4703,
   input         match_out4704,
   input         match_out4705,
   input         match_out4706,
   input         match_out4707,
   input         match_out4708,
   input         match_out4709,
   input         match_out4710,
   input         match_out4711,
   input         match_out4712,
   input         match_out4713,
   input         match_out4714,
   input         match_out4715,
   input         match_out4716,
   input         match_out4717,
   input         match_out4718,
   input         match_out4719,
   input         match_out4720,
   input         match_out4721,
   input         match_out4722,
   input         match_out4723,
   input         match_out4724,
   input         match_out4725,
   input         match_out4726,
   input         match_out4727,
   input         match_out4728,
   input         match_out4729,
   input         match_out4730,
   input         match_out4731,
   input         match_out4732,
   input         match_out4733,
   input         match_out4734,
   input         match_out4735,
   input         match_out4736,
   input         match_out4737,
   input         match_out4738,
   input         match_out4739,
   input         match_out4740,
   input         match_out4741,
   input         match_out4742,
   input         match_out4743,
   input         match_out4744,
   input         match_out4745,
   input         match_out4746,
   input         match_out4747,
   input         match_out4748,
   input         match_out4749,
   input         match_out4750,
   input         match_out4751,
   input         match_out4752,
   input         match_out4753,
   input         match_out4754,
   input         match_out4755,
   input         match_out4756,
   input         match_out4757,
   input         match_out4758,
   input         match_out4759,
   input         match_out4760,
   input         match_out4761,
   input         match_out4762,
   input         match_out4763,
   input         match_out4764,
   input         match_out4765,
   input         match_out4766,
   input         match_out4767,
   input         match_out4768,
   input         match_out4769,
   input         match_out4770,
   input         match_out4771,
   input         match_out4772,
   input         match_out4773,
   input         match_out4774,
   input         match_out4775,
   input         match_out4776,
   input         match_out4777,
   input         match_out4778,
   input         match_out4779,
   input         match_out4780,
   input         match_out4781,
   input         match_out4782,
   input         match_out4783,
   input         match_out4784,
   input         match_out4785,
   input         match_out4786,
   input         match_out4787,
   input         match_out4788,
   input         match_out4789,
   input         match_out4790,
   input         match_out4791,
   input         match_out4792,
   input         match_out4793,
   input         match_out4794,
   input         match_out4795,
   input         match_out4796,
   input         match_out4797,
   input         match_out4798,
   input         match_out4799,
   input         match_out4800,
   input         match_out4801,
   input         match_out4802,
   input         match_out4803,
   input         match_out4804,
   input         match_out4805,
   input         match_out4806,
   input         match_out4807,
   input         match_out4808,
   input         match_out4809,
   input         match_out4810,
   input         match_out4811,
   input         match_out4812,
   input         match_out4813,
   input         match_out4814,
   input         match_out4815,
   input         match_out4816,
   input         match_out4817,
   input         match_out4818,
   input         match_out4819,
   input         match_out4820,
   input         match_out4821,
   input         match_out4822,
   input         match_out4823,
   input         match_out4824,
   input         match_out4825,
   input         match_out4826,
   input         match_out4827,
   input         match_out4828,
   input         match_out4829,
   input         match_out4830,
   input         match_out4831,
   input         match_out4832,
   input         match_out4833,
   input         match_out4834,
   input         match_out4835,
   input         match_out4836,
   input         match_out4837,
   input         match_out4838,
   input         match_out4839,
   input         match_out4840,
   input         match_out4841,
   input         match_out4842,
   input         match_out4843,
   input         match_out4844,
   input         match_out4845,
   input         match_out4846,
   input         match_out4847,
   input         match_out4848,
   input         match_out4849,
   input         match_out4850,
   input         match_out4851,
   input         match_out4852,
   input         match_out4853,
   input         match_out4854,
   input         match_out4855,
   input         match_out4856,
   input         match_out4857,
   input         match_out4858,
   input         match_out4859,
   input         match_out4860,
   input         match_out4861,
   input         match_out4862,
   input         match_out4863,
   input         match_out4864,
   input         match_out4865,
   input         match_out4866,
   input         match_out4867,
   input         match_out4868,
   input         match_out4869,
   input         match_out4870,
   input         match_out4871,
   input         match_out4872,
   input         match_out4873,
   input         match_out4874,
   input         match_out4875,
   input         match_out4876,
   input         match_out4877,
   input         match_out4878,
   input         match_out4879,
   input         match_out4880,
   input         match_out4881,
   input         match_out4882,
   input         match_out4883,
   input         match_out4884,
   input         match_out4885,
   input         match_out4886,
   input         match_out4887,
   input         match_out4888,
   input         match_out4889,
   input         match_out4890,
   input         match_out4891,
   input         match_out4892,
   input         match_out4893,
   input         match_out4894,
   input         match_out4895,
   input         match_out4896,
   input         match_out4897,
   input         match_out4898,
   input         match_out4899,
   input         match_out4900,
   input         match_out4901,
   input         match_out4902,
   input         match_out4903,
   input         match_out4904,
   input         match_out4905,
   input         match_out4906,
   input         match_out4907,
   input         match_out4908,
   input         match_out4909,
   input         match_out4910,
   input         match_out4911,
   input         match_out4912,
   input         match_out4913,
   input         match_out4914,
   input         match_out4915,
   input         match_out4916,
   input         match_out4917,
   input         match_out4918,
   input         match_out4919,
   input         match_out4920,
   input         match_out4921,
   input         match_out4922,
   input         match_out4923,
   input         match_out4924,
   input         match_out4925,
   input         match_out4926,
   input         match_out4927,
   input         match_out4928,
   input         match_out4929,
   input         match_out4930,
   input         match_out4931,
   input         match_out4932,
   input         match_out4933,
   input         match_out4934,
   input         match_out4935,
   input         match_out4936,
   input         match_out4937,
   input         match_out4938,
   input         match_out4939,
   input         match_out4940,
   input         match_out4941,
   input         match_out4942,
   input         match_out4943,
   input         match_out4944,
   input         match_out4945,
   input         match_out4946,
   input         match_out4947,
   input         match_out4948,
   input         match_out4949,
   input         match_out4950,
   input         match_out4951,
   input         match_out4952,
   input         match_out4953,
   input         match_out4954,
   input         match_out4955,
   input         match_out4956,
   input         match_out4957,
   input         match_out4958,
   input         match_out4959,
   input         match_out4960,
   input         match_out4961,
   input         match_out4962,
   input         match_out4963,
   input         match_out4964,
   input         match_out4965,
   input         match_out4966,
   input         match_out4967,
   input         match_out4968,
   input         match_out4969,
   input         match_out4970,
   input         match_out4971,
   input         match_out4972,
   input         match_out4973,
   input         match_out4974,
   input         match_out4975,
   input         match_out4976,
   input         match_out4977,
   input         match_out4978,
   input         match_out4979,
   input         match_out4980,
   input         match_out4981,
   input         match_out4982,
   input         match_out4983,
   input         match_out4984,
   input         match_out4985,
   input         match_out4986,
   input         match_out4987,
   input         match_out4988,
   input         match_out4989,
   input         match_out4990,
   input         match_out4991,
   input         match_out4992,
   input         match_out4993,
   input         match_out4994,
   input         match_out4995,
   input         match_out4996,
   input         match_out4997,
   input         match_out4998,
   input         match_out4999,
   input         match_out5000,
   input         match_out5001,
   input         match_out5002,
   input         match_out5003,
   input         match_out5004,
   input         match_out5005,
   input         match_out5006,
   input         match_out5007,
   input         match_out5008,
   input         match_out5009,
   input         match_out5010,
   input         match_out5011,
   input         match_out5012,
   input         match_out5013,
   input         match_out5014,
   input         match_out5015,
   input         match_out5016,
   input         match_out5017,
   input         match_out5018,
   input         match_out5019,
   input         match_out5020,
   input         match_out5021,
   input         match_out5022,
   input         match_out5023,
   input         match_out5024,
   input         match_out5025,
   input         match_out5026,
   input         match_out5027,
   input         match_out5028,
   input         match_out5029,
   input         match_out5030,
   input         match_out5031,
   input         match_out5032,
   input         match_out5033,
   input         match_out5034,
   input         match_out5035,
   input         match_out5036,
   input         match_out5037,
   input         match_out5038,
   input         match_out5039,
   input         match_out5040,
   input         match_out5041,
   input         match_out5042,
   input         match_out5043,
   input         match_out5044,
   input         match_out5045,
   input         match_out5046,
   input         match_out5047,
   input         match_out5048,
   input         match_out5049,
   input         match_out5050,
   input         match_out5051,
   input         match_out5052,
   input         match_out5053,
   input         match_out5054,
   input         match_out5055,
   input         match_out5056,
   input         match_out5057,
   input         match_out5058,
   input         match_out5059,
   input         match_out5060,
   input         match_out5061,
   input         match_out5062,
   input         match_out5063,
   input         match_out5064,
   input         match_out5065,
   input         match_out5066,
   input         match_out5067,
   input         match_out5068,
   input         match_out5069,
   input         match_out5070,
   input         match_out5071,
   input         match_out5072,
   input         match_out5073,
   input         match_out5074,
   input         match_out5075,
   input         match_out5076,
   input         match_out5077,
   input         match_out5078,
   input         match_out5079,
   input         match_out5080,
   input         match_out5081,
   input         match_out5082,
   input         match_out5083,
   input         match_out5084,
   input         match_out5085,
   input         match_out5086,
   input         match_out5087,
   input         match_out5088,
   input         match_out5089,
   input         match_out5090,
   input         match_out5091,
   input         match_out5092,
   input         match_out5093,
   input         match_out5094,
   input         match_out5095,
   input         match_out5096,
   input         match_out5097,
   input         match_out5098,
   input         match_out5099,
   input         match_out5100,
   input         match_out5101,
   input         match_out5102,
   input         match_out5103,
   input         match_out5104,
   input         match_out5105,
   input         match_out5106,
   input         match_out5107,
   input         match_out5108,
   input         match_out5109,
   input         match_out5110,
   input         match_out5111,
   input         match_out5112,
   input         match_out5113,
   input         match_out5114,
   input         match_out5115,
   input         match_out5116,
   input         match_out5117,
   input         match_out5118,
   input         match_out5119,
   input         match_out5120,
   input         match_out5121,
   input         match_out5122,
   input         match_out5123,
   input         match_out5124,
   input         match_out5125,
   input         match_out5126,
   input         match_out5127,
   input         match_out5128,
   input         match_out5129,
   input         match_out5130,
   input         match_out5131,
   input         match_out5132,
   input         match_out5133,
   input         match_out5134,
   input         match_out5135,
   input         match_out5136,
   input         match_out5137,
   input         match_out5138,
   input         match_out5139,
   input         match_out5140,
   input         match_out5141,
   input         match_out5142,
   input         match_out5143,
   input         match_out5144,
   input         match_out5145,
   input         match_out5146,
   input         match_out5147,
   input         match_out5148,
   input         match_out5149,
   input         match_out5150,
   input         match_out5151,
   input         match_out5152,
   input         match_out5153,
   input         match_out5154,
   input         match_out5155,
   input         match_out5156,
   input         match_out5157,
   input         match_out5158,
   input         match_out5159,
   input         match_out5160,
   input         match_out5161,
   input         match_out5162,
   input         match_out5163,
   input         match_out5164,
   input         match_out5165,
   input         match_out5166,
   input         match_out5167,
   input         match_out5168,
   input         match_out5169,
   input         match_out5170,
   input         match_out5171,
   input         match_out5172,
   input         match_out5173,
   input         match_out5174,
   input         match_out5175,
   input         match_out5176,
   input         match_out5177,
   input         match_out5178,
   input         match_out5179,
   input         match_out5180,
   input         match_out5181,
   input         match_out5182,
   input         match_out5183,
   input         match_out5184,
   input         match_out5185,
   input         match_out5186,
   input         match_out5187,
   input         match_out5188,
   input         match_out5189,
   input         match_out5190,
   input         match_out5191,
   input         match_out5192,
   input         match_out5193,
   input         match_out5194,
   input         match_out5195,
   input         match_out5196,
   input         match_out5197,
   input         match_out5198,
   input         match_out5199,
   input         match_out5200,
   input         match_out5201,
   input         match_out5202,
   input         match_out5203,
   input         match_out5204,
   input         match_out5205,
   input         match_out5206,
   input         match_out5207,
   input         match_out5208,
   input         match_out5209,
   input         match_out5210,
   input         match_out5211,
   input         match_out5212,
   input         match_out5213,
   input         match_out5214,
   input         match_out5215,
   input         match_out5216,
   input         match_out5217,
   input         match_out5218,
   input         match_out5219,
   input         match_out5220,
   input         match_out5221,
   input         match_out5222,
   input         match_out5223,
   input         match_out5224,
   input         match_out5225,
   input         match_out5226,
   input         match_out5227,
   input         match_out5228,
   input         match_out5229,
   input         match_out5230,
   input         match_out5231,
   input         match_out5232,
   input         match_out5233,
   input         match_out5234,
   input         match_out5235,
   input         match_out5236,
   input         match_out5237,
   input         match_out5238,
   input         match_out5239,
   input         match_out5240,
   input         match_out5241,
   input         match_out5242,
   input         match_out5243,
   input         match_out5244,
   input         match_out5245,
   input         match_out5246,
   input         match_out5247,
   input         match_out5248,
   input         match_out5249,
   input         match_out5250,
   input         match_out5251,
   input         match_out5252,
   input         match_out5253,
   input         match_out5254,
   input         match_out5255,
   input         match_out5256,
   input         match_out5257,
   input         match_out5258,
   input         match_out5259,
   input         match_out5260,
   input         match_out5261,
   input         match_out5262,
   input         match_out5263,
   input         match_out5264,
   input         match_out5265,
   input         match_out5266,
   input         match_out5267,
   input         match_out5268,
   input         match_out5269,
   input         match_out5270,
   input         match_out5271,
   input         match_out5272,
   input         match_out5273,
   input         match_out5274,
   input         match_out5275,
   input         match_out5276,
   input         match_out5277,
   input         match_out5278,
   input         match_out5279,
   input         match_out5280,
   input         match_out5281,
   input         match_out5282,
   input         match_out5283,
   input         match_out5284,
   input         match_out5285,
   input         match_out5286,
   input         match_out5287,
   input         match_out5288,
   input         match_out5289,
   input         match_out5290,
   input         match_out5291,
   input         match_out5292,
   input         match_out5293,
   input         match_out5294,
   input         match_out5295,
   input         match_out5296,
   input         match_out5297,
   input         match_out5298,
   input         match_out5299,
   input         match_out5300,
   input         match_out5301,
   input         match_out5302,
   input         match_out5303,
   input         match_out5304,
   input         match_out5305,
   input         match_out5306,
   input         match_out5307,
   input         match_out5308,
   input         match_out5309,
   input         match_out5310,
   input         match_out5311,
   input         match_out5312,
   input         match_out5313,
   input         match_out5314,
   input         match_out5315,
   input         match_out5316,
   input         match_out5317,
   input         match_out5318,
   input         match_out5319,
   input         match_out5320,
   input         match_out5321,
   input         match_out5322,
   input         match_out5323,
   input         match_out5324,
   input         match_out5325,
   input         match_out5326,
   input         match_out5327,
   input         match_out5328,
   input         match_out5329,
   input         match_out5330,
   input         match_out5331,
   input         match_out5332,
   input         match_out5333,
   input         match_out5334,
   input         match_out5335,
   input         match_out5336,
   input         match_out5337,
   input         match_out5338,
   input         match_out5339,
   input         match_out5340,
   input         match_out5341,
   input         match_out5342,
   input         match_out5343,
   input         match_out5344,
   input         match_out5345,
   input         match_out5346,
   input         match_out5347,
   input         match_out5348,
   input         match_out5349,
   input         match_out5350,
   input         match_out5351,
   input         match_out5352,
   input         match_out5353,
   input         match_out5354,
   input         match_out5355,
   input         match_out5356,
   input         match_out5357,
   input         match_out5358,
   input         match_out5359,
   input         match_out5360,
   input         match_out5361,
   input         match_out5362,
   input         match_out5363,
   input         match_out5364,
   input         match_out5365,
   input         match_out5366,
   input         match_out5367,
   input         match_out5368,
   input         match_out5369,
   input         match_out5370,
   input         match_out5371,
   input         match_out5372,
   input         match_out5373,
   input         match_out5374,
   input         match_out5375,
   input         match_out5376,
   input         match_out5377,
   input         match_out5378,
   input         match_out5379,
   input         match_out5380,
   input         match_out5381,
   input         match_out5382,
   input         match_out5383,
   input         match_out5384,
   input         match_out5385,
   input         match_out5386,
   input         match_out5387,
   input         match_out5388,
   input         match_out5389,
   input         match_out5390,
   input         match_out5391,
   input         match_out5392,
   input         match_out5393,
   input         match_out5394,
   input         match_out5395,
   input         match_out5396,
   input         match_out5397,
   input         match_out5398,
   input         match_out5399,
   input         match_out5400,
   input         match_out5401,
   input         match_out5402,
   input         match_out5403,
   input         match_out5404,
   input         match_out5405,
   input         match_out5406,
   input         match_out5407,
   input         match_out5408,
   input         match_out5409,
   input         match_out5410,
   input         match_out5411,
   input         match_out5412,
   input         match_out5413,
   input         match_out5414,
   input         match_out5415,
   input         match_out5416,
   input         match_out5417,
   input         match_out5418,
   input         match_out5419,
   input         match_out5420,
   input         match_out5421,
   input         match_out5422,
   input         match_out5423,
   input         match_out5424,
   input         match_out5425,
   input         match_out5426,
   input         match_out5427,
   input         match_out5428,
   input         match_out5429,
   input         match_out5430,
   input         match_out5431,
   input         match_out5432,
   input         match_out5433,
   input         match_out5434,
   input         match_out5435,
   input         match_out5436,
   input         match_out5437,
   input         match_out5438,
   input         match_out5439,
   input         match_out5440,
   input         match_out5441,
   input         match_out5442,
   input         match_out5443,
   input         match_out5444,
   input         match_out5445,
   input         match_out5446,
   input         match_out5447,
   input         match_out5448,
   input         match_out5449,
   input         match_out5450,
   input         match_out5451,
   input         match_out5452,
   input         match_out5453,
   input         match_out5454,
   input         match_out5455,
   input         match_out5456,
   input         match_out5457,
   input         match_out5458,
   input         match_out5459,
   input         match_out5460,
   input         match_out5461,
   input         match_out5462,
   input         match_out5463,
   input         match_out5464,
   input         match_out5465,
   input         match_out5466,
   input         match_out5467,
   input         match_out5468,
   input         match_out5469,
   input         match_out5470,
   input         match_out5471,
   input         match_out5472,
   input         match_out5473,
   input         match_out5474,
   input         match_out5475,
   input         match_out5476,
   input         match_out5477,
   input         match_out5478,
   input         match_out5479,
   input         match_out5480,
   input         match_out5481,
   input         match_out5482,
   input         match_out5483,
   input         match_out5484,
   input         match_out5485,
   input         match_out5486,
   input         match_out5487,
   input         match_out5488,
   input         match_out5489,
   input         match_out5490,
   input         match_out5491,
   input         match_out5492,
   input         match_out5493,
   input         match_out5494,
   input         match_out5495,
   input         match_out5496,
   input         match_out5497,
   input         match_out5498,
   input         match_out5499,
   input         match_out5500,
   input         match_out5501,
   input         match_out5502,
   input         match_out5503,
   input         match_out5504,
   input         match_out5505,
   input         match_out5506,
   input         match_out5507,
   input         match_out5508,
   input         match_out5509,
   input         match_out5510,
   input         match_out5511,
   input         match_out5512,
   input         match_out5513,
   input         match_out5514,
   input         match_out5515,
   input         match_out5516,
   input         match_out5517,
   input         match_out5518,
   input         match_out5519,
   input         match_out5520,
   input         match_out5521,
   input         match_out5522,
   input         match_out5523,
   input         match_out5524,
   input         match_out5525,
   input         match_out5526,
   input         match_out5527,
   input         match_out5528,
   input         match_out5529,
   input         match_out5530,
   input         match_out5531,
   input         match_out5532,
   input         match_out5533,
   input         match_out5534,
   input         match_out5535,
   input         match_out5536,
   input         match_out5537,
   input         match_out5538,
   input         match_out5539,
   input         match_out5540,
   input         match_out5541,
   input         match_out5542,
   input         match_out5543,
   input         match_out5544,
   input         match_out5545,
   input         match_out5546,
   input         match_out5547,
   input         match_out5548,
   input         match_out5549,
   input         match_out5550,
   input         match_out5551,
   input         match_out5552,
   input         match_out5553,
   input         match_out5554,
   input         match_out5555,
   input         match_out5556,
   input         match_out5557,
   input         match_out5558,
   input         match_out5559,
   input         match_out5560,
   input         match_out5561,
   input         match_out5562,
   input         match_out5563,
   input         match_out5564,
   input         match_out5565,
   input         match_out5566,
   input         match_out5567,
   input         match_out5568,
   input         match_out5569,
   input         match_out5570,
   input         match_out5571,
   input         match_out5572,
   input         match_out5573,
   input         match_out5574,
   input         match_out5575,
   input         match_out5576,
   input         match_out5577,
   input         match_out5578,
   input         match_out5579,
   input         match_out5580,
   input         match_out5581,
   input         match_out5582,
   input         match_out5583,
   input         match_out5584,
   input         match_out5585,
   input         match_out5586,
   input         match_out5587,
   input         match_out5588,
   input         match_out5589,
   input         match_out5590,
   input         match_out5591,
   input         match_out5592,
   input         match_out5593,
   input         match_out5594,
   input         match_out5595,
   input         match_out5596,
   input         match_out5597,
   input         match_out5598,
   input         match_out5599,
   input         match_out5600,
   input         match_out5601,
   input         match_out5602,
   input         match_out5603,
   input         match_out5604,
   input         match_out5605,
   input         match_out5606,
   input         match_out5607,
   input         match_out5608,
   input         match_out5609,
   input         match_out5610,
   input         match_out5611,
   input         match_out5612,
   input         match_out5613,
   input         match_out5614,
   input         match_out5615,
   input         match_out5616,
   input         match_out5617,
   input         match_out5618,
   input         match_out5619,
   input         match_out5620,
   input         match_out5621,
   input         match_out5622,
   input         match_out5623,
   input         match_out5624,
   input         match_out5625,
   input         match_out5626,
   input         match_out5627,
   input         match_out5628,
   input         match_out5629,
   input         match_out5630,
   input         match_out5631,
   input         match_out5632,
   input         match_out5633,
   input         match_out5634,
   input         match_out5635,
   input         match_out5636,
   input         match_out5637,
   input         match_out5638,
   input         match_out5639,
   input         match_out5640,
   input         match_out5641,
   input         match_out5642,
   input         match_out5643,
   input         match_out5644,
   input         match_out5645,
   input         match_out5646,
   input         match_out5647,
   input         match_out5648,
   input         match_out5649,
   input         match_out5650,
   input         match_out5651,
   input         match_out5652,
   input         match_out5653,
   input         match_out5654,
   input         match_out5655,
   input         match_out5656,
   input         match_out5657,
   input         match_out5658,
   input         match_out5659,
   input         match_out5660,
   input         match_out5661,
   input         match_out5662,
   input         match_out5663,
   input         match_out5664,
   input         match_out5665,
   input         match_out5666,
   input         match_out5667,
   input         match_out5668,
   input         match_out5669,
   input         match_out5670,
   input         match_out5671,
   input         match_out5672,
   input         match_out5673,
   input         match_out5674,
   input         match_out5675,
   input         match_out5676,
   input         match_out5677,
   input         match_out5678,
   input         match_out5679,
   input         match_out5680,
   input         match_out5681,
   input         match_out5682,
   input         match_out5683,
   input         match_out5684,
   input         match_out5685,
   input         match_out5686,
   input         match_out5687,
   input         match_out5688,
   input         match_out5689,
   input         match_out5690,
   input         match_out5691,
   input         match_out5692,
   input         match_out5693,
   input         match_out5694,
   input         match_out5695,
   input         match_out5696,
   input         match_out5697,
   input         match_out5698,
   input         match_out5699,
   input         match_out5700,
   input         match_out5701,
   input         match_out5702,
   input         match_out5703,
   input         match_out5704,
   input         match_out5705,
   input         match_out5706,
   input         match_out5707,
   input         match_out5708,
   input         match_out5709,
   input         match_out5710,
   input         match_out5711,
   input         match_out5712,
   input         match_out5713,
   input         match_out5714,
   input         match_out5715,
   input         match_out5716,
   input         match_out5717,
   input         match_out5718,
   input         match_out5719,
   input         match_out5720,
   input         match_out5721,
   input         match_out5722,
   input         match_out5723,
   input         match_out5724,
   input         match_out5725,
   input         match_out5726,
   input         match_out5727,
   input         match_out5728,
   input         match_out5729,
   input         match_out5730,
   input         match_out5731,
   input         match_out5732,
   input         match_out5733,
   input         match_out5734,
   input         match_out5735,
   input         match_out5736,
   input         match_out5737,
   input         match_out5738,
   input         match_out5739,
   input         match_out5740,
   input         match_out5741,
   input         match_out5742,
   input         match_out5743,
   input         match_out5744,
   input         match_out5745,
   input         match_out5746,
   input         match_out5747,
   input         match_out5748,
   input         match_out5749,
   input         match_out5750,
   input         match_out5751,
   input         match_out5752,
   input         match_out5753,
   input         match_out5754,
   input         match_out5755,
   input         match_out5756,
   input         match_out5757,
   input         match_out5758,
   input         match_out5759,
   input         match_out5760,
   input         match_out5761,
   input         match_out5762,
   input         match_out5763,
   input         match_out5764,
   input         match_out5765,
   input         match_out5766,
   input         match_out5767,
   input         match_out5768,
   input         match_out5769,
   input         match_out5770,
   input         match_out5771,
   input         match_out5772,
   input         match_out5773,
   input         match_out5774,
   input         match_out5775,
   input         match_out5776,
   input         match_out5777,
   input         match_out5778,
   input         match_out5779,
   input         match_out5780,
   input         match_out5781,
   input         match_out5782,
   input         match_out5783,
   input         match_out5784,
   input         match_out5785,
   input         match_out5786,
   input         match_out5787,
   input         match_out5788,
   input         match_out5789,
   input         match_out5790,
   input         match_out5791,
   input         match_out5792,
   input         match_out5793,
   input         match_out5794,
   input         match_out5795,
   input         match_out5796,
   input         match_out5797,
   input         match_out5798,
   input         match_out5799,
   input         match_out5800,
   input         match_out5801,
   input         match_out5802,
   input         match_out5803,
   input         match_out5804,
   input         match_out5805,
   input         match_out5806,
   input         match_out5807,
   input         match_out5808,
   input         match_out5809,
   input         match_out5810,
   input         match_out5811,
   input         match_out5812,
   input         match_out5813,
   input         match_out5814,
   input         match_out5815,
   input         match_out5816,
   input         match_out5817,
   input         match_out5818,
   input         match_out5819,
   input         match_out5820,
   input         match_out5821,
   input         match_out5822,
   input         match_out5823,
   input         match_out5824,
   input         match_out5825,
   input         match_out5826,
   input         match_out5827,
   input         match_out5828,
   input         match_out5829,
   input         match_out5830,
   input         match_out5831,
   input         match_out5832,
   input         match_out5833,
   input         match_out5834,
   input         match_out5835,
   input         match_out5836,
   input         match_out5837,
   input         match_out5838,
   input         match_out5839,
   input         match_out5840,
   input         match_out5841,
   input         match_out5842,
   input         match_out5843,
   input         match_out5844,
   input         match_out5845,
   input         match_out5846,
   input         match_out5847,
   input         match_out5848,
   input         match_out5849,
   input         match_out5850,
   input         match_out5851,
   input         match_out5852,
   input         match_out5853,
   input         match_out5854,
   input         match_out5855,
   input         match_out5856,
   input         match_out5857,
   input         match_out5858,
   input         match_out5859,
   input         match_out5860,
   input         match_out5861,
   input         match_out5862,
   input         match_out5863,
   input         match_out5864,
   input         match_out5865,
   input         match_out5866,
   input         match_out5867,
   input         match_out5868,
   input         match_out5869,
   input         match_out5870,
   input         match_out5871,
   input         match_out5872,
   input         match_out5873,
   input         match_out5874,
   input         match_out5875,
   input         match_out5876,
   input         match_out5877,
   input         match_out5878,
   input         match_out5879,
   input         match_out5880,
   input         match_out5881,
   input         match_out5882,
   input         match_out5883,
   input         match_out5884,
   input         match_out5885,
   input         match_out5886,
   input         match_out5887,
   input         match_out5888,
   input         match_out5889,
   input         match_out5890,
   input         match_out5891,
   input         match_out5892,
   input         match_out5893,
   input         match_out5894,
   input         match_out5895,
   input         match_out5896,
   input         match_out5897,
   input         match_out5898,
   input         match_out5899,
   input         match_out5900,
   input         match_out5901,
   input         match_out5902,
   input         match_out5903,
   input         match_out5904,
   input         match_out5905,
   input         match_out5906,
   input         match_out5907,
   input         match_out5908,
   input         match_out5909,
   input         match_out5910,
   input         match_out5911,
   input         match_out5912,
   input         match_out5913,
   input         match_out5914,
   input         match_out5915,
   input         match_out5916,
   input         match_out5917,
   input         match_out5918,
   input         match_out5919,
   input         match_out5920,
   input         match_out5921,
   input         match_out5922,
   input         match_out5923,
   input         match_out5924,
   input         match_out5925,
   input         match_out5926,
   input         match_out5927,
   input         match_out5928,
   input         match_out5929,
   input         match_out5930,
   input         match_out5931,
   input         match_out5932,
   input         match_out5933,
   input         match_out5934,
   input         match_out5935,
   input         match_out5936,
   input         match_out5937,
   input         match_out5938,
   input         match_out5939,
   input         match_out5940,
   input         match_out5941,
   input         match_out5942,
   input         match_out5943,
   input         match_out5944,
   input         match_out5945,
   input         match_out5946,
   input         match_out5947,
   input         match_out5948,
   input         match_out5949,
   input         match_out5950,
   input         match_out5951,
   input         match_out5952,
   input         match_out5953,
   input         match_out5954,
   input         match_out5955,
   input         match_out5956,
   input         match_out5957,
   input         match_out5958,
   input         match_out5959,
   input         match_out5960,
   input         match_out5961,
   input         match_out5962,
   input         match_out5963,
   input         match_out5964,
   input         match_out5965,
   input         match_out5966,
   input         match_out5967,
   input         match_out5968,
   input         match_out5969,
   input         match_out5970,
   input         match_out5971,
   input         match_out5972,
   input         match_out5973,
   input         match_out5974,
   input         match_out5975,
   input         match_out5976,
   input         match_out5977,
   input         match_out5978,
   input         match_out5979,
   input         match_out5980,
   input         match_out5981,
   input         match_out5982,
   input         match_out5983,
   input         match_out5984,
   input         match_out5985,
   input         match_out5986,
   input         match_out5987,
   input         match_out5988,
   input         match_out5989,
   input         match_out5990,
   input         match_out5991,
   input         match_out5992,
   input         match_out5993,
   input         match_out5994,
   input         match_out5995,
   input         match_out5996,
   input         match_out5997,
   input         match_out5998,
   input         match_out5999,
   input         match_out6000,
   input         match_out6001,
   input         match_out6002,
   input         match_out6003,
   input         match_out6004,
   input         match_out6005,
   input         match_out6006,
   input         match_out6007,
   input         match_out6008,
   input         match_out6009,
   input         match_out6010,
   input         match_out6011,
   input         match_out6012,
   input         match_out6013,
   input         match_out6014,
   input         match_out6015,
   input         match_out6016,
   input         match_out6017,
   input         match_out6018,
   input         match_out6019,
   input         match_out6020,
   input         match_out6021,
   input         match_out6022,
   input         match_out6023,
   input         match_out6024,
   input         match_out6025,
   input         match_out6026,
   input         match_out6027,
   input         match_out6028,
   input         match_out6029,
   input         match_out6030,
   input         match_out6031,
   input         match_out6032,
   input         match_out6033,
   input         match_out6034,
   input         match_out6035,
   input         match_out6036,
   input         match_out6037,
   input         match_out6038,
   input         match_out6039,
   input         match_out6040,
   input         match_out6041,
   input         match_out6042,
   input         match_out6043,
   input         match_out6044,
   input         match_out6045,
   input         match_out6046,
   input         match_out6047,
   input         match_out6048,
   input         match_out6049,
   input         match_out6050,
   input         match_out6051,
   input         match_out6052,
   input         match_out6053,
   input         match_out6054,
   input         match_out6055,
   input         match_out6056,
   input         match_out6057,
   input         match_out6058,
   input         match_out6059,
   input         match_out6060,
   input         match_out6061,
   input         match_out6062,
   input         match_out6063,
   input         match_out6064,
   input         match_out6065,
   input         match_out6066,
   input         match_out6067,
   input         match_out6068,
   input         match_out6069,
   input         match_out6070,
   input         match_out6071,
   input         match_out6072,
   input         match_out6073,
   input         match_out6074,
   input         match_out6075,
   input         match_out6076,
   input         match_out6077,
   input         match_out6078,
   input         match_out6079,
   input         match_out6080,
   input         match_out6081,
   input         match_out6082,
   input         match_out6083,
   input         match_out6084,
   input         match_out6085,
   input         match_out6086,
   input         match_out6087,
   input         match_out6088,
   input         match_out6089,
   input         match_out6090,
   input         match_out6091,
   input         match_out6092,
   input         match_out6093,
   input         match_out6094,
   input         match_out6095,
   input         match_out6096,
   input         match_out6097,
   input         match_out6098,
   input         match_out6099,
   input         match_out6100,
   input         match_out6101,
   input         match_out6102,
   input         match_out6103,
   input         match_out6104,
   input         match_out6105,
   input         match_out6106,
   input         match_out6107,
   input         match_out6108,
   input         match_out6109,
   input         match_out6110,
   input         match_out6111,
   input         match_out6112,
   input         match_out6113,
   input         match_out6114,
   input         match_out6115,
   input         match_out6116,
   input         match_out6117,
   input         match_out6118,
   input         match_out6119,
   input         match_out6120,
   input         match_out6121,
   input         match_out6122,
   input         match_out6123,
   input         match_out6124,
   input         match_out6125,
   input         match_out6126,
   input         match_out6127,
   input         match_out6128,
   input         match_out6129,
   input         match_out6130,
   input         match_out6131,
   input         match_out6132,
   input         match_out6133,
   input         match_out6134,
   input         match_out6135,
   input         match_out6136,
   input         match_out6137,
   input         match_out6138,
   input         match_out6139,
   input         match_out6140,
   input         match_out6141,
   input         match_out6142,
   input         match_out6143,
   input         match_out6144,
   input         match_out6145,
   input         match_out6146,
   input         match_out6147,
   input         match_out6148,
   input         match_out6149,
   input         match_out6150,
   input         match_out6151,
   input         match_out6152,
   input         match_out6153,
   input         match_out6154,
   input         match_out6155,
   input         match_out6156,
   input         match_out6157,
   input         match_out6158,
   input         match_out6159,
   input         match_out6160,
   input         match_out6161,
   input         match_out6162,
   input         match_out6163,
   input         match_out6164,
   input         match_out6165,
   input         match_out6166,
   input         match_out6167,
   input         match_out6168,
   input         match_out6169,
   input         match_out6170,
   input         match_out6171,
   input         match_out6172,
   input         match_out6173,
   input         match_out6174,
   input         match_out6175,
   input         match_out6176,
   input         match_out6177,
   input         match_out6178,
   input         match_out6179,
   input         match_out6180,
   input         match_out6181,
   input         match_out6182,
   input         match_out6183,
   input         match_out6184,
   input         match_out6185,
   input         match_out6186,
   input         match_out6187,
   input         match_out6188,
   input         match_out6189,
   input         match_out6190,
   input         match_out6191,
   input         match_out6192,
   input         match_out6193,
   input         match_out6194,
   input         match_out6195,
   input         match_out6196,
   input         match_out6197,
   input         match_out6198,
   input         match_out6199,
   input         match_out6200,
   input         match_out6201,
   input         match_out6202,
   input         match_out6203,
   input         match_out6204,
   input         match_out6205,
   input         match_out6206,
   input         match_out6207,
   input         match_out6208,
   input         match_out6209,
   input         match_out6210,
   input         match_out6211,
   input         match_out6212,
   input         match_out6213,
   input         match_out6214,
   input         match_out6215,
   input         match_out6216,
   input         match_out6217,
   input         match_out6218,
   input         match_out6219,
   input         match_out6220,
   input         match_out6221,
   input         match_out6222,
   input         match_out6223,
   input         match_out6224,
   input         match_out6225,
   input         match_out6226,
   input         match_out6227,
   input         match_out6228,
   input         match_out6229,
   input         match_out6230,
   input         match_out6231,
   input         match_out6232,
   input         match_out6233,
   input         match_out6234,
   input         match_out6235,
   input         match_out6236,
   input         match_out6237,
   input         match_out6238,
   input         match_out6239,
   input         match_out6240,
   input         match_out6241,
   input         match_out6242,
   input         match_out6243,
   input         match_out6244,
   input         match_out6245,
   input         match_out6246,
   input         match_out6247,
   input         match_out6248,
   input         match_out6249,
   input         match_out6250,
   input         match_out6251,
   input         match_out6252,
   input         match_out6253,
   input         match_out6254,
   input         match_out6255,
   input         match_out6256,
   input         match_out6257,
   input         match_out6258,
   input         match_out6259,
   input         match_out6260,
   input         match_out6261,
   input         match_out6262,
   input         match_out6263,
   input         match_out6264,
   input         match_out6265,
   input         match_out6266,
   input         match_out6267,
   input         match_out6268,
   input         match_out6269,
   input         match_out6270,
   input         match_out6271,
   input         match_out6272,
   input         match_out6273,
   input         match_out6274,
   input         match_out6275,
   input         match_out6276,
   input         match_out6277,
   input         match_out6278,
   input         match_out6279,
   input         match_out6280,
   input         match_out6281,
   input         match_out6282,
   input         match_out6283,
   input         match_out6284,
   input         match_out6285,
   input         match_out6286,
   input         match_out6287,
   input         match_out6288,
   input         match_out6289,
   input         match_out6290,
   input         match_out6291,
   input         match_out6292,
   input         match_out6293,
   input         match_out6294,
   input         match_out6295,
   input         match_out6296,
   input         match_out6297,
   input         match_out6298,
   input         match_out6299,
   input         match_out6300,
   input         match_out6301,
   input         match_out6302,
   input         match_out6303,
   input         match_out6304,
   input         match_out6305,
   input         match_out6306,
   input         match_out6307,
   input         match_out6308,
   input         match_out6309,
   input         match_out6310,
   input         match_out6311,
   input         match_out6312,
   input         match_out6313,
   input         match_out6314,
   input         match_out6315,
   input         match_out6316,
   input         match_out6317,
   input         match_out6318,
   input         match_out6319,
   input         match_out6320,
   input         match_out6321,
   input         match_out6322,
   input         match_out6323,
   input         match_out6324,
   input         match_out6325,
   input         match_out6326,
   input         match_out6327,
   input         match_out6328,
   input         match_out6329,
   input         match_out6330,
   input         match_out6331,
   input         match_out6332,
   input         match_out6333,
   input         match_out6334,
   input         match_out6335,
   input         match_out6336,
   input         match_out6337,
   input         match_out6338,
   input         match_out6339,
   input         match_out6340,
   input         match_out6341,
   input         match_out6342,
   input         match_out6343,
   input         match_out6344,
   input         match_out6345,
   input         match_out6346,
   input         match_out6347,
   input         match_out6348,
   input         match_out6349,
   input         match_out6350,
   input         match_out6351,
   input         match_out6352,
   input         match_out6353,
   input         match_out6354,
   input         match_out6355,
   input         match_out6356,
   input         match_out6357,
   input         match_out6358,
   input         match_out6359,
   input         match_out6360,
   input         match_out6361,
   input         match_out6362,
   input         match_out6363,
   input         match_out6364,
   input         match_out6365,
   input         match_out6366,
   input         match_out6367,
   input         match_out6368,
   input         match_out6369,
   input         match_out6370,
   input         match_out6371,
   input         match_out6372,
   input         match_out6373,
   input         match_out6374,
   input         match_out6375,
   input         match_out6376,
   input         match_out6377,
   input         match_out6378,
   input         match_out6379,
   input         match_out6380,
   input         match_out6381,
   input         match_out6382,
   input         match_out6383,
   input         match_out6384,
   input         match_out6385,
   input         match_out6386,
   input         match_out6387,
   input         match_out6388,
   input         match_out6389,
   input         match_out6390,
   input         match_out6391,
   input         match_out6392,
   input         match_out6393,
   input         match_out6394,
   input         match_out6395,
   input         match_out6396,
   input         match_out6397,
   input         match_out6398,
   input         match_out6399,
   input         match_out6400,
   input         match_out6401,
   input         match_out6402,
   input         match_out6403,
   input         match_out6404,
   input         match_out6405,
   input         match_out6406,
   input         match_out6407,
   input         match_out6408,
   input         match_out6409,
   input         match_out6410,
   input         match_out6411,
   input         match_out6412,
   input         match_out6413,
   input         match_out6414,
   input         match_out6415,
   input         match_out6416,
   input         match_out6417,
   input         match_out6418,
   input         match_out6419,
   input         match_out6420,
   input         match_out6421,
   input         match_out6422,
   input         match_out6423,
   input         match_out6424,
   input         match_out6425,
   input         match_out6426,
   input         match_out6427,
   input         match_out6428,
   input         match_out6429,
   input         match_out6430,
   input         match_out6431,
   input         match_out6432,
   input         match_out6433,
   input         match_out6434,
   input         match_out6435,
   input         match_out6436,
   input         match_out6437,
   input         match_out6438,
   input         match_out6439,
   input         match_out6440,
   input         match_out6441,
   input         match_out6442,
   input         match_out6443,
   input         match_out6444,
   input         match_out6445,
   input         match_out6446,
   input         match_out6447,
   input         match_out6448,
   input         match_out6449,
   input         match_out6450,
   input         match_out6451,
   input         match_out6452,
   input         match_out6453,
   input         match_out6454,
   input         match_out6455,
   input         match_out6456,
   input         match_out6457,
   input         match_out6458,
   input         match_out6459,
   input         match_out6460,
   input         match_out6461,
   input         match_out6462,
   input         match_out6463,
   input         match_out6464,
   input         match_out6465,
   input         match_out6466,
   input         match_out6467,
   input         match_out6468,
   input         match_out6469,
   input         match_out6470,
   input         match_out6471,
   input         match_out6472,
   input         match_out6473,
   input         match_out6474,
   input         match_out6475,
   input         match_out6476,
   input         match_out6477,
   input         match_out6478,
   input         match_out6479,
   input         match_out6480,
   input         match_out6481,
   input         match_out6482,
   input         match_out6483,
   input         match_out6484,
   input         match_out6485,
   input         match_out6486,
   input         match_out6487,
   input         match_out6488,
   input         match_out6489,
   input         match_out6490,
   input         match_out6491,
   input         match_out6492,
   input         match_out6493,
   input         match_out6494,
   input         match_out6495,
   input         match_out6496,
   input         match_out6497,
   input         match_out6498,
   input         match_out6499,
   input         match_out6500,
   input         match_out6501,
   input         match_out6502,
   input         match_out6503,
   input         match_out6504,
   input         match_out6505,
   input         match_out6506,
   input         match_out6507,
   input         match_out6508,
   input         match_out6509,
   input         match_out6510,
   input         match_out6511,
   input         match_out6512,
   input         match_out6513,
   input         match_out6514,
   input         match_out6515,
   input         match_out6516,
   input         match_out6517,
   input         match_out6518,
   input         match_out6519,
   input         match_out6520,
   input         match_out6521,
   input         match_out6522,
   input         match_out6523,
   input         match_out6524,
   input         match_out6525,
   input         match_out6526,
   input         match_out6527,
   input         match_out6528,
   input         match_out6529,
   input         match_out6530,
   input         match_out6531,
   input         match_out6532,
   input         match_out6533,
   input         match_out6534,
   input         match_out6535,
   input         match_out6536,
   input         match_out6537,
   input         match_out6538,
   input         match_out6539,
   input         match_out6540,
   input         match_out6541,
   input         match_out6542,
   input         match_out6543,
   input         match_out6544,
   input         match_out6545,
   input         match_out6546,
   input         match_out6547,
   input         match_out6548,
   input         match_out6549,
   input         match_out6550,
   input         match_out6551,
   input         match_out6552,
   input         match_out6553,
   input         match_out6554,
   input         match_out6555,
   input         match_out6556,
   input         match_out6557,
   input         match_out6558,
   input         match_out6559,
   input         match_out6560,
   input         match_out6561,
   input         match_out6562,
   input         match_out6563,
   input         match_out6564,
   input         match_out6565,
   input         match_out6566,
   input         match_out6567,
   input         match_out6568,
   input         match_out6569,
   input         match_out6570,
   input         match_out6571,
   input         match_out6572,
   input         match_out6573,
   input         match_out6574,
   input         match_out6575,
   input         match_out6576,
   input         match_out6577,
   input         match_out6578,
   input         match_out6579,
   input         match_out6580,
   input         match_out6581,
   input         match_out6582,
   input         match_out6583,
   input         match_out6584,
   input         match_out6585,
   input         match_out6586,
   input         match_out6587,
   input         match_out6588,
   input         match_out6589,
   input         match_out6590,
   input         match_out6591,
   input         match_out6592,
   input         match_out6593,
   input         match_out6594,
   input         match_out6595,
   input         match_out6596,
   input         match_out6597,
   input         match_out6598,
   input         match_out6599,
   input         match_out6600,
   input         match_out6601,
   input         match_out6602,
   input         match_out6603,
   input         match_out6604,
   input         match_out6605,
   input         match_out6606,
   input         match_out6607,
   input         match_out6608,
   input         match_out6609,
   input         match_out6610,
   input         match_out6611,
   input         match_out6612,
   input         match_out6613,
   input         match_out6614,
   input         match_out6615,
   input         match_out6616,
   input         match_out6617,
   input         match_out6618,
   input         match_out6619,
   input         match_out6620,
   input         match_out6621,
   input         match_out6622,
   input         match_out6623,
   input         match_out6624,
   input         match_out6625,
   input         match_out6626,
   input         match_out6627,
   input         match_out6628,
   input         match_out6629,
   input         match_out6630,
   input         match_out6631,
   input         match_out6632,
   input         match_out6633,
   input         match_out6634,
   input         match_out6635,
   input         match_out6636,
   input         match_out6637,
   input         match_out6638,
   input         match_out6639,
   input         match_out6640,
   input         match_out6641,
   input         match_out6642,
   input         match_out6643,
   input         match_out6644,
   input         match_out6645,
   input         match_out6646,
   input         match_out6647,
   input         match_out6648,
   input         match_out6649,
   input         match_out6650,
   input         match_out6651,
   input         match_out6652,
   input         match_out6653,
   input         match_out6654,
   input         match_out6655,
   input         match_out6656,
   input         match_out6657,
   input         match_out6658,
   input         match_out6659,
   input         match_out6660,
   input         match_out6661,
   input         match_out6662,
   input         match_out6663,
   input         match_out6664,
   input         match_out6665,
   input         match_out6666,
   input         match_out6667,
   input         match_out6668,
   input         match_out6669,
   input         match_out6670,
   input         match_out6671,
   input         match_out6672,
   input         match_out6673,
   input         match_out6674,
   input         match_out6675,
   input         match_out6676,
   input         match_out6677,
   input         match_out6678,
   input         match_out6679,
   input         match_out6680,
   input         match_out6681,
   input         match_out6682,
   input         match_out6683,
   input         match_out6684,
   input         match_out6685,
   input         match_out6686,
   input         match_out6687,
   input         match_out6688,
   input         match_out6689,
   input         match_out6690,
   input         match_out6691,
   input         match_out6692,
   input         match_out6693,
   input         match_out6694,
   input         match_out6695,
   input         match_out6696,
   input         match_out6697,
   input         match_out6698,
   input         match_out6699,
   input         match_out6700,
   input         match_out6701,
   input         match_out6702,
   input         match_out6703,
   input         match_out6704,
   input         match_out6705,
   input         match_out6706,
   input         match_out6707,
   input         match_out6708,
   input         match_out6709,
   input         match_out6710,
   input         match_out6711,
   input         match_out6712,
   input         match_out6713,
   input         match_out6714,
   input         match_out6715,
   input         match_out6716,
   input         match_out6717,
   input         match_out6718,
   input         match_out6719,
   input         match_out6720,
   input         match_out6721,
   input         match_out6722,
   input         match_out6723,
   input         match_out6724,
   input         match_out6725,
   input         match_out6726,
   input         match_out6727,
   input         match_out6728,
   input         match_out6729,
   input         match_out6730,
   input         match_out6731,
   input         match_out6732,
   input         match_out6733,
   input         match_out6734,
   input         match_out6735,
   input         match_out6736,
   input         match_out6737,
   input         match_out6738,
   input         match_out6739,
   input         match_out6740,
   input         match_out6741,
   input         match_out6742,
   input         match_out6743,
   input         match_out6744,
   input         match_out6745,
   input         match_out6746,
   input         match_out6747,
   input         match_out6748,
   input         match_out6749,
   input         match_out6750,
   input         match_out6751,
   input         match_out6752,
   input         match_out6753,
   input         match_out6754,
   input         match_out6755,
   input         match_out6756,
   input         match_out6757,
   input         match_out6758,
   input         match_out6759,
   input         match_out6760,
   input         match_out6761,
   input         match_out6762,
   input         match_out6763,
   input         match_out6764,
   input         match_out6765,
   input         match_out6766,
   input         match_out6767,
   input         match_out6768,
   input         match_out6769,
   input         match_out6770,
   input         match_out6771,
   input         match_out6772,
   input         match_out6773,
   input         match_out6774,
   input         match_out6775,
   input         match_out6776,
   input         match_out6777,
   input         match_out6778,
   input         match_out6779,
   input         match_out6780,
   input         match_out6781,
   input         match_out6782,
   input         match_out6783,
   input         match_out6784,
   input         match_out6785,
   input         match_out6786,
   input         match_out6787,
   input         match_out6788,
   input         match_out6789,
   input         match_out6790,
   input         match_out6791,
   input         match_out6792,
   input         match_out6793,
   input         match_out6794,
   input         match_out6795,
   input         match_out6796,
   input         match_out6797,
   input         match_out6798,
   input         match_out6799,
   input         match_out6800,
   input         match_out6801,
   input         match_out6802,
   input         match_out6803,
   input         match_out6804,
   input         match_out6805,
   input         match_out6806,
   input         match_out6807,
   input         match_out6808,
   input         match_out6809,
   input         match_out6810,
   input         match_out6811,
   input         match_out6812,
   input         match_out6813,
   input         match_out6814,
   input         match_out6815,
   input         match_out6816,
   input         match_out6817,
   input         match_out6818,
   input         match_out6819,
   input         match_out6820,
   input         match_out6821,
   input         match_out6822,
   input         match_out6823,
   input         match_out6824,
   input         match_out6825,
   input         match_out6826,
   input         match_out6827,
   input         match_out6828,
   input         match_out6829,
   input         match_out6830,
   input         match_out6831,
   input         match_out6832,
   input         match_out6833,
   input         match_out6834,
   input         match_out6835,
   input         match_out6836,
   input         match_out6837,
   input         match_out6838,
   input         match_out6839,
   input         match_out6840,
   input         match_out6841,
   input         match_out6842,
   input         match_out6843,
   input         match_out6844,
   input         match_out6845,
   input         match_out6846,
   input         match_out6847,
   input         match_out6848,
   input         match_out6849,
   input         match_out6850,
   input         match_out6851,
   input         match_out6852,
   input         match_out6853,
   input         match_out6854,
   input         match_out6855,
   input         match_out6856,
   input         match_out6857,
   input         match_out6858,
   input         match_out6859,
   input         match_out6860,
   input         match_out6861,
   input         match_out6862,
   input         match_out6863,
   input         match_out6864,
   input         match_out6865,
   input         match_out6866,
   input         match_out6867,
   input         match_out6868,
   input         match_out6869,
   input         match_out6870,
   input         match_out6871,
   input         match_out6872,
   input         match_out6873,
   input         match_out6874,
   input         match_out6875,
   input         match_out6876,
   input         match_out6877,
   input         match_out6878,
   input         match_out6879,
   input         match_out6880,
   input         match_out6881,
   input         match_out6882,
   input         match_out6883,
   input         match_out6884,
   input         match_out6885,
   input         match_out6886,
   input         match_out6887,
   input         match_out6888,
   input         match_out6889,
   input         match_out6890,
   input         match_out6891,
   input         match_out6892,
   input         match_out6893,
   input         match_out6894,
   input         match_out6895,
   input         match_out6896,
   input         match_out6897,
   input         match_out6898,
   input         match_out6899,
   input         match_out6900,
   input         match_out6901,
   input         match_out6902,
   input         match_out6903,
   input         match_out6904,
   input         match_out6905,
   input         match_out6906,
   input         match_out6907,
   input         match_out6908,
   input         match_out6909,
   input         match_out6910,
   input         match_out6911,
   input         match_out6912,
   input         match_out6913,
   input         match_out6914,
   input         match_out6915,
   input         match_out6916,
   input         match_out6917,
   input         match_out6918,
   input         match_out6919,
   input         match_out6920,
   input         match_out6921,
   input         match_out6922,
   input         match_out6923,
   input         match_out6924,
   input         match_out6925,
   input         match_out6926,
   input         match_out6927,
   input         match_out6928,
   input         match_out6929,
   input         match_out6930,
   input         match_out6931,
   input         match_out6932,
   input         match_out6933,
   input         match_out6934,
   input         match_out6935,
   input         match_out6936,
   input         match_out6937,
   input         match_out6938,
   input         match_out6939,
   input         match_out6940,
   input         match_out6941,
   input         match_out6942,
   input         match_out6943,
   input         match_out6944,
   input         match_out6945,
   input         match_out6946,
   input         match_out6947,
   input         match_out6948,
   input         match_out6949,
   input         match_out6950,
   input         match_out6951,
   input         match_out6952,
   input         match_out6953,
   input         match_out6954,
   input         match_out6955,
   input         match_out6956,
   input         match_out6957,
   input         match_out6958,
   input         match_out6959,
   input         match_out6960,
   input         match_out6961,
   input         match_out6962,
   input         match_out6963,
   input         match_out6964,
   input         match_out6965,
   input         match_out6966,
   input         match_out6967,
   input         match_out6968,
   input         match_out6969,
   input         match_out6970,
   input         match_out6971,
   input         match_out6972,
   input         match_out6973,
   input         match_out6974,
   input         match_out6975,
   input         match_out6976,
   input         match_out6977,
   input         match_out6978,
   input         match_out6979,
   input         match_out6980,
   input         match_out6981,
   input         match_out6982,
   input         match_out6983,
   input         match_out6984,
   input         match_out6985,
   input         match_out6986,
   input         match_out6987,
   input         match_out6988,
   input         match_out6989,
   input         match_out6990,
   input         match_out6991,
   input         match_out6992,
   input         match_out6993,
   input         match_out6994,
   input         match_out6995,
   input         match_out6996,
   input         match_out6997,
   input         match_out6998,
   input         match_out6999,
   input         match_out7000,
   input         match_out7001,
   input         match_out7002,
   input         match_out7003,
   input         match_out7004,
   input         match_out7005,
   input         match_out7006,
   input         match_out7007,
   input         match_out7008,
   input         match_out7009,
   input         match_out7010,
   input         match_out7011,
   input         match_out7012,
   input         match_out7013,
   input         match_out7014,
   input         match_out7015,
   input         match_out7016,
   input         match_out7017,
   input         match_out7018,
   input         match_out7019,
   input         match_out7020,
   input         match_out7021,
   input         match_out7022,
   input         match_out7023,
   input         match_out7024,
   input         match_out7025,
   input         match_out7026,
   input         match_out7027,
   input         match_out7028,
   input         match_out7029,
   input         match_out7030,
   input         match_out7031,
   input         match_out7032,
   input         match_out7033,
   input         match_out7034,
   input         match_out7035,
   input         match_out7036,
   input         match_out7037,
   input         match_out7038,
   input         match_out7039,
   input         match_out7040,
   input         match_out7041,
   input         match_out7042,
   input         match_out7043,
   input         match_out7044,
   input         match_out7045,
   input         match_out7046,
   input         match_out7047,
   input         match_out7048,
   input         match_out7049,
   input         match_out7050,
   input         match_out7051,
   input         match_out7052,
   input         match_out7053,
   input         match_out7054,
   input         match_out7055,
   input         match_out7056,
   input         match_out7057,
   input         match_out7058,
   input         match_out7059,
   input         match_out7060,
   input         match_out7061,
   input         match_out7062,
   input         match_out7063,
   input         match_out7064,
   input         match_out7065,
   input         match_out7066,
   input         match_out7067,
   input         match_out7068,
   input         match_out7069,
   input         match_out7070,
   input         match_out7071,
   input         match_out7072,
   input         match_out7073,
   input         match_out7074,
   input         match_out7075,
   input         match_out7076,
   input         match_out7077,
   input         match_out7078,
   input         match_out7079,
   input         match_out7080,
   input         match_out7081,
   input         match_out7082,
   input         match_out7083,
   input         match_out7084,
   input         match_out7085,
   input         match_out7086,
   input         match_out7087,
   input         match_out7088,
   input         match_out7089,
   input         match_out7090,
   input         match_out7091,
   input         match_out7092,
   input         match_out7093,
   input         match_out7094,
   input         match_out7095,
   input         match_out7096,
   input         match_out7097,
   input         match_out7098,
   input         match_out7099,
   input         match_out7100,
   input         match_out7101,
   input         match_out7102,
   input         match_out7103,
   input         match_out7104,
   input         match_out7105,
   input         match_out7106,
   input         match_out7107,
   input         match_out7108,
   input         match_out7109,
   input         match_out7110,
   input         match_out7111,
   input         match_out7112,
   input         match_out7113,
   input         match_out7114,
   input         match_out7115,
   input         match_out7116,
   input         match_out7117,
   input         match_out7118,
   input         match_out7119,
   input         match_out7120,
   input         match_out7121,
   input         match_out7122,
   input         match_out7123,
   input         match_out7124,
   input         match_out7125,
   input         match_out7126,
   input         match_out7127,
   input         match_out7128,
   input         match_out7129,
   input         match_out7130,
   input         match_out7131,
   input         match_out7132,
   input         match_out7133,
   input         match_out7134,
   input         match_out7135,
   input         match_out7136,
   input         match_out7137,
   input         match_out7138,
   input         match_out7139,
   input         match_out7140,
   input         match_out7141,
   input         match_out7142,
   input         match_out7143,
   input         match_out7144,
   input         match_out7145,
   input         match_out7146,
   input         match_out7147,
   input         match_out7148,
   input         match_out7149,
   input         match_out7150,
   input         match_out7151,
   input         match_out7152,
   input         match_out7153,
   input         match_out7154,
   input         match_out7155,
   input         match_out7156,
   input         match_out7157,
   input         match_out7158,
   input         match_out7159,
   input         match_out7160,
   input         match_out7161,
   input         match_out7162,
   input         match_out7163,
   input         match_out7164,
   input         match_out7165,
   input         match_out7166,
   input         match_out7167,
   input         match_out7168,
   input         match_out7169,
   input         match_out7170,
   input         match_out7171,
   input         match_out7172,
   input         match_out7173,
   input         match_out7174,
   input         match_out7175,
   input         match_out7176,
   input         match_out7177,
   input         match_out7178,
   input         match_out7179,
   input         match_out7180,
   input         match_out7181,
   input         match_out7182,
   input         match_out7183,
   input         match_out7184,
   input         match_out7185,
   input         match_out7186,
   input         match_out7187,
   input         match_out7188,
   input         match_out7189,
   input         match_out7190,
   input         match_out7191,
   input         match_out7192,
   input         match_out7193,
   input         match_out7194,
   input         match_out7195,
   input         match_out7196,
   input         match_out7197,
   input         match_out7198,
   input         match_out7199,
   input         match_out7200,
   input         match_out7201,
   input         match_out7202,
   input         match_out7203,
   input         match_out7204,
   input         match_out7205,
   input         match_out7206,
   input         match_out7207,
   input         match_out7208,
   input         match_out7209,
   input         match_out7210,
   input         match_out7211,
   input         match_out7212,
   input         match_out7213,
   input         match_out7214,
   input         match_out7215,
   input         match_out7216,
   input         match_out7217,
   input         match_out7218,
   input         match_out7219,
   input         match_out7220,
   input         match_out7221,
   input         match_out7222,
   input         match_out7223,
   input         match_out7224,
   input         match_out7225,
   input         match_out7226,
   input         match_out7227,
   input         match_out7228,
   input         match_out7229,
   input         match_out7230,
   input         match_out7231,
   input         match_out7232,
   input         match_out7233,
   input         match_out7234,
   input         match_out7235,
   input         match_out7236,
   input         match_out7237,
   input         match_out7238,
   input         match_out7239,
   input         match_out7240,
   input         match_out7241,
   input         match_out7242,
   input         match_out7243,
   input         match_out7244,
   input         match_out7245,
   input         match_out7246,
   input         match_out7247,
   input         match_out7248,
   input         match_out7249,
   input         match_out7250,
   input         match_out7251,
   input         match_out7252,
   input         match_out7253,
   input         match_out7254,
   input         match_out7255,
   input         match_out7256,
   input         match_out7257,
   input         match_out7258,
   input         match_out7259,
   input         match_out7260,
   input         match_out7261,
   input         match_out7262,
   input         match_out7263,
   input         match_out7264,
   input         match_out7265,
   input         match_out7266,
   input         match_out7267,
   input         match_out7268,
   input         match_out7269,
   input         match_out7270,
   input         match_out7271,
   input         match_out7272,
   input         match_out7273,
   input         match_out7274,
   input         match_out7275,
   input         match_out7276,
   input         match_out7277,
   input         match_out7278,
   input         match_out7279,
   input         match_out7280,
   input         match_out7281,
   input         match_out7282,
   input         match_out7283,
   input         match_out7284,
   input         match_out7285,
   input         match_out7286,
   input         match_out7287,
   input         match_out7288,
   input         match_out7289,
   input         match_out7290,
   input         match_out7291,
   input         match_out7292,
   input         match_out7293,
   input         match_out7294,
   input         match_out7295,
   input         match_out7296,
   input         match_out7297,
   input         match_out7298,
   input         match_out7299,
   input         match_out7300,
   input         match_out7301,
   input         match_out7302,
   input         match_out7303,
   input         match_out7304,
   input         match_out7305,
   input         match_out7306,
   input         match_out7307,
   input         match_out7308,
   input         match_out7309,
   input         match_out7310,
   input         match_out7311,
   input         match_out7312,
   input         match_out7313,
   input         match_out7314,
   input         match_out7315,
   input         match_out7316,
   input         match_out7317,
   input         match_out7318,
   input         match_out7319,
   input         match_out7320,
   input         match_out7321,
   input         match_out7322,
   input         match_out7323,
   input         match_out7324,
   input         match_out7325,
   input         match_out7326,
   input         match_out7327,
   input         match_out7328,
   input         match_out7329,
   input         match_out7330,
   input         match_out7331,
   input         match_out7332,
   input         match_out7333,
   input         match_out7334,
   input         match_out7335,
   input         match_out7336,
   input         match_out7337,
   input         match_out7338,
   input         match_out7339,
   input         match_out7340,
   input         match_out7341,
   input         match_out7342,
   input         match_out7343,
   input         match_out7344,
   input         match_out7345,
   input         match_out7346,
   input         match_out7347,
   input         match_out7348,
   input         match_out7349,
   input         match_out7350,
   input         match_out7351,
   input         match_out7352,
   input         match_out7353,
   input         match_out7354,
   input         match_out7355,
   input         match_out7356,
   input         match_out7357,
   input         match_out7358,
   input         match_out7359,
   input         match_out7360,
   input         match_out7361,
   input         match_out7362,
   input         match_out7363,
   input         match_out7364,
   input         match_out7365,
   input         match_out7366,
   input         match_out7367,
   input         match_out7368,
   input         match_out7369,
   input         match_out7370,
   input         match_out7371,
   input         match_out7372,
   input         match_out7373,
   input         match_out7374,
   input         match_out7375,
   input         match_out7376,
   input         match_out7377,
   input         match_out7378,
   input         match_out7379,
   input         match_out7380,
   input         match_out7381,
   input         match_out7382,
   input         match_out7383,
   input         match_out7384,
   input         match_out7385,
   input         match_out7386,
   input         match_out7387,
   input         match_out7388,
   input         match_out7389,
   input         match_out7390,
   input         match_out7391,
   input         match_out7392,
   input         match_out7393,
   input         match_out7394,
   input         match_out7395,
   input         match_out7396,
   input         match_out7397,
   input         match_out7398,
   input         match_out7399,
   input         match_out7400,
   input         match_out7401,
   input         match_out7402,
   input         match_out7403,
   input         match_out7404,
   input         match_out7405,
   input         match_out7406,
   input         match_out7407,
   input         match_out7408,
   input         match_out7409,
   input         match_out7410,
   input         match_out7411,
   input         match_out7412,
   input         match_out7413,
   input         match_out7414,
   input         match_out7415,
   input         match_out7416,
   input         match_out7417,
   input         match_out7418,
   input         match_out7419,
   input         match_out7420,
   input         match_out7421,
   input         match_out7422,
   input         match_out7423,
   input         match_out7424,
   input         match_out7425,
   input         match_out7426,
   input         match_out7427,
   input         match_out7428,
   input         match_out7429,
   input         match_out7430,
   input         match_out7431,
   input         match_out7432,
   input         match_out7433,
   input         match_out7434,
   input         match_out7435,
   input         match_out7436,
   input         match_out7437,
   input         match_out7438,
   input         match_out7439,
   input         match_out7440,
   input         match_out7441,
   input         match_out7442,
   input         match_out7443,
   input         match_out7444,
   input         match_out7445,
   input         match_out7446,
   input         match_out7447,
   input         match_out7448,
   input         match_out7449,
   input         match_out7450,
   input         match_out7451,
   input         match_out7452,
   input         match_out7453,
   input         match_out7454,
   input         match_out7455,
   input         match_out7456,
   input         match_out7457,
   input         match_out7458,
   input         match_out7459,
   input         match_out7460,
   input         match_out7461,
   input         match_out7462,
   input         match_out7463,
   input         match_out7464,
   input         match_out7465,
   input         match_out7466,
   input         match_out7467,
   input         match_out7468,
   input         match_out7469,
   input         match_out7470,
   input         match_out7471,
   input         match_out7472,
   input         match_out7473,
   input         match_out7474,
   input         match_out7475,
   input         match_out7476,
   input         match_out7477,
   input         match_out7478,
   input         match_out7479,
   input         match_out7480,
   input         match_out7481,
   input         match_out7482,
   input         match_out7483,
   input         match_out7484,
   input         match_out7485,
   input         match_out7486,
   input         match_out7487,
   input         match_out7488,
   input         match_out7489,
   input         match_out7490,
   input         match_out7491,
   input         match_out7492,
   input         match_out7493,
   input         match_out7494,
   input         match_out7495,
   input         match_out7496,
   input         match_out7497,
   input         match_out7498,
   input         match_out7499,
   input         match_out7500,
   input         match_out7501,
   input         match_out7502,
   input         match_out7503,
   input         match_out7504,
   input         match_out7505,
   input         match_out7506,
   input         match_out7507,
   input         match_out7508,
   input         match_out7509,
   input         match_out7510,
   input         match_out7511,
   input         match_out7512,
   input         match_out7513,
   input         match_out7514,
   input         match_out7515,
   input         match_out7516,
   input         match_out7517,
   input         match_out7518,
   input         match_out7519,
   input         match_out7520,
   input         match_out7521,
   input         match_out7522,
   input         match_out7523,
   input         match_out7524,
   input         match_out7525,
   input         match_out7526,
   input         match_out7527,
   input         match_out7528,
   input         match_out7529,
   input         match_out7530,
   input         match_out7531,
   input         match_out7532,
   input         match_out7533,
   input         match_out7534,
   input         match_out7535,
   input         match_out7536,
   input         match_out7537,
   input         match_out7538,
   input         match_out7539,
   input         match_out7540,
   input         match_out7541,
   input         match_out7542,
   input         match_out7543,
   input         match_out7544,
   input         match_out7545,
   input         match_out7546,
   input         match_out7547,
   input         match_out7548,
   input         match_out7549,
   input         match_out7550,
   input         match_out7551,
   input         match_out7552,
   input         match_out7553,
   input         match_out7554,
   input         match_out7555,
   input         match_out7556,
   input         match_out7557,
   input         match_out7558,
   input         match_out7559,
   input         match_out7560,
   input         match_out7561,
   input         match_out7562,
   input         match_out7563,
   input         match_out7564,
   input         match_out7565,
   input         match_out7566,
   input         match_out7567,
   input         match_out7568,
   input         match_out7569,
   input         match_out7570,
   input         match_out7571,
   input         match_out7572,
   input         match_out7573,
   input         match_out7574,
   input         match_out7575,
   input         match_out7576,
   input         match_out7577,
   input         match_out7578,
   input         match_out7579,
   input         match_out7580,
   input         match_out7581,
   input         match_out7582,
   input         match_out7583,
   input         match_out7584,
   input         match_out7585,
   input         match_out7586,
   input         match_out7587,
   input         match_out7588,
   input         match_out7589,
   input         match_out7590,
   input         match_out7591,
   input         match_out7592,
   input         match_out7593,
   input         match_out7594,
   input         match_out7595,
   input         match_out7596,
   input         match_out7597,
   input         match_out7598,
   input         match_out7599,
   input         match_out7600,
   input         match_out7601,
   input         match_out7602,
   input         match_out7603,
   input         match_out7604,
   input         match_out7605,
   input         match_out7606,
   input         match_out7607,
   input         match_out7608,
   input         match_out7609,
   input         match_out7610,
   input         match_out7611,
   input         match_out7612,
   input         match_out7613,
   input         match_out7614,
   input         match_out7615,
   input         match_out7616,
   input         match_out7617,
   input         match_out7618,
   input         match_out7619,
   input         match_out7620,
   input         match_out7621,
   input         match_out7622,
   input         match_out7623,
   input         match_out7624,
   input         match_out7625,
   input         match_out7626,
   input         match_out7627,
   input         match_out7628,
   input         match_out7629,
   input         match_out7630,
   input         match_out7631,
   input         match_out7632,
   input         match_out7633,
   input         match_out7634,
   input         match_out7635,
   input         match_out7636,
   input         match_out7637,
   input         match_out7638,
   input         match_out7639,
   input         match_out7640,
   input         match_out7641,
   input         match_out7642,
   input         match_out7643,
   input         match_out7644,
   input         match_out7645,
   input         match_out7646,
   input         match_out7647,
   input         match_out7648,
   input         match_out7649,
   input         match_out7650,
   input         match_out7651,
   input         match_out7652,
   input         match_out7653,
   input         match_out7654,
   input         match_out7655,
   input         match_out7656,
   input         match_out7657,
   input         match_out7658,
   input         match_out7659,
   input         match_out7660,
   input         match_out7661,
   input         match_out7662,
   input         match_out7663,
   input         match_out7664,
   input         match_out7665,
   input         match_out7666,
   input         match_out7667,
   input         match_out7668,
   input         match_out7669,
   input         match_out7670,
   input         match_out7671,
   input         match_out7672,
   input         match_out7673,
   input         match_out7674,
   input         match_out7675,
   input         match_out7676,
   input         match_out7677,
   input         match_out7678,
   input         match_out7679,
   input         match_out7680,
   input         match_out7681,
   input         match_out7682,
   input         match_out7683,
   input         match_out7684,
   input         match_out7685,
   input         match_out7686,
   input         match_out7687,
   input         match_out7688,
   input         match_out7689,
   input         match_out7690,
   input         match_out7691,
   input         match_out7692,
   input         match_out7693,
   input         match_out7694,
   input         match_out7695,
   input         match_out7696,
   input         match_out7697,
   input         match_out7698,
   input         match_out7699,
   input         match_out7700,
   input         match_out7701,
   input         match_out7702,
   input         match_out7703,
   input         match_out7704,
   input         match_out7705,
   input         match_out7706,
   input         match_out7707,
   input         match_out7708,
   input         match_out7709,
   input         match_out7710,
   input         match_out7711,
   input         match_out7712,
   input         match_out7713,
   input         match_out7714,
   input         match_out7715,
   input         match_out7716,
   input         match_out7717,
   input         match_out7718,
   input         match_out7719,
   input         match_out7720,
   input         match_out7721,
   input         match_out7722,
   input         match_out7723,
   input         match_out7724,
   input         match_out7725,
   input         match_out7726,
   input         match_out7727,
   input         match_out7728,
   input         match_out7729,
   input         match_out7730,
   input         match_out7731,
   input         match_out7732,
   input         match_out7733,
   input         match_out7734,
   input         match_out7735,
   input         match_out7736,
   input         match_out7737,
   input         match_out7738,
   input         match_out7739,
   input         match_out7740,
   input         match_out7741,
   input         match_out7742,
   input         match_out7743,
   input         match_out7744,
   input         match_out7745,
   input         match_out7746,
   input         match_out7747,
   input         match_out7748,
   input         match_out7749,
   input         match_out7750,
   input         match_out7751,
   input         match_out7752,
   input         match_out7753,
   input         match_out7754,
   input         match_out7755,
   input         match_out7756,
   input         match_out7757,
   input         match_out7758,
   input         match_out7759,
   input         match_out7760,
   input         match_out7761,
   input         match_out7762,
   input         match_out7763,
   input         match_out7764,
   input         match_out7765,
   input         match_out7766,
   input         match_out7767,
   input         match_out7768,
   input         match_out7769,
   input         match_out7770,
   input         match_out7771,
   input         match_out7772,
   input         match_out7773,
   input         match_out7774,
   input         match_out7775,
   input         match_out7776,
   input         match_out7777,
   input         match_out7778,
   input         match_out7779,
   input         match_out7780,
   input         match_out7781,
   input         match_out7782,
   input         match_out7783,
   input         match_out7784,
   input         match_out7785,
   input         match_out7786,
   input         match_out7787,
   input         match_out7788,
   input         match_out7789,
   input         match_out7790,
   input         match_out7791,
   input         match_out7792,
   input         match_out7793,
   input         match_out7794,
   input         match_out7795,
   input         match_out7796,
   input         match_out7797,
   input         match_out7798,
   input         match_out7799,
   input         match_out7800,
   input         match_out7801,
   input         match_out7802,
   input         match_out7803,
   input         match_out7804,
   input         match_out7805,
   input         match_out7806,
   input         match_out7807,
   input         match_out7808,
   input         match_out7809,
   input         match_out7810,
   input         match_out7811,
   input         match_out7812,
   input         match_out7813,
   input         match_out7814,
   input         match_out7815,
   input         match_out7816,
   input         match_out7817,
   input         match_out7818,
   input         match_out7819,
   input         match_out7820,
   input         match_out7821,
   input         match_out7822,
   input         match_out7823,
   input         match_out7824,
   input         match_out7825,
   input         match_out7826,
   input         match_out7827,
   input         match_out7828,
   input         match_out7829,
   input         match_out7830,
   input         match_out7831,
   input         match_out7832,
   input         match_out7833,
   input         match_out7834,
   input         match_out7835,
   input         match_out7836,
   input         match_out7837,
   input         match_out7838,
   input         match_out7839,
   input         match_out7840,
   input         match_out7841,
   input         match_out7842,
   input         match_out7843,
   input         match_out7844,
   input         match_out7845,
   input         match_out7846,
   input         match_out7847,
   input         match_out7848,
   input         match_out7849,
   input         match_out7850,
   input         match_out7851,
   input         match_out7852,
   input         match_out7853,
   input         match_out7854,
   input         match_out7855,
   input         match_out7856,
   input         match_out7857,
   input         match_out7858,
   input         match_out7859,
   input         match_out7860,
   input         match_out7861,
   input         match_out7862,
   input         match_out7863,
   input         match_out7864,
   input         match_out7865,
   input         match_out7866,
   input         match_out7867,
   input         match_out7868,
   input         match_out7869,
   input         match_out7870,
   input         match_out7871,
   input         match_out7872,
   input         match_out7873,
   input         match_out7874,
   input         match_out7875,
   input         match_out7876,
   input         match_out7877,
   input         match_out7878,
   input         match_out7879,
   input         match_out7880,
   input         match_out7881,
   input         match_out7882,
   input         match_out7883,
   input         match_out7884,
   input         match_out7885,
   input         match_out7886,
   input         match_out7887,
   input         match_out7888,
   input         match_out7889,
   input         match_out7890,
   input         match_out7891,
   input         match_out7892,
   input         match_out7893,
   input         match_out7894,
   input         match_out7895,
   input         match_out7896,
   input         match_out7897,
   input         match_out7898,
   input         match_out7899,
   input         match_out7900,
   input         match_out7901,
   input         match_out7902,
   input         match_out7903,
   input         match_out7904,
   input         match_out7905,
   input         match_out7906,
   input         match_out7907,
   input         match_out7908,
   input         match_out7909,
   input         match_out7910,
   input         match_out7911,
   input         match_out7912,
   input         match_out7913,
   input         match_out7914,
   input         match_out7915,
   input         match_out7916,
   input         match_out7917,
   input         match_out7918,
   input         match_out7919,
   input         match_out7920,
   input         match_out7921,
   input         match_out7922,
   input         match_out7923,
   input         match_out7924,
   input         match_out7925,
   input         match_out7926,
   input         match_out7927,
   input         match_out7928,
   input         match_out7929,
   input         match_out7930,
   input         match_out7931,
   input         match_out7932,
   input         match_out7933,
   input         match_out7934,
   input         match_out7935,
   input         match_out7936,
   input         match_out7937,
   input         match_out7938,
   input         match_out7939,
   input         match_out7940,
   input         match_out7941,
   input         match_out7942,
   input         match_out7943,
   input         match_out7944,
   input         match_out7945,
   input         match_out7946,
   input         match_out7947,
   input         match_out7948,
   input         match_out7949,
   input         match_out7950,
   input         match_out7951,
   input         match_out7952,
   input         match_out7953,
   input         match_out7954,
   input         match_out7955,
   input         match_out7956,
   input         match_out7957,
   input         match_out7958,
   input         match_out7959,
   input         match_out7960,
   input         match_out7961,
   input         match_out7962,
   input         match_out7963,
   input         match_out7964,
   input         match_out7965,
   input         match_out7966,
   input         match_out7967,
   input         match_out7968,
   input         match_out7969,
   input         match_out7970,
   input         match_out7971,
   input         match_out7972,
   input         match_out7973,
   input         match_out7974,
   input         match_out7975,
   input         match_out7976,
   input         match_out7977,
   input         match_out7978,
   input         match_out7979,
   input         match_out7980,
   input         match_out7981,
   input         match_out7982,
   input         match_out7983,
   input         match_out7984,
   input         match_out7985,
   input         match_out7986,
   input         match_out7987,
   input         match_out7988,
   input         match_out7989,
   input         match_out7990,
   input         match_out7991,
   input         match_out7992,
   input         match_out7993,
   input         match_out7994,
   input         match_out7995,
   input         match_out7996,
   input         match_out7997,
   input         match_out7998,
   input         match_out7999,
   input         match_out8000,
   input         match_out8001,
   input         match_out8002,
   input         match_out8003,
   input         match_out8004,
   input         match_out8005,
   input         match_out8006,
   input         match_out8007,
   input         match_out8008,
   input         match_out8009,
   input         match_out8010,
   input         match_out8011,
   input         match_out8012,
   input         match_out8013,
   input         match_out8014,
   input         match_out8015,
   input         match_out8016,
   input         match_out8017,
   input         match_out8018,
   input         match_out8019,
   input         match_out8020,
   input         match_out8021,
   input         match_out8022,
   input         match_out8023,
   input         match_out8024,
   input         match_out8025,
   input         match_out8026,
   input         match_out8027,
   input         match_out8028,
   input         match_out8029,
   input         match_out8030,
   input         match_out8031,
   input         match_out8032,
   input         match_out8033,
   input         match_out8034,
   input         match_out8035,
   input         match_out8036,
   input         match_out8037,
   input         match_out8038,
   input         match_out8039,
   input         match_out8040,
   input         match_out8041,
   input         match_out8042,
   input         match_out8043,
   input         match_out8044,
   input         match_out8045,
   input         match_out8046,
   input         match_out8047,
   input         match_out8048,
   input         match_out8049,
   input         match_out8050,
   input         match_out8051,
   input         match_out8052,
   input         match_out8053,
   input         match_out8054,
   input         match_out8055,
   input         match_out8056,
   input         match_out8057,
   input         match_out8058,
   input         match_out8059,
   input         match_out8060,
   input         match_out8061,
   input         match_out8062,
   input         match_out8063,
   input         match_out8064,
   input         match_out8065,
   input         match_out8066,
   input         match_out8067,
   input         match_out8068,
   input         match_out8069,
   input         match_out8070,
   input         match_out8071,
   input         match_out8072,
   input         match_out8073,
   input         match_out8074,
   input         match_out8075,
   input         match_out8076,
   input         match_out8077,
   input         match_out8078,
   input         match_out8079,
   input         match_out8080,
   input         match_out8081,
   input         match_out8082,
   input         match_out8083,
   input         match_out8084,
   input         match_out8085,
   input         match_out8086,
   input         match_out8087,
   input         match_out8088,
   input         match_out8089,
   input         match_out8090,
   input         match_out8091,
   input         match_out8092,
   input         match_out8093,
   input         match_out8094,
   input         match_out8095,
   input         match_out8096,
   input         match_out8097,
   input         match_out8098,
   input         match_out8099,
   input         match_out8100,
   input         match_out8101,
   input         match_out8102,
   input         match_out8103,
   input         match_out8104,
   input         match_out8105,
   input         match_out8106,
   input         match_out8107,
   input         match_out8108,
   input         match_out8109,
   input         match_out8110,
   input         match_out8111,
   input         match_out8112,
   input         match_out8113,
   input         match_out8114,
   input         match_out8115,
   input         match_out8116,
   input         match_out8117,
   input         match_out8118,
   input         match_out8119,
   input         match_out8120,
   input         match_out8121,
   input         match_out8122,
   input         match_out8123,
   input         match_out8124,
   input         match_out8125,
   input         match_out8126,
   input         match_out8127,
   input         match_out8128,
   input         match_out8129,
   input         match_out8130,
   input         match_out8131,
   input         match_out8132,
   input         match_out8133,
   input         match_out8134,
   input         match_out8135,
   input         match_out8136,
   input         match_out8137,
   input         match_out8138,
   input         match_out8139,
   input         match_out8140,
   input         match_out8141,
   input         match_out8142,
   input         match_out8143,
   input         match_out8144,
   input         match_out8145,
   input         match_out8146,
   input         match_out8147,
   input         match_out8148,
   input         match_out8149,
   input         match_out8150,
   input         match_out8151,
   input         match_out8152,
   input         match_out8153,
   input         match_out8154,
   input         match_out8155,
   input         match_out8156,
   input         match_out8157,
   input         match_out8158,
   input         match_out8159,
   input         match_out8160,
   input         match_out8161,
   input         match_out8162,
   input         match_out8163,
   input         match_out8164,
   input         match_out8165,
   input         match_out8166,
   input         match_out8167,
   input         match_out8168,
   input         match_out8169,
   input         match_out8170,
   input         match_out8171,
   input         match_out8172,
   input         match_out8173,
   input         match_out8174,
   input         match_out8175,
   input         match_out8176,
   input         match_out8177,
   input         match_out8178,
   input         match_out8179,
   input         match_out8180,
   input         match_out8181,
   input         match_out8182,
   input         match_out8183,
   input         match_out8184,
   input         match_out8185,
   input         match_out8186,
   input         match_out8187,
   input         match_out8188,
   input         match_out8189,
   input         match_out8190,
   input         match_out8191,
   output        cfg_en0,
   output        cfg_en1,
   output        cfg_en2,
   output        cfg_en3,
   output        cfg_en4,
   output        cfg_en5,
   output        cfg_en6,
   output        cfg_en7,
   output        cfg_en8,
   output        cfg_en9,
   output        cfg_en10,
   output        cfg_en11,
   output        cfg_en12,
   output        cfg_en13,
   output        cfg_en14,
   output        cfg_en15,
   output        cfg_en16,
   output        cfg_en17,
   output        cfg_en18,
   output        cfg_en19,
   output        cfg_en20,
   output        cfg_en21,
   output        cfg_en22,
   output        cfg_en23,
   output        cfg_en24,
   output        cfg_en25,
   output        cfg_en26,
   output        cfg_en27,
   output        cfg_en28,
   output        cfg_en29,
   output        cfg_en30,
   output        cfg_en31,
   output        cfg_en32,
   output        cfg_en33,
   output        cfg_en34,
   output        cfg_en35,
   output        cfg_en36,
   output        cfg_en37,
   output        cfg_en38,
   output        cfg_en39,
   output        cfg_en40,
   output        cfg_en41,
   output        cfg_en42,
   output        cfg_en43,
   output        cfg_en44,
   output        cfg_en45,
   output        cfg_en46,
   output        cfg_en47,
   output        cfg_en48,
   output        cfg_en49,
   output        cfg_en50,
   output        cfg_en51,
   output        cfg_en52,
   output        cfg_en53,
   output        cfg_en54,
   output        cfg_en55,
   output        cfg_en56,
   output        cfg_en57,
   output        cfg_en58,
   output        cfg_en59,
   output        cfg_en60,
   output        cfg_en61,
   output        cfg_en62,
   output        cfg_en63,
   output        cfg_en64,
   output        cfg_en65,
   output        cfg_en66,
   output        cfg_en67,
   output        cfg_en68,
   output        cfg_en69,
   output        cfg_en70,
   output        cfg_en71,
   output        cfg_en72,
   output        cfg_en73,
   output        cfg_en74,
   output        cfg_en75,
   output        cfg_en76,
   output        cfg_en77,
   output        cfg_en78,
   output        cfg_en79,
   output        cfg_en80,
   output        cfg_en81,
   output        cfg_en82,
   output        cfg_en83,
   output        cfg_en84,
   output        cfg_en85,
   output        cfg_en86,
   output        cfg_en87,
   output        cfg_en88,
   output        cfg_en89,
   output        cfg_en90,
   output        cfg_en91,
   output        cfg_en92,
   output        cfg_en93,
   output        cfg_en94,
   output        cfg_en95,
   output        cfg_en96,
   output        cfg_en97,
   output        cfg_en98,
   output        cfg_en99,
   output        cfg_en100,
   output        cfg_en101,
   output        cfg_en102,
   output        cfg_en103,
   output        cfg_en104,
   output        cfg_en105,
   output        cfg_en106,
   output        cfg_en107,
   output        cfg_en108,
   output        cfg_en109,
   output        cfg_en110,
   output        cfg_en111,
   output        cfg_en112,
   output        cfg_en113,
   output        cfg_en114,
   output        cfg_en115,
   output        cfg_en116,
   output        cfg_en117,
   output        cfg_en118,
   output        cfg_en119,
   output        cfg_en120,
   output        cfg_en121,
   output        cfg_en122,
   output        cfg_en123,
   output        cfg_en124,
   output        cfg_en125,
   output        cfg_en126,
   output        cfg_en127,
   output        cfg_en128,
   output        cfg_en129,
   output        cfg_en130,
   output        cfg_en131,
   output        cfg_en132,
   output        cfg_en133,
   output        cfg_en134,
   output        cfg_en135,
   output        cfg_en136,
   output        cfg_en137,
   output        cfg_en138,
   output        cfg_en139,
   output        cfg_en140,
   output        cfg_en141,
   output        cfg_en142,
   output        cfg_en143,
   output        cfg_en144,
   output        cfg_en145,
   output        cfg_en146,
   output        cfg_en147,
   output        cfg_en148,
   output        cfg_en149,
   output        cfg_en150,
   output        cfg_en151,
   output        cfg_en152,
   output        cfg_en153,
   output        cfg_en154,
   output        cfg_en155,
   output        cfg_en156,
   output        cfg_en157,
   output        cfg_en158,
   output        cfg_en159,
   output        cfg_en160,
   output        cfg_en161,
   output        cfg_en162,
   output        cfg_en163,
   output        cfg_en164,
   output        cfg_en165,
   output        cfg_en166,
   output        cfg_en167,
   output        cfg_en168,
   output        cfg_en169,
   output        cfg_en170,
   output        cfg_en171,
   output        cfg_en172,
   output        cfg_en173,
   output        cfg_en174,
   output        cfg_en175,
   output        cfg_en176,
   output        cfg_en177,
   output        cfg_en178,
   output        cfg_en179,
   output        cfg_en180,
   output        cfg_en181,
   output        cfg_en182,
   output        cfg_en183,
   output        cfg_en184,
   output        cfg_en185,
   output        cfg_en186,
   output        cfg_en187,
   output        cfg_en188,
   output        cfg_en189,
   output        cfg_en190,
   output        cfg_en191,
   output        cfg_en192,
   output        cfg_en193,
   output        cfg_en194,
   output        cfg_en195,
   output        cfg_en196,
   output        cfg_en197,
   output        cfg_en198,
   output        cfg_en199,
   output        cfg_en200,
   output        cfg_en201,
   output        cfg_en202,
   output        cfg_en203,
   output        cfg_en204,
   output        cfg_en205,
   output        cfg_en206,
   output        cfg_en207,
   output        cfg_en208,
   output        cfg_en209,
   output        cfg_en210,
   output        cfg_en211,
   output        cfg_en212,
   output        cfg_en213,
   output        cfg_en214,
   output        cfg_en215,
   output        cfg_en216,
   output        cfg_en217,
   output        cfg_en218,
   output        cfg_en219,
   output        cfg_en220,
   output        cfg_en221,
   output        cfg_en222,
   output        cfg_en223,
   output        cfg_en224,
   output        cfg_en225,
   output        cfg_en226,
   output        cfg_en227,
   output        cfg_en228,
   output        cfg_en229,
   output        cfg_en230,
   output        cfg_en231,
   output        cfg_en232,
   output        cfg_en233,
   output        cfg_en234,
   output        cfg_en235,
   output        cfg_en236,
   output        cfg_en237,
   output        cfg_en238,
   output        cfg_en239,
   output        cfg_en240,
   output        cfg_en241,
   output        cfg_en242,
   output        cfg_en243,
   output        cfg_en244,
   output        cfg_en245,
   output        cfg_en246,
   output        cfg_en247,
   output        cfg_en248,
   output        cfg_en249,
   output        cfg_en250,
   output        cfg_en251,
   output        cfg_en252,
   output        cfg_en253,
   output        cfg_en254,
   output        cfg_en255,
   output        cfg_en256,
   output        cfg_en257,
   output        cfg_en258,
   output        cfg_en259,
   output        cfg_en260,
   output        cfg_en261,
   output        cfg_en262,
   output        cfg_en263,
   output        cfg_en264,
   output        cfg_en265,
   output        cfg_en266,
   output        cfg_en267,
   output        cfg_en268,
   output        cfg_en269,
   output        cfg_en270,
   output        cfg_en271,
   output        cfg_en272,
   output        cfg_en273,
   output        cfg_en274,
   output        cfg_en275,
   output        cfg_en276,
   output        cfg_en277,
   output        cfg_en278,
   output        cfg_en279,
   output        cfg_en280,
   output        cfg_en281,
   output        cfg_en282,
   output        cfg_en283,
   output        cfg_en284,
   output        cfg_en285,
   output        cfg_en286,
   output        cfg_en287,
   output        cfg_en288,
   output        cfg_en289,
   output        cfg_en290,
   output        cfg_en291,
   output        cfg_en292,
   output        cfg_en293,
   output        cfg_en294,
   output        cfg_en295,
   output        cfg_en296,
   output        cfg_en297,
   output        cfg_en298,
   output        cfg_en299,
   output        cfg_en300,
   output        cfg_en301,
   output        cfg_en302,
   output        cfg_en303,
   output        cfg_en304,
   output        cfg_en305,
   output        cfg_en306,
   output        cfg_en307,
   output        cfg_en308,
   output        cfg_en309,
   output        cfg_en310,
   output        cfg_en311,
   output        cfg_en312,
   output        cfg_en313,
   output        cfg_en314,
   output        cfg_en315,
   output        cfg_en316,
   output        cfg_en317,
   output        cfg_en318,
   output        cfg_en319,
   output        cfg_en320,
   output        cfg_en321,
   output        cfg_en322,
   output        cfg_en323,
   output        cfg_en324,
   output        cfg_en325,
   output        cfg_en326,
   output        cfg_en327,
   output        cfg_en328,
   output        cfg_en329,
   output        cfg_en330,
   output        cfg_en331,
   output        cfg_en332,
   output        cfg_en333,
   output        cfg_en334,
   output        cfg_en335,
   output        cfg_en336,
   output        cfg_en337,
   output        cfg_en338,
   output        cfg_en339,
   output        cfg_en340,
   output        cfg_en341,
   output        cfg_en342,
   output        cfg_en343,
   output        cfg_en344,
   output        cfg_en345,
   output        cfg_en346,
   output        cfg_en347,
   output        cfg_en348,
   output        cfg_en349,
   output        cfg_en350,
   output        cfg_en351,
   output        cfg_en352,
   output        cfg_en353,
   output        cfg_en354,
   output        cfg_en355,
   output        cfg_en356,
   output        cfg_en357,
   output        cfg_en358,
   output        cfg_en359,
   output        cfg_en360,
   output        cfg_en361,
   output        cfg_en362,
   output        cfg_en363,
   output        cfg_en364,
   output        cfg_en365,
   output        cfg_en366,
   output        cfg_en367,
   output        cfg_en368,
   output        cfg_en369,
   output        cfg_en370,
   output        cfg_en371,
   output        cfg_en372,
   output        cfg_en373,
   output        cfg_en374,
   output        cfg_en375,
   output        cfg_en376,
   output        cfg_en377,
   output        cfg_en378,
   output        cfg_en379,
   output        cfg_en380,
   output        cfg_en381,
   output        cfg_en382,
   output        cfg_en383,
   output        cfg_en384,
   output        cfg_en385,
   output        cfg_en386,
   output        cfg_en387,
   output        cfg_en388,
   output        cfg_en389,
   output        cfg_en390,
   output        cfg_en391,
   output        cfg_en392,
   output        cfg_en393,
   output        cfg_en394,
   output        cfg_en395,
   output        cfg_en396,
   output        cfg_en397,
   output        cfg_en398,
   output        cfg_en399,
   output        cfg_en400,
   output        cfg_en401,
   output        cfg_en402,
   output        cfg_en403,
   output        cfg_en404,
   output        cfg_en405,
   output        cfg_en406,
   output        cfg_en407,
   output        cfg_en408,
   output        cfg_en409,
   output        cfg_en410,
   output        cfg_en411,
   output        cfg_en412,
   output        cfg_en413,
   output        cfg_en414,
   output        cfg_en415,
   output        cfg_en416,
   output        cfg_en417,
   output        cfg_en418,
   output        cfg_en419,
   output        cfg_en420,
   output        cfg_en421,
   output        cfg_en422,
   output        cfg_en423,
   output        cfg_en424,
   output        cfg_en425,
   output        cfg_en426,
   output        cfg_en427,
   output        cfg_en428,
   output        cfg_en429,
   output        cfg_en430,
   output        cfg_en431,
   output        cfg_en432,
   output        cfg_en433,
   output        cfg_en434,
   output        cfg_en435,
   output        cfg_en436,
   output        cfg_en437,
   output        cfg_en438,
   output        cfg_en439,
   output        cfg_en440,
   output        cfg_en441,
   output        cfg_en442,
   output        cfg_en443,
   output        cfg_en444,
   output        cfg_en445,
   output        cfg_en446,
   output        cfg_en447,
   output        cfg_en448,
   output        cfg_en449,
   output        cfg_en450,
   output        cfg_en451,
   output        cfg_en452,
   output        cfg_en453,
   output        cfg_en454,
   output        cfg_en455,
   output        cfg_en456,
   output        cfg_en457,
   output        cfg_en458,
   output        cfg_en459,
   output        cfg_en460,
   output        cfg_en461,
   output        cfg_en462,
   output        cfg_en463,
   output        cfg_en464,
   output        cfg_en465,
   output        cfg_en466,
   output        cfg_en467,
   output        cfg_en468,
   output        cfg_en469,
   output        cfg_en470,
   output        cfg_en471,
   output        cfg_en472,
   output        cfg_en473,
   output        cfg_en474,
   output        cfg_en475,
   output        cfg_en476,
   output        cfg_en477,
   output        cfg_en478,
   output        cfg_en479,
   output        cfg_en480,
   output        cfg_en481,
   output        cfg_en482,
   output        cfg_en483,
   output        cfg_en484,
   output        cfg_en485,
   output        cfg_en486,
   output        cfg_en487,
   output        cfg_en488,
   output        cfg_en489,
   output        cfg_en490,
   output        cfg_en491,
   output        cfg_en492,
   output        cfg_en493,
   output        cfg_en494,
   output        cfg_en495,
   output        cfg_en496,
   output        cfg_en497,
   output        cfg_en498,
   output        cfg_en499,
   output        cfg_en500,
   output        cfg_en501,
   output        cfg_en502,
   output        cfg_en503,
   output        cfg_en504,
   output        cfg_en505,
   output        cfg_en506,
   output        cfg_en507,
   output        cfg_en508,
   output        cfg_en509,
   output        cfg_en510,
   output        cfg_en511,
   output        cfg_en512,
   output        cfg_en513,
   output        cfg_en514,
   output        cfg_en515,
   output        cfg_en516,
   output        cfg_en517,
   output        cfg_en518,
   output        cfg_en519,
   output        cfg_en520,
   output        cfg_en521,
   output        cfg_en522,
   output        cfg_en523,
   output        cfg_en524,
   output        cfg_en525,
   output        cfg_en526,
   output        cfg_en527,
   output        cfg_en528,
   output        cfg_en529,
   output        cfg_en530,
   output        cfg_en531,
   output        cfg_en532,
   output        cfg_en533,
   output        cfg_en534,
   output        cfg_en535,
   output        cfg_en536,
   output        cfg_en537,
   output        cfg_en538,
   output        cfg_en539,
   output        cfg_en540,
   output        cfg_en541,
   output        cfg_en542,
   output        cfg_en543,
   output        cfg_en544,
   output        cfg_en545,
   output        cfg_en546,
   output        cfg_en547,
   output        cfg_en548,
   output        cfg_en549,
   output        cfg_en550,
   output        cfg_en551,
   output        cfg_en552,
   output        cfg_en553,
   output        cfg_en554,
   output        cfg_en555,
   output        cfg_en556,
   output        cfg_en557,
   output        cfg_en558,
   output        cfg_en559,
   output        cfg_en560,
   output        cfg_en561,
   output        cfg_en562,
   output        cfg_en563,
   output        cfg_en564,
   output        cfg_en565,
   output        cfg_en566,
   output        cfg_en567,
   output        cfg_en568,
   output        cfg_en569,
   output        cfg_en570,
   output        cfg_en571,
   output        cfg_en572,
   output        cfg_en573,
   output        cfg_en574,
   output        cfg_en575,
   output        cfg_en576,
   output        cfg_en577,
   output        cfg_en578,
   output        cfg_en579,
   output        cfg_en580,
   output        cfg_en581,
   output        cfg_en582,
   output        cfg_en583,
   output        cfg_en584,
   output        cfg_en585,
   output        cfg_en586,
   output        cfg_en587,
   output        cfg_en588,
   output        cfg_en589,
   output        cfg_en590,
   output        cfg_en591,
   output        cfg_en592,
   output        cfg_en593,
   output        cfg_en594,
   output        cfg_en595,
   output        cfg_en596,
   output        cfg_en597,
   output        cfg_en598,
   output        cfg_en599,
   output        cfg_en600,
   output        cfg_en601,
   output        cfg_en602,
   output        cfg_en603,
   output        cfg_en604,
   output        cfg_en605,
   output        cfg_en606,
   output        cfg_en607,
   output        cfg_en608,
   output        cfg_en609,
   output        cfg_en610,
   output        cfg_en611,
   output        cfg_en612,
   output        cfg_en613,
   output        cfg_en614,
   output        cfg_en615,
   output        cfg_en616,
   output        cfg_en617,
   output        cfg_en618,
   output        cfg_en619,
   output        cfg_en620,
   output        cfg_en621,
   output        cfg_en622,
   output        cfg_en623,
   output        cfg_en624,
   output        cfg_en625,
   output        cfg_en626,
   output        cfg_en627,
   output        cfg_en628,
   output        cfg_en629,
   output        cfg_en630,
   output        cfg_en631,
   output        cfg_en632,
   output        cfg_en633,
   output        cfg_en634,
   output        cfg_en635,
   output        cfg_en636,
   output        cfg_en637,
   output        cfg_en638,
   output        cfg_en639,
   output        cfg_en640,
   output        cfg_en641,
   output        cfg_en642,
   output        cfg_en643,
   output        cfg_en644,
   output        cfg_en645,
   output        cfg_en646,
   output        cfg_en647,
   output        cfg_en648,
   output        cfg_en649,
   output        cfg_en650,
   output        cfg_en651,
   output        cfg_en652,
   output        cfg_en653,
   output        cfg_en654,
   output        cfg_en655,
   output        cfg_en656,
   output        cfg_en657,
   output        cfg_en658,
   output        cfg_en659,
   output        cfg_en660,
   output        cfg_en661,
   output        cfg_en662,
   output        cfg_en663,
   output        cfg_en664,
   output        cfg_en665,
   output        cfg_en666,
   output        cfg_en667,
   output        cfg_en668,
   output        cfg_en669,
   output        cfg_en670,
   output        cfg_en671,
   output        cfg_en672,
   output        cfg_en673,
   output        cfg_en674,
   output        cfg_en675,
   output        cfg_en676,
   output        cfg_en677,
   output        cfg_en678,
   output        cfg_en679,
   output        cfg_en680,
   output        cfg_en681,
   output        cfg_en682,
   output        cfg_en683,
   output        cfg_en684,
   output        cfg_en685,
   output        cfg_en686,
   output        cfg_en687,
   output        cfg_en688,
   output        cfg_en689,
   output        cfg_en690,
   output        cfg_en691,
   output        cfg_en692,
   output        cfg_en693,
   output        cfg_en694,
   output        cfg_en695,
   output        cfg_en696,
   output        cfg_en697,
   output        cfg_en698,
   output        cfg_en699,
   output        cfg_en700,
   output        cfg_en701,
   output        cfg_en702,
   output        cfg_en703,
   output        cfg_en704,
   output        cfg_en705,
   output        cfg_en706,
   output        cfg_en707,
   output        cfg_en708,
   output        cfg_en709,
   output        cfg_en710,
   output        cfg_en711,
   output        cfg_en712,
   output        cfg_en713,
   output        cfg_en714,
   output        cfg_en715,
   output        cfg_en716,
   output        cfg_en717,
   output        cfg_en718,
   output        cfg_en719,
   output        cfg_en720,
   output        cfg_en721,
   output        cfg_en722,
   output        cfg_en723,
   output        cfg_en724,
   output        cfg_en725,
   output        cfg_en726,
   output        cfg_en727,
   output        cfg_en728,
   output        cfg_en729,
   output        cfg_en730,
   output        cfg_en731,
   output        cfg_en732,
   output        cfg_en733,
   output        cfg_en734,
   output        cfg_en735,
   output        cfg_en736,
   output        cfg_en737,
   output        cfg_en738,
   output        cfg_en739,
   output        cfg_en740,
   output        cfg_en741,
   output        cfg_en742,
   output        cfg_en743,
   output        cfg_en744,
   output        cfg_en745,
   output        cfg_en746,
   output        cfg_en747,
   output        cfg_en748,
   output        cfg_en749,
   output        cfg_en750,
   output        cfg_en751,
   output        cfg_en752,
   output        cfg_en753,
   output        cfg_en754,
   output        cfg_en755,
   output        cfg_en756,
   output        cfg_en757,
   output        cfg_en758,
   output        cfg_en759,
   output        cfg_en760,
   output        cfg_en761,
   output        cfg_en762,
   output        cfg_en763,
   output        cfg_en764,
   output        cfg_en765,
   output        cfg_en766,
   output        cfg_en767,
   output        cfg_en768,
   output        cfg_en769,
   output        cfg_en770,
   output        cfg_en771,
   output        cfg_en772,
   output        cfg_en773,
   output        cfg_en774,
   output        cfg_en775,
   output        cfg_en776,
   output        cfg_en777,
   output        cfg_en778,
   output        cfg_en779,
   output        cfg_en780,
   output        cfg_en781,
   output        cfg_en782,
   output        cfg_en783,
   output        cfg_en784,
   output        cfg_en785,
   output        cfg_en786,
   output        cfg_en787,
   output        cfg_en788,
   output        cfg_en789,
   output        cfg_en790,
   output        cfg_en791,
   output        cfg_en792,
   output        cfg_en793,
   output        cfg_en794,
   output        cfg_en795,
   output        cfg_en796,
   output        cfg_en797,
   output        cfg_en798,
   output        cfg_en799,
   output        cfg_en800,
   output        cfg_en801,
   output        cfg_en802,
   output        cfg_en803,
   output        cfg_en804,
   output        cfg_en805,
   output        cfg_en806,
   output        cfg_en807,
   output        cfg_en808,
   output        cfg_en809,
   output        cfg_en810,
   output        cfg_en811,
   output        cfg_en812,
   output        cfg_en813,
   output        cfg_en814,
   output        cfg_en815,
   output        cfg_en816,
   output        cfg_en817,
   output        cfg_en818,
   output        cfg_en819,
   output        cfg_en820,
   output        cfg_en821,
   output        cfg_en822,
   output        cfg_en823,
   output        cfg_en824,
   output        cfg_en825,
   output        cfg_en826,
   output        cfg_en827,
   output        cfg_en828,
   output        cfg_en829,
   output        cfg_en830,
   output        cfg_en831,
   output        cfg_en832,
   output        cfg_en833,
   output        cfg_en834,
   output        cfg_en835,
   output        cfg_en836,
   output        cfg_en837,
   output        cfg_en838,
   output        cfg_en839,
   output        cfg_en840,
   output        cfg_en841,
   output        cfg_en842,
   output        cfg_en843,
   output        cfg_en844,
   output        cfg_en845,
   output        cfg_en846,
   output        cfg_en847,
   output        cfg_en848,
   output        cfg_en849,
   output        cfg_en850,
   output        cfg_en851,
   output        cfg_en852,
   output        cfg_en853,
   output        cfg_en854,
   output        cfg_en855,
   output        cfg_en856,
   output        cfg_en857,
   output        cfg_en858,
   output        cfg_en859,
   output        cfg_en860,
   output        cfg_en861,
   output        cfg_en862,
   output        cfg_en863,
   output        cfg_en864,
   output        cfg_en865,
   output        cfg_en866,
   output        cfg_en867,
   output        cfg_en868,
   output        cfg_en869,
   output        cfg_en870,
   output        cfg_en871,
   output        cfg_en872,
   output        cfg_en873,
   output        cfg_en874,
   output        cfg_en875,
   output        cfg_en876,
   output        cfg_en877,
   output        cfg_en878,
   output        cfg_en879,
   output        cfg_en880,
   output        cfg_en881,
   output        cfg_en882,
   output        cfg_en883,
   output        cfg_en884,
   output        cfg_en885,
   output        cfg_en886,
   output        cfg_en887,
   output        cfg_en888,
   output        cfg_en889,
   output        cfg_en890,
   output        cfg_en891,
   output        cfg_en892,
   output        cfg_en893,
   output        cfg_en894,
   output        cfg_en895,
   output        cfg_en896,
   output        cfg_en897,
   output        cfg_en898,
   output        cfg_en899,
   output        cfg_en900,
   output        cfg_en901,
   output        cfg_en902,
   output        cfg_en903,
   output        cfg_en904,
   output        cfg_en905,
   output        cfg_en906,
   output        cfg_en907,
   output        cfg_en908,
   output        cfg_en909,
   output        cfg_en910,
   output        cfg_en911,
   output        cfg_en912,
   output        cfg_en913,
   output        cfg_en914,
   output        cfg_en915,
   output        cfg_en916,
   output        cfg_en917,
   output        cfg_en918,
   output        cfg_en919,
   output        cfg_en920,
   output        cfg_en921,
   output        cfg_en922,
   output        cfg_en923,
   output        cfg_en924,
   output        cfg_en925,
   output        cfg_en926,
   output        cfg_en927,
   output        cfg_en928,
   output        cfg_en929,
   output        cfg_en930,
   output        cfg_en931,
   output        cfg_en932,
   output        cfg_en933,
   output        cfg_en934,
   output        cfg_en935,
   output        cfg_en936,
   output        cfg_en937,
   output        cfg_en938,
   output        cfg_en939,
   output        cfg_en940,
   output        cfg_en941,
   output        cfg_en942,
   output        cfg_en943,
   output        cfg_en944,
   output        cfg_en945,
   output        cfg_en946,
   output        cfg_en947,
   output        cfg_en948,
   output        cfg_en949,
   output        cfg_en950,
   output        cfg_en951,
   output        cfg_en952,
   output        cfg_en953,
   output        cfg_en954,
   output        cfg_en955,
   output        cfg_en956,
   output        cfg_en957,
   output        cfg_en958,
   output        cfg_en959,
   output        cfg_en960,
   output        cfg_en961,
   output        cfg_en962,
   output        cfg_en963,
   output        cfg_en964,
   output        cfg_en965,
   output        cfg_en966,
   output        cfg_en967,
   output        cfg_en968,
   output        cfg_en969,
   output        cfg_en970,
   output        cfg_en971,
   output        cfg_en972,
   output        cfg_en973,
   output        cfg_en974,
   output        cfg_en975,
   output        cfg_en976,
   output        cfg_en977,
   output        cfg_en978,
   output        cfg_en979,
   output        cfg_en980,
   output        cfg_en981,
   output        cfg_en982,
   output        cfg_en983,
   output        cfg_en984,
   output        cfg_en985,
   output        cfg_en986,
   output        cfg_en987,
   output        cfg_en988,
   output        cfg_en989,
   output        cfg_en990,
   output        cfg_en991,
   output        cfg_en992,
   output        cfg_en993,
   output        cfg_en994,
   output        cfg_en995,
   output        cfg_en996,
   output        cfg_en997,
   output        cfg_en998,
   output        cfg_en999,
   output        cfg_en1000,
   output        cfg_en1001,
   output        cfg_en1002,
   output        cfg_en1003,
   output        cfg_en1004,
   output        cfg_en1005,
   output        cfg_en1006,
   output        cfg_en1007,
   output        cfg_en1008,
   output        cfg_en1009,
   output        cfg_en1010,
   output        cfg_en1011,
   output        cfg_en1012,
   output        cfg_en1013,
   output        cfg_en1014,
   output        cfg_en1015,
   output        cfg_en1016,
   output        cfg_en1017,
   output        cfg_en1018,
   output        cfg_en1019,
   output        cfg_en1020,
   output        cfg_en1021,
   output        cfg_en1022,
   output        cfg_en1023,
   output        cfg_en1024,
   output        cfg_en1025,
   output        cfg_en1026,
   output        cfg_en1027,
   output        cfg_en1028,
   output        cfg_en1029,
   output        cfg_en1030,
   output        cfg_en1031,
   output        cfg_en1032,
   output        cfg_en1033,
   output        cfg_en1034,
   output        cfg_en1035,
   output        cfg_en1036,
   output        cfg_en1037,
   output        cfg_en1038,
   output        cfg_en1039,
   output        cfg_en1040,
   output        cfg_en1041,
   output        cfg_en1042,
   output        cfg_en1043,
   output        cfg_en1044,
   output        cfg_en1045,
   output        cfg_en1046,
   output        cfg_en1047,
   output        cfg_en1048,
   output        cfg_en1049,
   output        cfg_en1050,
   output        cfg_en1051,
   output        cfg_en1052,
   output        cfg_en1053,
   output        cfg_en1054,
   output        cfg_en1055,
   output        cfg_en1056,
   output        cfg_en1057,
   output        cfg_en1058,
   output        cfg_en1059,
   output        cfg_en1060,
   output        cfg_en1061,
   output        cfg_en1062,
   output        cfg_en1063,
   output        cfg_en1064,
   output        cfg_en1065,
   output        cfg_en1066,
   output        cfg_en1067,
   output        cfg_en1068,
   output        cfg_en1069,
   output        cfg_en1070,
   output        cfg_en1071,
   output        cfg_en1072,
   output        cfg_en1073,
   output        cfg_en1074,
   output        cfg_en1075,
   output        cfg_en1076,
   output        cfg_en1077,
   output        cfg_en1078,
   output        cfg_en1079,
   output        cfg_en1080,
   output        cfg_en1081,
   output        cfg_en1082,
   output        cfg_en1083,
   output        cfg_en1084,
   output        cfg_en1085,
   output        cfg_en1086,
   output        cfg_en1087,
   output        cfg_en1088,
   output        cfg_en1089,
   output        cfg_en1090,
   output        cfg_en1091,
   output        cfg_en1092,
   output        cfg_en1093,
   output        cfg_en1094,
   output        cfg_en1095,
   output        cfg_en1096,
   output        cfg_en1097,
   output        cfg_en1098,
   output        cfg_en1099,
   output        cfg_en1100,
   output        cfg_en1101,
   output        cfg_en1102,
   output        cfg_en1103,
   output        cfg_en1104,
   output        cfg_en1105,
   output        cfg_en1106,
   output        cfg_en1107,
   output        cfg_en1108,
   output        cfg_en1109,
   output        cfg_en1110,
   output        cfg_en1111,
   output        cfg_en1112,
   output        cfg_en1113,
   output        cfg_en1114,
   output        cfg_en1115,
   output        cfg_en1116,
   output        cfg_en1117,
   output        cfg_en1118,
   output        cfg_en1119,
   output        cfg_en1120,
   output        cfg_en1121,
   output        cfg_en1122,
   output        cfg_en1123,
   output        cfg_en1124,
   output        cfg_en1125,
   output        cfg_en1126,
   output        cfg_en1127,
   output        cfg_en1128,
   output        cfg_en1129,
   output        cfg_en1130,
   output        cfg_en1131,
   output        cfg_en1132,
   output        cfg_en1133,
   output        cfg_en1134,
   output        cfg_en1135,
   output        cfg_en1136,
   output        cfg_en1137,
   output        cfg_en1138,
   output        cfg_en1139,
   output        cfg_en1140,
   output        cfg_en1141,
   output        cfg_en1142,
   output        cfg_en1143,
   output        cfg_en1144,
   output        cfg_en1145,
   output        cfg_en1146,
   output        cfg_en1147,
   output        cfg_en1148,
   output        cfg_en1149,
   output        cfg_en1150,
   output        cfg_en1151,
   output        cfg_en1152,
   output        cfg_en1153,
   output        cfg_en1154,
   output        cfg_en1155,
   output        cfg_en1156,
   output        cfg_en1157,
   output        cfg_en1158,
   output        cfg_en1159,
   output        cfg_en1160,
   output        cfg_en1161,
   output        cfg_en1162,
   output        cfg_en1163,
   output        cfg_en1164,
   output        cfg_en1165,
   output        cfg_en1166,
   output        cfg_en1167,
   output        cfg_en1168,
   output        cfg_en1169,
   output        cfg_en1170,
   output        cfg_en1171,
   output        cfg_en1172,
   output        cfg_en1173,
   output        cfg_en1174,
   output        cfg_en1175,
   output        cfg_en1176,
   output        cfg_en1177,
   output        cfg_en1178,
   output        cfg_en1179,
   output        cfg_en1180,
   output        cfg_en1181,
   output        cfg_en1182,
   output        cfg_en1183,
   output        cfg_en1184,
   output        cfg_en1185,
   output        cfg_en1186,
   output        cfg_en1187,
   output        cfg_en1188,
   output        cfg_en1189,
   output        cfg_en1190,
   output        cfg_en1191,
   output        cfg_en1192,
   output        cfg_en1193,
   output        cfg_en1194,
   output        cfg_en1195,
   output        cfg_en1196,
   output        cfg_en1197,
   output        cfg_en1198,
   output        cfg_en1199,
   output        cfg_en1200,
   output        cfg_en1201,
   output        cfg_en1202,
   output        cfg_en1203,
   output        cfg_en1204,
   output        cfg_en1205,
   output        cfg_en1206,
   output        cfg_en1207,
   output        cfg_en1208,
   output        cfg_en1209,
   output        cfg_en1210,
   output        cfg_en1211,
   output        cfg_en1212,
   output        cfg_en1213,
   output        cfg_en1214,
   output        cfg_en1215,
   output        cfg_en1216,
   output        cfg_en1217,
   output        cfg_en1218,
   output        cfg_en1219,
   output        cfg_en1220,
   output        cfg_en1221,
   output        cfg_en1222,
   output        cfg_en1223,
   output        cfg_en1224,
   output        cfg_en1225,
   output        cfg_en1226,
   output        cfg_en1227,
   output        cfg_en1228,
   output        cfg_en1229,
   output        cfg_en1230,
   output        cfg_en1231,
   output        cfg_en1232,
   output        cfg_en1233,
   output        cfg_en1234,
   output        cfg_en1235,
   output        cfg_en1236,
   output        cfg_en1237,
   output        cfg_en1238,
   output        cfg_en1239,
   output        cfg_en1240,
   output        cfg_en1241,
   output        cfg_en1242,
   output        cfg_en1243,
   output        cfg_en1244,
   output        cfg_en1245,
   output        cfg_en1246,
   output        cfg_en1247,
   output        cfg_en1248,
   output        cfg_en1249,
   output        cfg_en1250,
   output        cfg_en1251,
   output        cfg_en1252,
   output        cfg_en1253,
   output        cfg_en1254,
   output        cfg_en1255,
   output        cfg_en1256,
   output        cfg_en1257,
   output        cfg_en1258,
   output        cfg_en1259,
   output        cfg_en1260,
   output        cfg_en1261,
   output        cfg_en1262,
   output        cfg_en1263,
   output        cfg_en1264,
   output        cfg_en1265,
   output        cfg_en1266,
   output        cfg_en1267,
   output        cfg_en1268,
   output        cfg_en1269,
   output        cfg_en1270,
   output        cfg_en1271,
   output        cfg_en1272,
   output        cfg_en1273,
   output        cfg_en1274,
   output        cfg_en1275,
   output        cfg_en1276,
   output        cfg_en1277,
   output        cfg_en1278,
   output        cfg_en1279,
   output        cfg_en1280,
   output        cfg_en1281,
   output        cfg_en1282,
   output        cfg_en1283,
   output        cfg_en1284,
   output        cfg_en1285,
   output        cfg_en1286,
   output        cfg_en1287,
   output        cfg_en1288,
   output        cfg_en1289,
   output        cfg_en1290,
   output        cfg_en1291,
   output        cfg_en1292,
   output        cfg_en1293,
   output        cfg_en1294,
   output        cfg_en1295,
   output        cfg_en1296,
   output        cfg_en1297,
   output        cfg_en1298,
   output        cfg_en1299,
   output        cfg_en1300,
   output        cfg_en1301,
   output        cfg_en1302,
   output        cfg_en1303,
   output        cfg_en1304,
   output        cfg_en1305,
   output        cfg_en1306,
   output        cfg_en1307,
   output        cfg_en1308,
   output        cfg_en1309,
   output        cfg_en1310,
   output        cfg_en1311,
   output        cfg_en1312,
   output        cfg_en1313,
   output        cfg_en1314,
   output        cfg_en1315,
   output        cfg_en1316,
   output        cfg_en1317,
   output        cfg_en1318,
   output        cfg_en1319,
   output        cfg_en1320,
   output        cfg_en1321,
   output        cfg_en1322,
   output        cfg_en1323,
   output        cfg_en1324,
   output        cfg_en1325,
   output        cfg_en1326,
   output        cfg_en1327,
   output        cfg_en1328,
   output        cfg_en1329,
   output        cfg_en1330,
   output        cfg_en1331,
   output        cfg_en1332,
   output        cfg_en1333,
   output        cfg_en1334,
   output        cfg_en1335,
   output        cfg_en1336,
   output        cfg_en1337,
   output        cfg_en1338,
   output        cfg_en1339,
   output        cfg_en1340,
   output        cfg_en1341,
   output        cfg_en1342,
   output        cfg_en1343,
   output        cfg_en1344,
   output        cfg_en1345,
   output        cfg_en1346,
   output        cfg_en1347,
   output        cfg_en1348,
   output        cfg_en1349,
   output        cfg_en1350,
   output        cfg_en1351,
   output        cfg_en1352,
   output        cfg_en1353,
   output        cfg_en1354,
   output        cfg_en1355,
   output        cfg_en1356,
   output        cfg_en1357,
   output        cfg_en1358,
   output        cfg_en1359,
   output        cfg_en1360,
   output        cfg_en1361,
   output        cfg_en1362,
   output        cfg_en1363,
   output        cfg_en1364,
   output        cfg_en1365,
   output        cfg_en1366,
   output        cfg_en1367,
   output        cfg_en1368,
   output        cfg_en1369,
   output        cfg_en1370,
   output        cfg_en1371,
   output        cfg_en1372,
   output        cfg_en1373,
   output        cfg_en1374,
   output        cfg_en1375,
   output        cfg_en1376,
   output        cfg_en1377,
   output        cfg_en1378,
   output        cfg_en1379,
   output        cfg_en1380,
   output        cfg_en1381,
   output        cfg_en1382,
   output        cfg_en1383,
   output        cfg_en1384,
   output        cfg_en1385,
   output        cfg_en1386,
   output        cfg_en1387,
   output        cfg_en1388,
   output        cfg_en1389,
   output        cfg_en1390,
   output        cfg_en1391,
   output        cfg_en1392,
   output        cfg_en1393,
   output        cfg_en1394,
   output        cfg_en1395,
   output        cfg_en1396,
   output        cfg_en1397,
   output        cfg_en1398,
   output        cfg_en1399,
   output        cfg_en1400,
   output        cfg_en1401,
   output        cfg_en1402,
   output        cfg_en1403,
   output        cfg_en1404,
   output        cfg_en1405,
   output        cfg_en1406,
   output        cfg_en1407,
   output        cfg_en1408,
   output        cfg_en1409,
   output        cfg_en1410,
   output        cfg_en1411,
   output        cfg_en1412,
   output        cfg_en1413,
   output        cfg_en1414,
   output        cfg_en1415,
   output        cfg_en1416,
   output        cfg_en1417,
   output        cfg_en1418,
   output        cfg_en1419,
   output        cfg_en1420,
   output        cfg_en1421,
   output        cfg_en1422,
   output        cfg_en1423,
   output        cfg_en1424,
   output        cfg_en1425,
   output        cfg_en1426,
   output        cfg_en1427,
   output        cfg_en1428,
   output        cfg_en1429,
   output        cfg_en1430,
   output        cfg_en1431,
   output        cfg_en1432,
   output        cfg_en1433,
   output        cfg_en1434,
   output        cfg_en1435,
   output        cfg_en1436,
   output        cfg_en1437,
   output        cfg_en1438,
   output        cfg_en1439,
   output        cfg_en1440,
   output        cfg_en1441,
   output        cfg_en1442,
   output        cfg_en1443,
   output        cfg_en1444,
   output        cfg_en1445,
   output        cfg_en1446,
   output        cfg_en1447,
   output        cfg_en1448,
   output        cfg_en1449,
   output        cfg_en1450,
   output        cfg_en1451,
   output        cfg_en1452,
   output        cfg_en1453,
   output        cfg_en1454,
   output        cfg_en1455,
   output        cfg_en1456,
   output        cfg_en1457,
   output        cfg_en1458,
   output        cfg_en1459,
   output        cfg_en1460,
   output        cfg_en1461,
   output        cfg_en1462,
   output        cfg_en1463,
   output        cfg_en1464,
   output        cfg_en1465,
   output        cfg_en1466,
   output        cfg_en1467,
   output        cfg_en1468,
   output        cfg_en1469,
   output        cfg_en1470,
   output        cfg_en1471,
   output        cfg_en1472,
   output        cfg_en1473,
   output        cfg_en1474,
   output        cfg_en1475,
   output        cfg_en1476,
   output        cfg_en1477,
   output        cfg_en1478,
   output        cfg_en1479,
   output        cfg_en1480,
   output        cfg_en1481,
   output        cfg_en1482,
   output        cfg_en1483,
   output        cfg_en1484,
   output        cfg_en1485,
   output        cfg_en1486,
   output        cfg_en1487,
   output        cfg_en1488,
   output        cfg_en1489,
   output        cfg_en1490,
   output        cfg_en1491,
   output        cfg_en1492,
   output        cfg_en1493,
   output        cfg_en1494,
   output        cfg_en1495,
   output        cfg_en1496,
   output        cfg_en1497,
   output        cfg_en1498,
   output        cfg_en1499,
   output        cfg_en1500,
   output        cfg_en1501,
   output        cfg_en1502,
   output        cfg_en1503,
   output        cfg_en1504,
   output        cfg_en1505,
   output        cfg_en1506,
   output        cfg_en1507,
   output        cfg_en1508,
   output        cfg_en1509,
   output        cfg_en1510,
   output        cfg_en1511,
   output        cfg_en1512,
   output        cfg_en1513,
   output        cfg_en1514,
   output        cfg_en1515,
   output        cfg_en1516,
   output        cfg_en1517,
   output        cfg_en1518,
   output        cfg_en1519,
   output        cfg_en1520,
   output        cfg_en1521,
   output        cfg_en1522,
   output        cfg_en1523,
   output        cfg_en1524,
   output        cfg_en1525,
   output        cfg_en1526,
   output        cfg_en1527,
   output        cfg_en1528,
   output        cfg_en1529,
   output        cfg_en1530,
   output        cfg_en1531,
   output        cfg_en1532,
   output        cfg_en1533,
   output        cfg_en1534,
   output        cfg_en1535,
   output        cfg_en1536,
   output        cfg_en1537,
   output        cfg_en1538,
   output        cfg_en1539,
   output        cfg_en1540,
   output        cfg_en1541,
   output        cfg_en1542,
   output        cfg_en1543,
   output        cfg_en1544,
   output        cfg_en1545,
   output        cfg_en1546,
   output        cfg_en1547,
   output        cfg_en1548,
   output        cfg_en1549,
   output        cfg_en1550,
   output        cfg_en1551,
   output        cfg_en1552,
   output        cfg_en1553,
   output        cfg_en1554,
   output        cfg_en1555,
   output        cfg_en1556,
   output        cfg_en1557,
   output        cfg_en1558,
   output        cfg_en1559,
   output        cfg_en1560,
   output        cfg_en1561,
   output        cfg_en1562,
   output        cfg_en1563,
   output        cfg_en1564,
   output        cfg_en1565,
   output        cfg_en1566,
   output        cfg_en1567,
   output        cfg_en1568,
   output        cfg_en1569,
   output        cfg_en1570,
   output        cfg_en1571,
   output        cfg_en1572,
   output        cfg_en1573,
   output        cfg_en1574,
   output        cfg_en1575,
   output        cfg_en1576,
   output        cfg_en1577,
   output        cfg_en1578,
   output        cfg_en1579,
   output        cfg_en1580,
   output        cfg_en1581,
   output        cfg_en1582,
   output        cfg_en1583,
   output        cfg_en1584,
   output        cfg_en1585,
   output        cfg_en1586,
   output        cfg_en1587,
   output        cfg_en1588,
   output        cfg_en1589,
   output        cfg_en1590,
   output        cfg_en1591,
   output        cfg_en1592,
   output        cfg_en1593,
   output        cfg_en1594,
   output        cfg_en1595,
   output        cfg_en1596,
   output        cfg_en1597,
   output        cfg_en1598,
   output        cfg_en1599,
   output        cfg_en1600,
   output        cfg_en1601,
   output        cfg_en1602,
   output        cfg_en1603,
   output        cfg_en1604,
   output        cfg_en1605,
   output        cfg_en1606,
   output        cfg_en1607,
   output        cfg_en1608,
   output        cfg_en1609,
   output        cfg_en1610,
   output        cfg_en1611,
   output        cfg_en1612,
   output        cfg_en1613,
   output        cfg_en1614,
   output        cfg_en1615,
   output        cfg_en1616,
   output        cfg_en1617,
   output        cfg_en1618,
   output        cfg_en1619,
   output        cfg_en1620,
   output        cfg_en1621,
   output        cfg_en1622,
   output        cfg_en1623,
   output        cfg_en1624,
   output        cfg_en1625,
   output        cfg_en1626,
   output        cfg_en1627,
   output        cfg_en1628,
   output        cfg_en1629,
   output        cfg_en1630,
   output        cfg_en1631,
   output        cfg_en1632,
   output        cfg_en1633,
   output        cfg_en1634,
   output        cfg_en1635,
   output        cfg_en1636,
   output        cfg_en1637,
   output        cfg_en1638,
   output        cfg_en1639,
   output        cfg_en1640,
   output        cfg_en1641,
   output        cfg_en1642,
   output        cfg_en1643,
   output        cfg_en1644,
   output        cfg_en1645,
   output        cfg_en1646,
   output        cfg_en1647,
   output        cfg_en1648,
   output        cfg_en1649,
   output        cfg_en1650,
   output        cfg_en1651,
   output        cfg_en1652,
   output        cfg_en1653,
   output        cfg_en1654,
   output        cfg_en1655,
   output        cfg_en1656,
   output        cfg_en1657,
   output        cfg_en1658,
   output        cfg_en1659,
   output        cfg_en1660,
   output        cfg_en1661,
   output        cfg_en1662,
   output        cfg_en1663,
   output        cfg_en1664,
   output        cfg_en1665,
   output        cfg_en1666,
   output        cfg_en1667,
   output        cfg_en1668,
   output        cfg_en1669,
   output        cfg_en1670,
   output        cfg_en1671,
   output        cfg_en1672,
   output        cfg_en1673,
   output        cfg_en1674,
   output        cfg_en1675,
   output        cfg_en1676,
   output        cfg_en1677,
   output        cfg_en1678,
   output        cfg_en1679,
   output        cfg_en1680,
   output        cfg_en1681,
   output        cfg_en1682,
   output        cfg_en1683,
   output        cfg_en1684,
   output        cfg_en1685,
   output        cfg_en1686,
   output        cfg_en1687,
   output        cfg_en1688,
   output        cfg_en1689,
   output        cfg_en1690,
   output        cfg_en1691,
   output        cfg_en1692,
   output        cfg_en1693,
   output        cfg_en1694,
   output        cfg_en1695,
   output        cfg_en1696,
   output        cfg_en1697,
   output        cfg_en1698,
   output        cfg_en1699,
   output        cfg_en1700,
   output        cfg_en1701,
   output        cfg_en1702,
   output        cfg_en1703,
   output        cfg_en1704,
   output        cfg_en1705,
   output        cfg_en1706,
   output        cfg_en1707,
   output        cfg_en1708,
   output        cfg_en1709,
   output        cfg_en1710,
   output        cfg_en1711,
   output        cfg_en1712,
   output        cfg_en1713,
   output        cfg_en1714,
   output        cfg_en1715,
   output        cfg_en1716,
   output        cfg_en1717,
   output        cfg_en1718,
   output        cfg_en1719,
   output        cfg_en1720,
   output        cfg_en1721,
   output        cfg_en1722,
   output        cfg_en1723,
   output        cfg_en1724,
   output        cfg_en1725,
   output        cfg_en1726,
   output        cfg_en1727,
   output        cfg_en1728,
   output        cfg_en1729,
   output        cfg_en1730,
   output        cfg_en1731,
   output        cfg_en1732,
   output        cfg_en1733,
   output        cfg_en1734,
   output        cfg_en1735,
   output        cfg_en1736,
   output        cfg_en1737,
   output        cfg_en1738,
   output        cfg_en1739,
   output        cfg_en1740,
   output        cfg_en1741,
   output        cfg_en1742,
   output        cfg_en1743,
   output        cfg_en1744,
   output        cfg_en1745,
   output        cfg_en1746,
   output        cfg_en1747,
   output        cfg_en1748,
   output        cfg_en1749,
   output        cfg_en1750,
   output        cfg_en1751,
   output        cfg_en1752,
   output        cfg_en1753,
   output        cfg_en1754,
   output        cfg_en1755,
   output        cfg_en1756,
   output        cfg_en1757,
   output        cfg_en1758,
   output        cfg_en1759,
   output        cfg_en1760,
   output        cfg_en1761,
   output        cfg_en1762,
   output        cfg_en1763,
   output        cfg_en1764,
   output        cfg_en1765,
   output        cfg_en1766,
   output        cfg_en1767,
   output        cfg_en1768,
   output        cfg_en1769,
   output        cfg_en1770,
   output        cfg_en1771,
   output        cfg_en1772,
   output        cfg_en1773,
   output        cfg_en1774,
   output        cfg_en1775,
   output        cfg_en1776,
   output        cfg_en1777,
   output        cfg_en1778,
   output        cfg_en1779,
   output        cfg_en1780,
   output        cfg_en1781,
   output        cfg_en1782,
   output        cfg_en1783,
   output        cfg_en1784,
   output        cfg_en1785,
   output        cfg_en1786,
   output        cfg_en1787,
   output        cfg_en1788,
   output        cfg_en1789,
   output        cfg_en1790,
   output        cfg_en1791,
   output        cfg_en1792,
   output        cfg_en1793,
   output        cfg_en1794,
   output        cfg_en1795,
   output        cfg_en1796,
   output        cfg_en1797,
   output        cfg_en1798,
   output        cfg_en1799,
   output        cfg_en1800,
   output        cfg_en1801,
   output        cfg_en1802,
   output        cfg_en1803,
   output        cfg_en1804,
   output        cfg_en1805,
   output        cfg_en1806,
   output        cfg_en1807,
   output        cfg_en1808,
   output        cfg_en1809,
   output        cfg_en1810,
   output        cfg_en1811,
   output        cfg_en1812,
   output        cfg_en1813,
   output        cfg_en1814,
   output        cfg_en1815,
   output        cfg_en1816,
   output        cfg_en1817,
   output        cfg_en1818,
   output        cfg_en1819,
   output        cfg_en1820,
   output        cfg_en1821,
   output        cfg_en1822,
   output        cfg_en1823,
   output        cfg_en1824,
   output        cfg_en1825,
   output        cfg_en1826,
   output        cfg_en1827,
   output        cfg_en1828,
   output        cfg_en1829,
   output        cfg_en1830,
   output        cfg_en1831,
   output        cfg_en1832,
   output        cfg_en1833,
   output        cfg_en1834,
   output        cfg_en1835,
   output        cfg_en1836,
   output        cfg_en1837,
   output        cfg_en1838,
   output        cfg_en1839,
   output        cfg_en1840,
   output        cfg_en1841,
   output        cfg_en1842,
   output        cfg_en1843,
   output        cfg_en1844,
   output        cfg_en1845,
   output        cfg_en1846,
   output        cfg_en1847,
   output        cfg_en1848,
   output        cfg_en1849,
   output        cfg_en1850,
   output        cfg_en1851,
   output        cfg_en1852,
   output        cfg_en1853,
   output        cfg_en1854,
   output        cfg_en1855,
   output        cfg_en1856,
   output        cfg_en1857,
   output        cfg_en1858,
   output        cfg_en1859,
   output        cfg_en1860,
   output        cfg_en1861,
   output        cfg_en1862,
   output        cfg_en1863,
   output        cfg_en1864,
   output        cfg_en1865,
   output        cfg_en1866,
   output        cfg_en1867,
   output        cfg_en1868,
   output        cfg_en1869,
   output        cfg_en1870,
   output        cfg_en1871,
   output        cfg_en1872,
   output        cfg_en1873,
   output        cfg_en1874,
   output        cfg_en1875,
   output        cfg_en1876,
   output        cfg_en1877,
   output        cfg_en1878,
   output        cfg_en1879,
   output        cfg_en1880,
   output        cfg_en1881,
   output        cfg_en1882,
   output        cfg_en1883,
   output        cfg_en1884,
   output        cfg_en1885,
   output        cfg_en1886,
   output        cfg_en1887,
   output        cfg_en1888,
   output        cfg_en1889,
   output        cfg_en1890,
   output        cfg_en1891,
   output        cfg_en1892,
   output        cfg_en1893,
   output        cfg_en1894,
   output        cfg_en1895,
   output        cfg_en1896,
   output        cfg_en1897,
   output        cfg_en1898,
   output        cfg_en1899,
   output        cfg_en1900,
   output        cfg_en1901,
   output        cfg_en1902,
   output        cfg_en1903,
   output        cfg_en1904,
   output        cfg_en1905,
   output        cfg_en1906,
   output        cfg_en1907,
   output        cfg_en1908,
   output        cfg_en1909,
   output        cfg_en1910,
   output        cfg_en1911,
   output        cfg_en1912,
   output        cfg_en1913,
   output        cfg_en1914,
   output        cfg_en1915,
   output        cfg_en1916,
   output        cfg_en1917,
   output        cfg_en1918,
   output        cfg_en1919,
   output        cfg_en1920,
   output        cfg_en1921,
   output        cfg_en1922,
   output        cfg_en1923,
   output        cfg_en1924,
   output        cfg_en1925,
   output        cfg_en1926,
   output        cfg_en1927,
   output        cfg_en1928,
   output        cfg_en1929,
   output        cfg_en1930,
   output        cfg_en1931,
   output        cfg_en1932,
   output        cfg_en1933,
   output        cfg_en1934,
   output        cfg_en1935,
   output        cfg_en1936,
   output        cfg_en1937,
   output        cfg_en1938,
   output        cfg_en1939,
   output        cfg_en1940,
   output        cfg_en1941,
   output        cfg_en1942,
   output        cfg_en1943,
   output        cfg_en1944,
   output        cfg_en1945,
   output        cfg_en1946,
   output        cfg_en1947,
   output        cfg_en1948,
   output        cfg_en1949,
   output        cfg_en1950,
   output        cfg_en1951,
   output        cfg_en1952,
   output        cfg_en1953,
   output        cfg_en1954,
   output        cfg_en1955,
   output        cfg_en1956,
   output        cfg_en1957,
   output        cfg_en1958,
   output        cfg_en1959,
   output        cfg_en1960,
   output        cfg_en1961,
   output        cfg_en1962,
   output        cfg_en1963,
   output        cfg_en1964,
   output        cfg_en1965,
   output        cfg_en1966,
   output        cfg_en1967,
   output        cfg_en1968,
   output        cfg_en1969,
   output        cfg_en1970,
   output        cfg_en1971,
   output        cfg_en1972,
   output        cfg_en1973,
   output        cfg_en1974,
   output        cfg_en1975,
   output        cfg_en1976,
   output        cfg_en1977,
   output        cfg_en1978,
   output        cfg_en1979,
   output        cfg_en1980,
   output        cfg_en1981,
   output        cfg_en1982,
   output        cfg_en1983,
   output        cfg_en1984,
   output        cfg_en1985,
   output        cfg_en1986,
   output        cfg_en1987,
   output        cfg_en1988,
   output        cfg_en1989,
   output        cfg_en1990,
   output        cfg_en1991,
   output        cfg_en1992,
   output        cfg_en1993,
   output        cfg_en1994,
   output        cfg_en1995,
   output        cfg_en1996,
   output        cfg_en1997,
   output        cfg_en1998,
   output        cfg_en1999,
   output        cfg_en2000,
   output        cfg_en2001,
   output        cfg_en2002,
   output        cfg_en2003,
   output        cfg_en2004,
   output        cfg_en2005,
   output        cfg_en2006,
   output        cfg_en2007,
   output        cfg_en2008,
   output        cfg_en2009,
   output        cfg_en2010,
   output        cfg_en2011,
   output        cfg_en2012,
   output        cfg_en2013,
   output        cfg_en2014,
   output        cfg_en2015,
   output        cfg_en2016,
   output        cfg_en2017,
   output        cfg_en2018,
   output        cfg_en2019,
   output        cfg_en2020,
   output        cfg_en2021,
   output        cfg_en2022,
   output        cfg_en2023,
   output        cfg_en2024,
   output        cfg_en2025,
   output        cfg_en2026,
   output        cfg_en2027,
   output        cfg_en2028,
   output        cfg_en2029,
   output        cfg_en2030,
   output        cfg_en2031,
   output        cfg_en2032,
   output        cfg_en2033,
   output        cfg_en2034,
   output        cfg_en2035,
   output        cfg_en2036,
   output        cfg_en2037,
   output        cfg_en2038,
   output        cfg_en2039,
   output        cfg_en2040,
   output        cfg_en2041,
   output        cfg_en2042,
   output        cfg_en2043,
   output        cfg_en2044,
   output        cfg_en2045,
   output        cfg_en2046,
   output        cfg_en2047,
   output        cfg_en2048,
   output        cfg_en2049,
   output        cfg_en2050,
   output        cfg_en2051,
   output        cfg_en2052,
   output        cfg_en2053,
   output        cfg_en2054,
   output        cfg_en2055,
   output        cfg_en2056,
   output        cfg_en2057,
   output        cfg_en2058,
   output        cfg_en2059,
   output        cfg_en2060,
   output        cfg_en2061,
   output        cfg_en2062,
   output        cfg_en2063,
   output        cfg_en2064,
   output        cfg_en2065,
   output        cfg_en2066,
   output        cfg_en2067,
   output        cfg_en2068,
   output        cfg_en2069,
   output        cfg_en2070,
   output        cfg_en2071,
   output        cfg_en2072,
   output        cfg_en2073,
   output        cfg_en2074,
   output        cfg_en2075,
   output        cfg_en2076,
   output        cfg_en2077,
   output        cfg_en2078,
   output        cfg_en2079,
   output        cfg_en2080,
   output        cfg_en2081,
   output        cfg_en2082,
   output        cfg_en2083,
   output        cfg_en2084,
   output        cfg_en2085,
   output        cfg_en2086,
   output        cfg_en2087,
   output        cfg_en2088,
   output        cfg_en2089,
   output        cfg_en2090,
   output        cfg_en2091,
   output        cfg_en2092,
   output        cfg_en2093,
   output        cfg_en2094,
   output        cfg_en2095,
   output        cfg_en2096,
   output        cfg_en2097,
   output        cfg_en2098,
   output        cfg_en2099,
   output        cfg_en2100,
   output        cfg_en2101,
   output        cfg_en2102,
   output        cfg_en2103,
   output        cfg_en2104,
   output        cfg_en2105,
   output        cfg_en2106,
   output        cfg_en2107,
   output        cfg_en2108,
   output        cfg_en2109,
   output        cfg_en2110,
   output        cfg_en2111,
   output        cfg_en2112,
   output        cfg_en2113,
   output        cfg_en2114,
   output        cfg_en2115,
   output        cfg_en2116,
   output        cfg_en2117,
   output        cfg_en2118,
   output        cfg_en2119,
   output        cfg_en2120,
   output        cfg_en2121,
   output        cfg_en2122,
   output        cfg_en2123,
   output        cfg_en2124,
   output        cfg_en2125,
   output        cfg_en2126,
   output        cfg_en2127,
   output        cfg_en2128,
   output        cfg_en2129,
   output        cfg_en2130,
   output        cfg_en2131,
   output        cfg_en2132,
   output        cfg_en2133,
   output        cfg_en2134,
   output        cfg_en2135,
   output        cfg_en2136,
   output        cfg_en2137,
   output        cfg_en2138,
   output        cfg_en2139,
   output        cfg_en2140,
   output        cfg_en2141,
   output        cfg_en2142,
   output        cfg_en2143,
   output        cfg_en2144,
   output        cfg_en2145,
   output        cfg_en2146,
   output        cfg_en2147,
   output        cfg_en2148,
   output        cfg_en2149,
   output        cfg_en2150,
   output        cfg_en2151,
   output        cfg_en2152,
   output        cfg_en2153,
   output        cfg_en2154,
   output        cfg_en2155,
   output        cfg_en2156,
   output        cfg_en2157,
   output        cfg_en2158,
   output        cfg_en2159,
   output        cfg_en2160,
   output        cfg_en2161,
   output        cfg_en2162,
   output        cfg_en2163,
   output        cfg_en2164,
   output        cfg_en2165,
   output        cfg_en2166,
   output        cfg_en2167,
   output        cfg_en2168,
   output        cfg_en2169,
   output        cfg_en2170,
   output        cfg_en2171,
   output        cfg_en2172,
   output        cfg_en2173,
   output        cfg_en2174,
   output        cfg_en2175,
   output        cfg_en2176,
   output        cfg_en2177,
   output        cfg_en2178,
   output        cfg_en2179,
   output        cfg_en2180,
   output        cfg_en2181,
   output        cfg_en2182,
   output        cfg_en2183,
   output        cfg_en2184,
   output        cfg_en2185,
   output        cfg_en2186,
   output        cfg_en2187,
   output        cfg_en2188,
   output        cfg_en2189,
   output        cfg_en2190,
   output        cfg_en2191,
   output        cfg_en2192,
   output        cfg_en2193,
   output        cfg_en2194,
   output        cfg_en2195,
   output        cfg_en2196,
   output        cfg_en2197,
   output        cfg_en2198,
   output        cfg_en2199,
   output        cfg_en2200,
   output        cfg_en2201,
   output        cfg_en2202,
   output        cfg_en2203,
   output        cfg_en2204,
   output        cfg_en2205,
   output        cfg_en2206,
   output        cfg_en2207,
   output        cfg_en2208,
   output        cfg_en2209,
   output        cfg_en2210,
   output        cfg_en2211,
   output        cfg_en2212,
   output        cfg_en2213,
   output        cfg_en2214,
   output        cfg_en2215,
   output        cfg_en2216,
   output        cfg_en2217,
   output        cfg_en2218,
   output        cfg_en2219,
   output        cfg_en2220,
   output        cfg_en2221,
   output        cfg_en2222,
   output        cfg_en2223,
   output        cfg_en2224,
   output        cfg_en2225,
   output        cfg_en2226,
   output        cfg_en2227,
   output        cfg_en2228,
   output        cfg_en2229,
   output        cfg_en2230,
   output        cfg_en2231,
   output        cfg_en2232,
   output        cfg_en2233,
   output        cfg_en2234,
   output        cfg_en2235,
   output        cfg_en2236,
   output        cfg_en2237,
   output        cfg_en2238,
   output        cfg_en2239,
   output        cfg_en2240,
   output        cfg_en2241,
   output        cfg_en2242,
   output        cfg_en2243,
   output        cfg_en2244,
   output        cfg_en2245,
   output        cfg_en2246,
   output        cfg_en2247,
   output        cfg_en2248,
   output        cfg_en2249,
   output        cfg_en2250,
   output        cfg_en2251,
   output        cfg_en2252,
   output        cfg_en2253,
   output        cfg_en2254,
   output        cfg_en2255,
   output        cfg_en2256,
   output        cfg_en2257,
   output        cfg_en2258,
   output        cfg_en2259,
   output        cfg_en2260,
   output        cfg_en2261,
   output        cfg_en2262,
   output        cfg_en2263,
   output        cfg_en2264,
   output        cfg_en2265,
   output        cfg_en2266,
   output        cfg_en2267,
   output        cfg_en2268,
   output        cfg_en2269,
   output        cfg_en2270,
   output        cfg_en2271,
   output        cfg_en2272,
   output        cfg_en2273,
   output        cfg_en2274,
   output        cfg_en2275,
   output        cfg_en2276,
   output        cfg_en2277,
   output        cfg_en2278,
   output        cfg_en2279,
   output        cfg_en2280,
   output        cfg_en2281,
   output        cfg_en2282,
   output        cfg_en2283,
   output        cfg_en2284,
   output        cfg_en2285,
   output        cfg_en2286,
   output        cfg_en2287,
   output        cfg_en2288,
   output        cfg_en2289,
   output        cfg_en2290,
   output        cfg_en2291,
   output        cfg_en2292,
   output        cfg_en2293,
   output        cfg_en2294,
   output        cfg_en2295,
   output        cfg_en2296,
   output        cfg_en2297,
   output        cfg_en2298,
   output        cfg_en2299,
   output        cfg_en2300,
   output        cfg_en2301,
   output        cfg_en2302,
   output        cfg_en2303,
   output        cfg_en2304,
   output        cfg_en2305,
   output        cfg_en2306,
   output        cfg_en2307,
   output        cfg_en2308,
   output        cfg_en2309,
   output        cfg_en2310,
   output        cfg_en2311,
   output        cfg_en2312,
   output        cfg_en2313,
   output        cfg_en2314,
   output        cfg_en2315,
   output        cfg_en2316,
   output        cfg_en2317,
   output        cfg_en2318,
   output        cfg_en2319,
   output        cfg_en2320,
   output        cfg_en2321,
   output        cfg_en2322,
   output        cfg_en2323,
   output        cfg_en2324,
   output        cfg_en2325,
   output        cfg_en2326,
   output        cfg_en2327,
   output        cfg_en2328,
   output        cfg_en2329,
   output        cfg_en2330,
   output        cfg_en2331,
   output        cfg_en2332,
   output        cfg_en2333,
   output        cfg_en2334,
   output        cfg_en2335,
   output        cfg_en2336,
   output        cfg_en2337,
   output        cfg_en2338,
   output        cfg_en2339,
   output        cfg_en2340,
   output        cfg_en2341,
   output        cfg_en2342,
   output        cfg_en2343,
   output        cfg_en2344,
   output        cfg_en2345,
   output        cfg_en2346,
   output        cfg_en2347,
   output        cfg_en2348,
   output        cfg_en2349,
   output        cfg_en2350,
   output        cfg_en2351,
   output        cfg_en2352,
   output        cfg_en2353,
   output        cfg_en2354,
   output        cfg_en2355,
   output        cfg_en2356,
   output        cfg_en2357,
   output        cfg_en2358,
   output        cfg_en2359,
   output        cfg_en2360,
   output        cfg_en2361,
   output        cfg_en2362,
   output        cfg_en2363,
   output        cfg_en2364,
   output        cfg_en2365,
   output        cfg_en2366,
   output        cfg_en2367,
   output        cfg_en2368,
   output        cfg_en2369,
   output        cfg_en2370,
   output        cfg_en2371,
   output        cfg_en2372,
   output        cfg_en2373,
   output        cfg_en2374,
   output        cfg_en2375,
   output        cfg_en2376,
   output        cfg_en2377,
   output        cfg_en2378,
   output        cfg_en2379,
   output        cfg_en2380,
   output        cfg_en2381,
   output        cfg_en2382,
   output        cfg_en2383,
   output        cfg_en2384,
   output        cfg_en2385,
   output        cfg_en2386,
   output        cfg_en2387,
   output        cfg_en2388,
   output        cfg_en2389,
   output        cfg_en2390,
   output        cfg_en2391,
   output        cfg_en2392,
   output        cfg_en2393,
   output        cfg_en2394,
   output        cfg_en2395,
   output        cfg_en2396,
   output        cfg_en2397,
   output        cfg_en2398,
   output        cfg_en2399,
   output        cfg_en2400,
   output        cfg_en2401,
   output        cfg_en2402,
   output        cfg_en2403,
   output        cfg_en2404,
   output        cfg_en2405,
   output        cfg_en2406,
   output        cfg_en2407,
   output        cfg_en2408,
   output        cfg_en2409,
   output        cfg_en2410,
   output        cfg_en2411,
   output        cfg_en2412,
   output        cfg_en2413,
   output        cfg_en2414,
   output        cfg_en2415,
   output        cfg_en2416,
   output        cfg_en2417,
   output        cfg_en2418,
   output        cfg_en2419,
   output        cfg_en2420,
   output        cfg_en2421,
   output        cfg_en2422,
   output        cfg_en2423,
   output        cfg_en2424,
   output        cfg_en2425,
   output        cfg_en2426,
   output        cfg_en2427,
   output        cfg_en2428,
   output        cfg_en2429,
   output        cfg_en2430,
   output        cfg_en2431,
   output        cfg_en2432,
   output        cfg_en2433,
   output        cfg_en2434,
   output        cfg_en2435,
   output        cfg_en2436,
   output        cfg_en2437,
   output        cfg_en2438,
   output        cfg_en2439,
   output        cfg_en2440,
   output        cfg_en2441,
   output        cfg_en2442,
   output        cfg_en2443,
   output        cfg_en2444,
   output        cfg_en2445,
   output        cfg_en2446,
   output        cfg_en2447,
   output        cfg_en2448,
   output        cfg_en2449,
   output        cfg_en2450,
   output        cfg_en2451,
   output        cfg_en2452,
   output        cfg_en2453,
   output        cfg_en2454,
   output        cfg_en2455,
   output        cfg_en2456,
   output        cfg_en2457,
   output        cfg_en2458,
   output        cfg_en2459,
   output        cfg_en2460,
   output        cfg_en2461,
   output        cfg_en2462,
   output        cfg_en2463,
   output        cfg_en2464,
   output        cfg_en2465,
   output        cfg_en2466,
   output        cfg_en2467,
   output        cfg_en2468,
   output        cfg_en2469,
   output        cfg_en2470,
   output        cfg_en2471,
   output        cfg_en2472,
   output        cfg_en2473,
   output        cfg_en2474,
   output        cfg_en2475,
   output        cfg_en2476,
   output        cfg_en2477,
   output        cfg_en2478,
   output        cfg_en2479,
   output        cfg_en2480,
   output        cfg_en2481,
   output        cfg_en2482,
   output        cfg_en2483,
   output        cfg_en2484,
   output        cfg_en2485,
   output        cfg_en2486,
   output        cfg_en2487,
   output        cfg_en2488,
   output        cfg_en2489,
   output        cfg_en2490,
   output        cfg_en2491,
   output        cfg_en2492,
   output        cfg_en2493,
   output        cfg_en2494,
   output        cfg_en2495,
   output        cfg_en2496,
   output        cfg_en2497,
   output        cfg_en2498,
   output        cfg_en2499,
   output        cfg_en2500,
   output        cfg_en2501,
   output        cfg_en2502,
   output        cfg_en2503,
   output        cfg_en2504,
   output        cfg_en2505,
   output        cfg_en2506,
   output        cfg_en2507,
   output        cfg_en2508,
   output        cfg_en2509,
   output        cfg_en2510,
   output        cfg_en2511,
   output        cfg_en2512,
   output        cfg_en2513,
   output        cfg_en2514,
   output        cfg_en2515,
   output        cfg_en2516,
   output        cfg_en2517,
   output        cfg_en2518,
   output        cfg_en2519,
   output        cfg_en2520,
   output        cfg_en2521,
   output        cfg_en2522,
   output        cfg_en2523,
   output        cfg_en2524,
   output        cfg_en2525,
   output        cfg_en2526,
   output        cfg_en2527,
   output        cfg_en2528,
   output        cfg_en2529,
   output        cfg_en2530,
   output        cfg_en2531,
   output        cfg_en2532,
   output        cfg_en2533,
   output        cfg_en2534,
   output        cfg_en2535,
   output        cfg_en2536,
   output        cfg_en2537,
   output        cfg_en2538,
   output        cfg_en2539,
   output        cfg_en2540,
   output        cfg_en2541,
   output        cfg_en2542,
   output        cfg_en2543,
   output        cfg_en2544,
   output        cfg_en2545,
   output        cfg_en2546,
   output        cfg_en2547,
   output        cfg_en2548,
   output        cfg_en2549,
   output        cfg_en2550,
   output        cfg_en2551,
   output        cfg_en2552,
   output        cfg_en2553,
   output        cfg_en2554,
   output        cfg_en2555,
   output        cfg_en2556,
   output        cfg_en2557,
   output        cfg_en2558,
   output        cfg_en2559,
   output        cfg_en2560,
   output        cfg_en2561,
   output        cfg_en2562,
   output        cfg_en2563,
   output        cfg_en2564,
   output        cfg_en2565,
   output        cfg_en2566,
   output        cfg_en2567,
   output        cfg_en2568,
   output        cfg_en2569,
   output        cfg_en2570,
   output        cfg_en2571,
   output        cfg_en2572,
   output        cfg_en2573,
   output        cfg_en2574,
   output        cfg_en2575,
   output        cfg_en2576,
   output        cfg_en2577,
   output        cfg_en2578,
   output        cfg_en2579,
   output        cfg_en2580,
   output        cfg_en2581,
   output        cfg_en2582,
   output        cfg_en2583,
   output        cfg_en2584,
   output        cfg_en2585,
   output        cfg_en2586,
   output        cfg_en2587,
   output        cfg_en2588,
   output        cfg_en2589,
   output        cfg_en2590,
   output        cfg_en2591,
   output        cfg_en2592,
   output        cfg_en2593,
   output        cfg_en2594,
   output        cfg_en2595,
   output        cfg_en2596,
   output        cfg_en2597,
   output        cfg_en2598,
   output        cfg_en2599,
   output        cfg_en2600,
   output        cfg_en2601,
   output        cfg_en2602,
   output        cfg_en2603,
   output        cfg_en2604,
   output        cfg_en2605,
   output        cfg_en2606,
   output        cfg_en2607,
   output        cfg_en2608,
   output        cfg_en2609,
   output        cfg_en2610,
   output        cfg_en2611,
   output        cfg_en2612,
   output        cfg_en2613,
   output        cfg_en2614,
   output        cfg_en2615,
   output        cfg_en2616,
   output        cfg_en2617,
   output        cfg_en2618,
   output        cfg_en2619,
   output        cfg_en2620,
   output        cfg_en2621,
   output        cfg_en2622,
   output        cfg_en2623,
   output        cfg_en2624,
   output        cfg_en2625,
   output        cfg_en2626,
   output        cfg_en2627,
   output        cfg_en2628,
   output        cfg_en2629,
   output        cfg_en2630,
   output        cfg_en2631,
   output        cfg_en2632,
   output        cfg_en2633,
   output        cfg_en2634,
   output        cfg_en2635,
   output        cfg_en2636,
   output        cfg_en2637,
   output        cfg_en2638,
   output        cfg_en2639,
   output        cfg_en2640,
   output        cfg_en2641,
   output        cfg_en2642,
   output        cfg_en2643,
   output        cfg_en2644,
   output        cfg_en2645,
   output        cfg_en2646,
   output        cfg_en2647,
   output        cfg_en2648,
   output        cfg_en2649,
   output        cfg_en2650,
   output        cfg_en2651,
   output        cfg_en2652,
   output        cfg_en2653,
   output        cfg_en2654,
   output        cfg_en2655,
   output        cfg_en2656,
   output        cfg_en2657,
   output        cfg_en2658,
   output        cfg_en2659,
   output        cfg_en2660,
   output        cfg_en2661,
   output        cfg_en2662,
   output        cfg_en2663,
   output        cfg_en2664,
   output        cfg_en2665,
   output        cfg_en2666,
   output        cfg_en2667,
   output        cfg_en2668,
   output        cfg_en2669,
   output        cfg_en2670,
   output        cfg_en2671,
   output        cfg_en2672,
   output        cfg_en2673,
   output        cfg_en2674,
   output        cfg_en2675,
   output        cfg_en2676,
   output        cfg_en2677,
   output        cfg_en2678,
   output        cfg_en2679,
   output        cfg_en2680,
   output        cfg_en2681,
   output        cfg_en2682,
   output        cfg_en2683,
   output        cfg_en2684,
   output        cfg_en2685,
   output        cfg_en2686,
   output        cfg_en2687,
   output        cfg_en2688,
   output        cfg_en2689,
   output        cfg_en2690,
   output        cfg_en2691,
   output        cfg_en2692,
   output        cfg_en2693,
   output        cfg_en2694,
   output        cfg_en2695,
   output        cfg_en2696,
   output        cfg_en2697,
   output        cfg_en2698,
   output        cfg_en2699,
   output        cfg_en2700,
   output        cfg_en2701,
   output        cfg_en2702,
   output        cfg_en2703,
   output        cfg_en2704,
   output        cfg_en2705,
   output        cfg_en2706,
   output        cfg_en2707,
   output        cfg_en2708,
   output        cfg_en2709,
   output        cfg_en2710,
   output        cfg_en2711,
   output        cfg_en2712,
   output        cfg_en2713,
   output        cfg_en2714,
   output        cfg_en2715,
   output        cfg_en2716,
   output        cfg_en2717,
   output        cfg_en2718,
   output        cfg_en2719,
   output        cfg_en2720,
   output        cfg_en2721,
   output        cfg_en2722,
   output        cfg_en2723,
   output        cfg_en2724,
   output        cfg_en2725,
   output        cfg_en2726,
   output        cfg_en2727,
   output        cfg_en2728,
   output        cfg_en2729,
   output        cfg_en2730,
   output        cfg_en2731,
   output        cfg_en2732,
   output        cfg_en2733,
   output        cfg_en2734,
   output        cfg_en2735,
   output        cfg_en2736,
   output        cfg_en2737,
   output        cfg_en2738,
   output        cfg_en2739,
   output        cfg_en2740,
   output        cfg_en2741,
   output        cfg_en2742,
   output        cfg_en2743,
   output        cfg_en2744,
   output        cfg_en2745,
   output        cfg_en2746,
   output        cfg_en2747,
   output        cfg_en2748,
   output        cfg_en2749,
   output        cfg_en2750,
   output        cfg_en2751,
   output        cfg_en2752,
   output        cfg_en2753,
   output        cfg_en2754,
   output        cfg_en2755,
   output        cfg_en2756,
   output        cfg_en2757,
   output        cfg_en2758,
   output        cfg_en2759,
   output        cfg_en2760,
   output        cfg_en2761,
   output        cfg_en2762,
   output        cfg_en2763,
   output        cfg_en2764,
   output        cfg_en2765,
   output        cfg_en2766,
   output        cfg_en2767,
   output        cfg_en2768,
   output        cfg_en2769,
   output        cfg_en2770,
   output        cfg_en2771,
   output        cfg_en2772,
   output        cfg_en2773,
   output        cfg_en2774,
   output        cfg_en2775,
   output        cfg_en2776,
   output        cfg_en2777,
   output        cfg_en2778,
   output        cfg_en2779,
   output        cfg_en2780,
   output        cfg_en2781,
   output        cfg_en2782,
   output        cfg_en2783,
   output        cfg_en2784,
   output        cfg_en2785,
   output        cfg_en2786,
   output        cfg_en2787,
   output        cfg_en2788,
   output        cfg_en2789,
   output        cfg_en2790,
   output        cfg_en2791,
   output        cfg_en2792,
   output        cfg_en2793,
   output        cfg_en2794,
   output        cfg_en2795,
   output        cfg_en2796,
   output        cfg_en2797,
   output        cfg_en2798,
   output        cfg_en2799,
   output        cfg_en2800,
   output        cfg_en2801,
   output        cfg_en2802,
   output        cfg_en2803,
   output        cfg_en2804,
   output        cfg_en2805,
   output        cfg_en2806,
   output        cfg_en2807,
   output        cfg_en2808,
   output        cfg_en2809,
   output        cfg_en2810,
   output        cfg_en2811,
   output        cfg_en2812,
   output        cfg_en2813,
   output        cfg_en2814,
   output        cfg_en2815,
   output        cfg_en2816,
   output        cfg_en2817,
   output        cfg_en2818,
   output        cfg_en2819,
   output        cfg_en2820,
   output        cfg_en2821,
   output        cfg_en2822,
   output        cfg_en2823,
   output        cfg_en2824,
   output        cfg_en2825,
   output        cfg_en2826,
   output        cfg_en2827,
   output        cfg_en2828,
   output        cfg_en2829,
   output        cfg_en2830,
   output        cfg_en2831,
   output        cfg_en2832,
   output        cfg_en2833,
   output        cfg_en2834,
   output        cfg_en2835,
   output        cfg_en2836,
   output        cfg_en2837,
   output        cfg_en2838,
   output        cfg_en2839,
   output        cfg_en2840,
   output        cfg_en2841,
   output        cfg_en2842,
   output        cfg_en2843,
   output        cfg_en2844,
   output        cfg_en2845,
   output        cfg_en2846,
   output        cfg_en2847,
   output        cfg_en2848,
   output        cfg_en2849,
   output        cfg_en2850,
   output        cfg_en2851,
   output        cfg_en2852,
   output        cfg_en2853,
   output        cfg_en2854,
   output        cfg_en2855,
   output        cfg_en2856,
   output        cfg_en2857,
   output        cfg_en2858,
   output        cfg_en2859,
   output        cfg_en2860,
   output        cfg_en2861,
   output        cfg_en2862,
   output        cfg_en2863,
   output        cfg_en2864,
   output        cfg_en2865,
   output        cfg_en2866,
   output        cfg_en2867,
   output        cfg_en2868,
   output        cfg_en2869,
   output        cfg_en2870,
   output        cfg_en2871,
   output        cfg_en2872,
   output        cfg_en2873,
   output        cfg_en2874,
   output        cfg_en2875,
   output        cfg_en2876,
   output        cfg_en2877,
   output        cfg_en2878,
   output        cfg_en2879,
   output        cfg_en2880,
   output        cfg_en2881,
   output        cfg_en2882,
   output        cfg_en2883,
   output        cfg_en2884,
   output        cfg_en2885,
   output        cfg_en2886,
   output        cfg_en2887,
   output        cfg_en2888,
   output        cfg_en2889,
   output        cfg_en2890,
   output        cfg_en2891,
   output        cfg_en2892,
   output        cfg_en2893,
   output        cfg_en2894,
   output        cfg_en2895,
   output        cfg_en2896,
   output        cfg_en2897,
   output        cfg_en2898,
   output        cfg_en2899,
   output        cfg_en2900,
   output        cfg_en2901,
   output        cfg_en2902,
   output        cfg_en2903,
   output        cfg_en2904,
   output        cfg_en2905,
   output        cfg_en2906,
   output        cfg_en2907,
   output        cfg_en2908,
   output        cfg_en2909,
   output        cfg_en2910,
   output        cfg_en2911,
   output        cfg_en2912,
   output        cfg_en2913,
   output        cfg_en2914,
   output        cfg_en2915,
   output        cfg_en2916,
   output        cfg_en2917,
   output        cfg_en2918,
   output        cfg_en2919,
   output        cfg_en2920,
   output        cfg_en2921,
   output        cfg_en2922,
   output        cfg_en2923,
   output        cfg_en2924,
   output        cfg_en2925,
   output        cfg_en2926,
   output        cfg_en2927,
   output        cfg_en2928,
   output        cfg_en2929,
   output        cfg_en2930,
   output        cfg_en2931,
   output        cfg_en2932,
   output        cfg_en2933,
   output        cfg_en2934,
   output        cfg_en2935,
   output        cfg_en2936,
   output        cfg_en2937,
   output        cfg_en2938,
   output        cfg_en2939,
   output        cfg_en2940,
   output        cfg_en2941,
   output        cfg_en2942,
   output        cfg_en2943,
   output        cfg_en2944,
   output        cfg_en2945,
   output        cfg_en2946,
   output        cfg_en2947,
   output        cfg_en2948,
   output        cfg_en2949,
   output        cfg_en2950,
   output        cfg_en2951,
   output        cfg_en2952,
   output        cfg_en2953,
   output        cfg_en2954,
   output        cfg_en2955,
   output        cfg_en2956,
   output        cfg_en2957,
   output        cfg_en2958,
   output        cfg_en2959,
   output        cfg_en2960,
   output        cfg_en2961,
   output        cfg_en2962,
   output        cfg_en2963,
   output        cfg_en2964,
   output        cfg_en2965,
   output        cfg_en2966,
   output        cfg_en2967,
   output        cfg_en2968,
   output        cfg_en2969,
   output        cfg_en2970,
   output        cfg_en2971,
   output        cfg_en2972,
   output        cfg_en2973,
   output        cfg_en2974,
   output        cfg_en2975,
   output        cfg_en2976,
   output        cfg_en2977,
   output        cfg_en2978,
   output        cfg_en2979,
   output        cfg_en2980,
   output        cfg_en2981,
   output        cfg_en2982,
   output        cfg_en2983,
   output        cfg_en2984,
   output        cfg_en2985,
   output        cfg_en2986,
   output        cfg_en2987,
   output        cfg_en2988,
   output        cfg_en2989,
   output        cfg_en2990,
   output        cfg_en2991,
   output        cfg_en2992,
   output        cfg_en2993,
   output        cfg_en2994,
   output        cfg_en2995,
   output        cfg_en2996,
   output        cfg_en2997,
   output        cfg_en2998,
   output        cfg_en2999,
   output        cfg_en3000,
   output        cfg_en3001,
   output        cfg_en3002,
   output        cfg_en3003,
   output        cfg_en3004,
   output        cfg_en3005,
   output        cfg_en3006,
   output        cfg_en3007,
   output        cfg_en3008,
   output        cfg_en3009,
   output        cfg_en3010,
   output        cfg_en3011,
   output        cfg_en3012,
   output        cfg_en3013,
   output        cfg_en3014,
   output        cfg_en3015,
   output        cfg_en3016,
   output        cfg_en3017,
   output        cfg_en3018,
   output        cfg_en3019,
   output        cfg_en3020,
   output        cfg_en3021,
   output        cfg_en3022,
   output        cfg_en3023,
   output        cfg_en3024,
   output        cfg_en3025,
   output        cfg_en3026,
   output        cfg_en3027,
   output        cfg_en3028,
   output        cfg_en3029,
   output        cfg_en3030,
   output        cfg_en3031,
   output        cfg_en3032,
   output        cfg_en3033,
   output        cfg_en3034,
   output        cfg_en3035,
   output        cfg_en3036,
   output        cfg_en3037,
   output        cfg_en3038,
   output        cfg_en3039,
   output        cfg_en3040,
   output        cfg_en3041,
   output        cfg_en3042,
   output        cfg_en3043,
   output        cfg_en3044,
   output        cfg_en3045,
   output        cfg_en3046,
   output        cfg_en3047,
   output        cfg_en3048,
   output        cfg_en3049,
   output        cfg_en3050,
   output        cfg_en3051,
   output        cfg_en3052,
   output        cfg_en3053,
   output        cfg_en3054,
   output        cfg_en3055,
   output        cfg_en3056,
   output        cfg_en3057,
   output        cfg_en3058,
   output        cfg_en3059,
   output        cfg_en3060,
   output        cfg_en3061,
   output        cfg_en3062,
   output        cfg_en3063,
   output        cfg_en3064,
   output        cfg_en3065,
   output        cfg_en3066,
   output        cfg_en3067,
   output        cfg_en3068,
   output        cfg_en3069,
   output        cfg_en3070,
   output        cfg_en3071,
   output        cfg_en3072,
   output        cfg_en3073,
   output        cfg_en3074,
   output        cfg_en3075,
   output        cfg_en3076,
   output        cfg_en3077,
   output        cfg_en3078,
   output        cfg_en3079,
   output        cfg_en3080,
   output        cfg_en3081,
   output        cfg_en3082,
   output        cfg_en3083,
   output        cfg_en3084,
   output        cfg_en3085,
   output        cfg_en3086,
   output        cfg_en3087,
   output        cfg_en3088,
   output        cfg_en3089,
   output        cfg_en3090,
   output        cfg_en3091,
   output        cfg_en3092,
   output        cfg_en3093,
   output        cfg_en3094,
   output        cfg_en3095,
   output        cfg_en3096,
   output        cfg_en3097,
   output        cfg_en3098,
   output        cfg_en3099,
   output        cfg_en3100,
   output        cfg_en3101,
   output        cfg_en3102,
   output        cfg_en3103,
   output        cfg_en3104,
   output        cfg_en3105,
   output        cfg_en3106,
   output        cfg_en3107,
   output        cfg_en3108,
   output        cfg_en3109,
   output        cfg_en3110,
   output        cfg_en3111,
   output        cfg_en3112,
   output        cfg_en3113,
   output        cfg_en3114,
   output        cfg_en3115,
   output        cfg_en3116,
   output        cfg_en3117,
   output        cfg_en3118,
   output        cfg_en3119,
   output        cfg_en3120,
   output        cfg_en3121,
   output        cfg_en3122,
   output        cfg_en3123,
   output        cfg_en3124,
   output        cfg_en3125,
   output        cfg_en3126,
   output        cfg_en3127,
   output        cfg_en3128,
   output        cfg_en3129,
   output        cfg_en3130,
   output        cfg_en3131,
   output        cfg_en3132,
   output        cfg_en3133,
   output        cfg_en3134,
   output        cfg_en3135,
   output        cfg_en3136,
   output        cfg_en3137,
   output        cfg_en3138,
   output        cfg_en3139,
   output        cfg_en3140,
   output        cfg_en3141,
   output        cfg_en3142,
   output        cfg_en3143,
   output        cfg_en3144,
   output        cfg_en3145,
   output        cfg_en3146,
   output        cfg_en3147,
   output        cfg_en3148,
   output        cfg_en3149,
   output        cfg_en3150,
   output        cfg_en3151,
   output        cfg_en3152,
   output        cfg_en3153,
   output        cfg_en3154,
   output        cfg_en3155,
   output        cfg_en3156,
   output        cfg_en3157,
   output        cfg_en3158,
   output        cfg_en3159,
   output        cfg_en3160,
   output        cfg_en3161,
   output        cfg_en3162,
   output        cfg_en3163,
   output        cfg_en3164,
   output        cfg_en3165,
   output        cfg_en3166,
   output        cfg_en3167,
   output        cfg_en3168,
   output        cfg_en3169,
   output        cfg_en3170,
   output        cfg_en3171,
   output        cfg_en3172,
   output        cfg_en3173,
   output        cfg_en3174,
   output        cfg_en3175,
   output        cfg_en3176,
   output        cfg_en3177,
   output        cfg_en3178,
   output        cfg_en3179,
   output        cfg_en3180,
   output        cfg_en3181,
   output        cfg_en3182,
   output        cfg_en3183,
   output        cfg_en3184,
   output        cfg_en3185,
   output        cfg_en3186,
   output        cfg_en3187,
   output        cfg_en3188,
   output        cfg_en3189,
   output        cfg_en3190,
   output        cfg_en3191,
   output        cfg_en3192,
   output        cfg_en3193,
   output        cfg_en3194,
   output        cfg_en3195,
   output        cfg_en3196,
   output        cfg_en3197,
   output        cfg_en3198,
   output        cfg_en3199,
   output        cfg_en3200,
   output        cfg_en3201,
   output        cfg_en3202,
   output        cfg_en3203,
   output        cfg_en3204,
   output        cfg_en3205,
   output        cfg_en3206,
   output        cfg_en3207,
   output        cfg_en3208,
   output        cfg_en3209,
   output        cfg_en3210,
   output        cfg_en3211,
   output        cfg_en3212,
   output        cfg_en3213,
   output        cfg_en3214,
   output        cfg_en3215,
   output        cfg_en3216,
   output        cfg_en3217,
   output        cfg_en3218,
   output        cfg_en3219,
   output        cfg_en3220,
   output        cfg_en3221,
   output        cfg_en3222,
   output        cfg_en3223,
   output        cfg_en3224,
   output        cfg_en3225,
   output        cfg_en3226,
   output        cfg_en3227,
   output        cfg_en3228,
   output        cfg_en3229,
   output        cfg_en3230,
   output        cfg_en3231,
   output        cfg_en3232,
   output        cfg_en3233,
   output        cfg_en3234,
   output        cfg_en3235,
   output        cfg_en3236,
   output        cfg_en3237,
   output        cfg_en3238,
   output        cfg_en3239,
   output        cfg_en3240,
   output        cfg_en3241,
   output        cfg_en3242,
   output        cfg_en3243,
   output        cfg_en3244,
   output        cfg_en3245,
   output        cfg_en3246,
   output        cfg_en3247,
   output        cfg_en3248,
   output        cfg_en3249,
   output        cfg_en3250,
   output        cfg_en3251,
   output        cfg_en3252,
   output        cfg_en3253,
   output        cfg_en3254,
   output        cfg_en3255,
   output        cfg_en3256,
   output        cfg_en3257,
   output        cfg_en3258,
   output        cfg_en3259,
   output        cfg_en3260,
   output        cfg_en3261,
   output        cfg_en3262,
   output        cfg_en3263,
   output        cfg_en3264,
   output        cfg_en3265,
   output        cfg_en3266,
   output        cfg_en3267,
   output        cfg_en3268,
   output        cfg_en3269,
   output        cfg_en3270,
   output        cfg_en3271,
   output        cfg_en3272,
   output        cfg_en3273,
   output        cfg_en3274,
   output        cfg_en3275,
   output        cfg_en3276,
   output        cfg_en3277,
   output        cfg_en3278,
   output        cfg_en3279,
   output        cfg_en3280,
   output        cfg_en3281,
   output        cfg_en3282,
   output        cfg_en3283,
   output        cfg_en3284,
   output        cfg_en3285,
   output        cfg_en3286,
   output        cfg_en3287,
   output        cfg_en3288,
   output        cfg_en3289,
   output        cfg_en3290,
   output        cfg_en3291,
   output        cfg_en3292,
   output        cfg_en3293,
   output        cfg_en3294,
   output        cfg_en3295,
   output        cfg_en3296,
   output        cfg_en3297,
   output        cfg_en3298,
   output        cfg_en3299,
   output        cfg_en3300,
   output        cfg_en3301,
   output        cfg_en3302,
   output        cfg_en3303,
   output        cfg_en3304,
   output        cfg_en3305,
   output        cfg_en3306,
   output        cfg_en3307,
   output        cfg_en3308,
   output        cfg_en3309,
   output        cfg_en3310,
   output        cfg_en3311,
   output        cfg_en3312,
   output        cfg_en3313,
   output        cfg_en3314,
   output        cfg_en3315,
   output        cfg_en3316,
   output        cfg_en3317,
   output        cfg_en3318,
   output        cfg_en3319,
   output        cfg_en3320,
   output        cfg_en3321,
   output        cfg_en3322,
   output        cfg_en3323,
   output        cfg_en3324,
   output        cfg_en3325,
   output        cfg_en3326,
   output        cfg_en3327,
   output        cfg_en3328,
   output        cfg_en3329,
   output        cfg_en3330,
   output        cfg_en3331,
   output        cfg_en3332,
   output        cfg_en3333,
   output        cfg_en3334,
   output        cfg_en3335,
   output        cfg_en3336,
   output        cfg_en3337,
   output        cfg_en3338,
   output        cfg_en3339,
   output        cfg_en3340,
   output        cfg_en3341,
   output        cfg_en3342,
   output        cfg_en3343,
   output        cfg_en3344,
   output        cfg_en3345,
   output        cfg_en3346,
   output        cfg_en3347,
   output        cfg_en3348,
   output        cfg_en3349,
   output        cfg_en3350,
   output        cfg_en3351,
   output        cfg_en3352,
   output        cfg_en3353,
   output        cfg_en3354,
   output        cfg_en3355,
   output        cfg_en3356,
   output        cfg_en3357,
   output        cfg_en3358,
   output        cfg_en3359,
   output        cfg_en3360,
   output        cfg_en3361,
   output        cfg_en3362,
   output        cfg_en3363,
   output        cfg_en3364,
   output        cfg_en3365,
   output        cfg_en3366,
   output        cfg_en3367,
   output        cfg_en3368,
   output        cfg_en3369,
   output        cfg_en3370,
   output        cfg_en3371,
   output        cfg_en3372,
   output        cfg_en3373,
   output        cfg_en3374,
   output        cfg_en3375,
   output        cfg_en3376,
   output        cfg_en3377,
   output        cfg_en3378,
   output        cfg_en3379,
   output        cfg_en3380,
   output        cfg_en3381,
   output        cfg_en3382,
   output        cfg_en3383,
   output        cfg_en3384,
   output        cfg_en3385,
   output        cfg_en3386,
   output        cfg_en3387,
   output        cfg_en3388,
   output        cfg_en3389,
   output        cfg_en3390,
   output        cfg_en3391,
   output        cfg_en3392,
   output        cfg_en3393,
   output        cfg_en3394,
   output        cfg_en3395,
   output        cfg_en3396,
   output        cfg_en3397,
   output        cfg_en3398,
   output        cfg_en3399,
   output        cfg_en3400,
   output        cfg_en3401,
   output        cfg_en3402,
   output        cfg_en3403,
   output        cfg_en3404,
   output        cfg_en3405,
   output        cfg_en3406,
   output        cfg_en3407,
   output        cfg_en3408,
   output        cfg_en3409,
   output        cfg_en3410,
   output        cfg_en3411,
   output        cfg_en3412,
   output        cfg_en3413,
   output        cfg_en3414,
   output        cfg_en3415,
   output        cfg_en3416,
   output        cfg_en3417,
   output        cfg_en3418,
   output        cfg_en3419,
   output        cfg_en3420,
   output        cfg_en3421,
   output        cfg_en3422,
   output        cfg_en3423,
   output        cfg_en3424,
   output        cfg_en3425,
   output        cfg_en3426,
   output        cfg_en3427,
   output        cfg_en3428,
   output        cfg_en3429,
   output        cfg_en3430,
   output        cfg_en3431,
   output        cfg_en3432,
   output        cfg_en3433,
   output        cfg_en3434,
   output        cfg_en3435,
   output        cfg_en3436,
   output        cfg_en3437,
   output        cfg_en3438,
   output        cfg_en3439,
   output        cfg_en3440,
   output        cfg_en3441,
   output        cfg_en3442,
   output        cfg_en3443,
   output        cfg_en3444,
   output        cfg_en3445,
   output        cfg_en3446,
   output        cfg_en3447,
   output        cfg_en3448,
   output        cfg_en3449,
   output        cfg_en3450,
   output        cfg_en3451,
   output        cfg_en3452,
   output        cfg_en3453,
   output        cfg_en3454,
   output        cfg_en3455,
   output        cfg_en3456,
   output        cfg_en3457,
   output        cfg_en3458,
   output        cfg_en3459,
   output        cfg_en3460,
   output        cfg_en3461,
   output        cfg_en3462,
   output        cfg_en3463,
   output        cfg_en3464,
   output        cfg_en3465,
   output        cfg_en3466,
   output        cfg_en3467,
   output        cfg_en3468,
   output        cfg_en3469,
   output        cfg_en3470,
   output        cfg_en3471,
   output        cfg_en3472,
   output        cfg_en3473,
   output        cfg_en3474,
   output        cfg_en3475,
   output        cfg_en3476,
   output        cfg_en3477,
   output        cfg_en3478,
   output        cfg_en3479,
   output        cfg_en3480,
   output        cfg_en3481,
   output        cfg_en3482,
   output        cfg_en3483,
   output        cfg_en3484,
   output        cfg_en3485,
   output        cfg_en3486,
   output        cfg_en3487,
   output        cfg_en3488,
   output        cfg_en3489,
   output        cfg_en3490,
   output        cfg_en3491,
   output        cfg_en3492,
   output        cfg_en3493,
   output        cfg_en3494,
   output        cfg_en3495,
   output        cfg_en3496,
   output        cfg_en3497,
   output        cfg_en3498,
   output        cfg_en3499,
   output        cfg_en3500,
   output        cfg_en3501,
   output        cfg_en3502,
   output        cfg_en3503,
   output        cfg_en3504,
   output        cfg_en3505,
   output        cfg_en3506,
   output        cfg_en3507,
   output        cfg_en3508,
   output        cfg_en3509,
   output        cfg_en3510,
   output        cfg_en3511,
   output        cfg_en3512,
   output        cfg_en3513,
   output        cfg_en3514,
   output        cfg_en3515,
   output        cfg_en3516,
   output        cfg_en3517,
   output        cfg_en3518,
   output        cfg_en3519,
   output        cfg_en3520,
   output        cfg_en3521,
   output        cfg_en3522,
   output        cfg_en3523,
   output        cfg_en3524,
   output        cfg_en3525,
   output        cfg_en3526,
   output        cfg_en3527,
   output        cfg_en3528,
   output        cfg_en3529,
   output        cfg_en3530,
   output        cfg_en3531,
   output        cfg_en3532,
   output        cfg_en3533,
   output        cfg_en3534,
   output        cfg_en3535,
   output        cfg_en3536,
   output        cfg_en3537,
   output        cfg_en3538,
   output        cfg_en3539,
   output        cfg_en3540,
   output        cfg_en3541,
   output        cfg_en3542,
   output        cfg_en3543,
   output        cfg_en3544,
   output        cfg_en3545,
   output        cfg_en3546,
   output        cfg_en3547,
   output        cfg_en3548,
   output        cfg_en3549,
   output        cfg_en3550,
   output        cfg_en3551,
   output        cfg_en3552,
   output        cfg_en3553,
   output        cfg_en3554,
   output        cfg_en3555,
   output        cfg_en3556,
   output        cfg_en3557,
   output        cfg_en3558,
   output        cfg_en3559,
   output        cfg_en3560,
   output        cfg_en3561,
   output        cfg_en3562,
   output        cfg_en3563,
   output        cfg_en3564,
   output        cfg_en3565,
   output        cfg_en3566,
   output        cfg_en3567,
   output        cfg_en3568,
   output        cfg_en3569,
   output        cfg_en3570,
   output        cfg_en3571,
   output        cfg_en3572,
   output        cfg_en3573,
   output        cfg_en3574,
   output        cfg_en3575,
   output        cfg_en3576,
   output        cfg_en3577,
   output        cfg_en3578,
   output        cfg_en3579,
   output        cfg_en3580,
   output        cfg_en3581,
   output        cfg_en3582,
   output        cfg_en3583,
   output        cfg_en3584,
   output        cfg_en3585,
   output        cfg_en3586,
   output        cfg_en3587,
   output        cfg_en3588,
   output        cfg_en3589,
   output        cfg_en3590,
   output        cfg_en3591,
   output        cfg_en3592,
   output        cfg_en3593,
   output        cfg_en3594,
   output        cfg_en3595,
   output        cfg_en3596,
   output        cfg_en3597,
   output        cfg_en3598,
   output        cfg_en3599,
   output        cfg_en3600,
   output        cfg_en3601,
   output        cfg_en3602,
   output        cfg_en3603,
   output        cfg_en3604,
   output        cfg_en3605,
   output        cfg_en3606,
   output        cfg_en3607,
   output        cfg_en3608,
   output        cfg_en3609,
   output        cfg_en3610,
   output        cfg_en3611,
   output        cfg_en3612,
   output        cfg_en3613,
   output        cfg_en3614,
   output        cfg_en3615,
   output        cfg_en3616,
   output        cfg_en3617,
   output        cfg_en3618,
   output        cfg_en3619,
   output        cfg_en3620,
   output        cfg_en3621,
   output        cfg_en3622,
   output        cfg_en3623,
   output        cfg_en3624,
   output        cfg_en3625,
   output        cfg_en3626,
   output        cfg_en3627,
   output        cfg_en3628,
   output        cfg_en3629,
   output        cfg_en3630,
   output        cfg_en3631,
   output        cfg_en3632,
   output        cfg_en3633,
   output        cfg_en3634,
   output        cfg_en3635,
   output        cfg_en3636,
   output        cfg_en3637,
   output        cfg_en3638,
   output        cfg_en3639,
   output        cfg_en3640,
   output        cfg_en3641,
   output        cfg_en3642,
   output        cfg_en3643,
   output        cfg_en3644,
   output        cfg_en3645,
   output        cfg_en3646,
   output        cfg_en3647,
   output        cfg_en3648,
   output        cfg_en3649,
   output        cfg_en3650,
   output        cfg_en3651,
   output        cfg_en3652,
   output        cfg_en3653,
   output        cfg_en3654,
   output        cfg_en3655,
   output        cfg_en3656,
   output        cfg_en3657,
   output        cfg_en3658,
   output        cfg_en3659,
   output        cfg_en3660,
   output        cfg_en3661,
   output        cfg_en3662,
   output        cfg_en3663,
   output        cfg_en3664,
   output        cfg_en3665,
   output        cfg_en3666,
   output        cfg_en3667,
   output        cfg_en3668,
   output        cfg_en3669,
   output        cfg_en3670,
   output        cfg_en3671,
   output        cfg_en3672,
   output        cfg_en3673,
   output        cfg_en3674,
   output        cfg_en3675,
   output        cfg_en3676,
   output        cfg_en3677,
   output        cfg_en3678,
   output        cfg_en3679,
   output        cfg_en3680,
   output        cfg_en3681,
   output        cfg_en3682,
   output        cfg_en3683,
   output        cfg_en3684,
   output        cfg_en3685,
   output        cfg_en3686,
   output        cfg_en3687,
   output        cfg_en3688,
   output        cfg_en3689,
   output        cfg_en3690,
   output        cfg_en3691,
   output        cfg_en3692,
   output        cfg_en3693,
   output        cfg_en3694,
   output        cfg_en3695,
   output        cfg_en3696,
   output        cfg_en3697,
   output        cfg_en3698,
   output        cfg_en3699,
   output        cfg_en3700,
   output        cfg_en3701,
   output        cfg_en3702,
   output        cfg_en3703,
   output        cfg_en3704,
   output        cfg_en3705,
   output        cfg_en3706,
   output        cfg_en3707,
   output        cfg_en3708,
   output        cfg_en3709,
   output        cfg_en3710,
   output        cfg_en3711,
   output        cfg_en3712,
   output        cfg_en3713,
   output        cfg_en3714,
   output        cfg_en3715,
   output        cfg_en3716,
   output        cfg_en3717,
   output        cfg_en3718,
   output        cfg_en3719,
   output        cfg_en3720,
   output        cfg_en3721,
   output        cfg_en3722,
   output        cfg_en3723,
   output        cfg_en3724,
   output        cfg_en3725,
   output        cfg_en3726,
   output        cfg_en3727,
   output        cfg_en3728,
   output        cfg_en3729,
   output        cfg_en3730,
   output        cfg_en3731,
   output        cfg_en3732,
   output        cfg_en3733,
   output        cfg_en3734,
   output        cfg_en3735,
   output        cfg_en3736,
   output        cfg_en3737,
   output        cfg_en3738,
   output        cfg_en3739,
   output        cfg_en3740,
   output        cfg_en3741,
   output        cfg_en3742,
   output        cfg_en3743,
   output        cfg_en3744,
   output        cfg_en3745,
   output        cfg_en3746,
   output        cfg_en3747,
   output        cfg_en3748,
   output        cfg_en3749,
   output        cfg_en3750,
   output        cfg_en3751,
   output        cfg_en3752,
   output        cfg_en3753,
   output        cfg_en3754,
   output        cfg_en3755,
   output        cfg_en3756,
   output        cfg_en3757,
   output        cfg_en3758,
   output        cfg_en3759,
   output        cfg_en3760,
   output        cfg_en3761,
   output        cfg_en3762,
   output        cfg_en3763,
   output        cfg_en3764,
   output        cfg_en3765,
   output        cfg_en3766,
   output        cfg_en3767,
   output        cfg_en3768,
   output        cfg_en3769,
   output        cfg_en3770,
   output        cfg_en3771,
   output        cfg_en3772,
   output        cfg_en3773,
   output        cfg_en3774,
   output        cfg_en3775,
   output        cfg_en3776,
   output        cfg_en3777,
   output        cfg_en3778,
   output        cfg_en3779,
   output        cfg_en3780,
   output        cfg_en3781,
   output        cfg_en3782,
   output        cfg_en3783,
   output        cfg_en3784,
   output        cfg_en3785,
   output        cfg_en3786,
   output        cfg_en3787,
   output        cfg_en3788,
   output        cfg_en3789,
   output        cfg_en3790,
   output        cfg_en3791,
   output        cfg_en3792,
   output        cfg_en3793,
   output        cfg_en3794,
   output        cfg_en3795,
   output        cfg_en3796,
   output        cfg_en3797,
   output        cfg_en3798,
   output        cfg_en3799,
   output        cfg_en3800,
   output        cfg_en3801,
   output        cfg_en3802,
   output        cfg_en3803,
   output        cfg_en3804,
   output        cfg_en3805,
   output        cfg_en3806,
   output        cfg_en3807,
   output        cfg_en3808,
   output        cfg_en3809,
   output        cfg_en3810,
   output        cfg_en3811,
   output        cfg_en3812,
   output        cfg_en3813,
   output        cfg_en3814,
   output        cfg_en3815,
   output        cfg_en3816,
   output        cfg_en3817,
   output        cfg_en3818,
   output        cfg_en3819,
   output        cfg_en3820,
   output        cfg_en3821,
   output        cfg_en3822,
   output        cfg_en3823,
   output        cfg_en3824,
   output        cfg_en3825,
   output        cfg_en3826,
   output        cfg_en3827,
   output        cfg_en3828,
   output        cfg_en3829,
   output        cfg_en3830,
   output        cfg_en3831,
   output        cfg_en3832,
   output        cfg_en3833,
   output        cfg_en3834,
   output        cfg_en3835,
   output        cfg_en3836,
   output        cfg_en3837,
   output        cfg_en3838,
   output        cfg_en3839,
   output        cfg_en3840,
   output        cfg_en3841,
   output        cfg_en3842,
   output        cfg_en3843,
   output        cfg_en3844,
   output        cfg_en3845,
   output        cfg_en3846,
   output        cfg_en3847,
   output        cfg_en3848,
   output        cfg_en3849,
   output        cfg_en3850,
   output        cfg_en3851,
   output        cfg_en3852,
   output        cfg_en3853,
   output        cfg_en3854,
   output        cfg_en3855,
   output        cfg_en3856,
   output        cfg_en3857,
   output        cfg_en3858,
   output        cfg_en3859,
   output        cfg_en3860,
   output        cfg_en3861,
   output        cfg_en3862,
   output        cfg_en3863,
   output        cfg_en3864,
   output        cfg_en3865,
   output        cfg_en3866,
   output        cfg_en3867,
   output        cfg_en3868,
   output        cfg_en3869,
   output        cfg_en3870,
   output        cfg_en3871,
   output        cfg_en3872,
   output        cfg_en3873,
   output        cfg_en3874,
   output        cfg_en3875,
   output        cfg_en3876,
   output        cfg_en3877,
   output        cfg_en3878,
   output        cfg_en3879,
   output        cfg_en3880,
   output        cfg_en3881,
   output        cfg_en3882,
   output        cfg_en3883,
   output        cfg_en3884,
   output        cfg_en3885,
   output        cfg_en3886,
   output        cfg_en3887,
   output        cfg_en3888,
   output        cfg_en3889,
   output        cfg_en3890,
   output        cfg_en3891,
   output        cfg_en3892,
   output        cfg_en3893,
   output        cfg_en3894,
   output        cfg_en3895,
   output        cfg_en3896,
   output        cfg_en3897,
   output        cfg_en3898,
   output        cfg_en3899,
   output        cfg_en3900,
   output        cfg_en3901,
   output        cfg_en3902,
   output        cfg_en3903,
   output        cfg_en3904,
   output        cfg_en3905,
   output        cfg_en3906,
   output        cfg_en3907,
   output        cfg_en3908,
   output        cfg_en3909,
   output        cfg_en3910,
   output        cfg_en3911,
   output        cfg_en3912,
   output        cfg_en3913,
   output        cfg_en3914,
   output        cfg_en3915,
   output        cfg_en3916,
   output        cfg_en3917,
   output        cfg_en3918,
   output        cfg_en3919,
   output        cfg_en3920,
   output        cfg_en3921,
   output        cfg_en3922,
   output        cfg_en3923,
   output        cfg_en3924,
   output        cfg_en3925,
   output        cfg_en3926,
   output        cfg_en3927,
   output        cfg_en3928,
   output        cfg_en3929,
   output        cfg_en3930,
   output        cfg_en3931,
   output        cfg_en3932,
   output        cfg_en3933,
   output        cfg_en3934,
   output        cfg_en3935,
   output        cfg_en3936,
   output        cfg_en3937,
   output        cfg_en3938,
   output        cfg_en3939,
   output        cfg_en3940,
   output        cfg_en3941,
   output        cfg_en3942,
   output        cfg_en3943,
   output        cfg_en3944,
   output        cfg_en3945,
   output        cfg_en3946,
   output        cfg_en3947,
   output        cfg_en3948,
   output        cfg_en3949,
   output        cfg_en3950,
   output        cfg_en3951,
   output        cfg_en3952,
   output        cfg_en3953,
   output        cfg_en3954,
   output        cfg_en3955,
   output        cfg_en3956,
   output        cfg_en3957,
   output        cfg_en3958,
   output        cfg_en3959,
   output        cfg_en3960,
   output        cfg_en3961,
   output        cfg_en3962,
   output        cfg_en3963,
   output        cfg_en3964,
   output        cfg_en3965,
   output        cfg_en3966,
   output        cfg_en3967,
   output        cfg_en3968,
   output        cfg_en3969,
   output        cfg_en3970,
   output        cfg_en3971,
   output        cfg_en3972,
   output        cfg_en3973,
   output        cfg_en3974,
   output        cfg_en3975,
   output        cfg_en3976,
   output        cfg_en3977,
   output        cfg_en3978,
   output        cfg_en3979,
   output        cfg_en3980,
   output        cfg_en3981,
   output        cfg_en3982,
   output        cfg_en3983,
   output        cfg_en3984,
   output        cfg_en3985,
   output        cfg_en3986,
   output        cfg_en3987,
   output        cfg_en3988,
   output        cfg_en3989,
   output        cfg_en3990,
   output        cfg_en3991,
   output        cfg_en3992,
   output        cfg_en3993,
   output        cfg_en3994,
   output        cfg_en3995,
   output        cfg_en3996,
   output        cfg_en3997,
   output        cfg_en3998,
   output        cfg_en3999,
   output        cfg_en4000,
   output        cfg_en4001,
   output        cfg_en4002,
   output        cfg_en4003,
   output        cfg_en4004,
   output        cfg_en4005,
   output        cfg_en4006,
   output        cfg_en4007,
   output        cfg_en4008,
   output        cfg_en4009,
   output        cfg_en4010,
   output        cfg_en4011,
   output        cfg_en4012,
   output        cfg_en4013,
   output        cfg_en4014,
   output        cfg_en4015,
   output        cfg_en4016,
   output        cfg_en4017,
   output        cfg_en4018,
   output        cfg_en4019,
   output        cfg_en4020,
   output        cfg_en4021,
   output        cfg_en4022,
   output        cfg_en4023,
   output        cfg_en4024,
   output        cfg_en4025,
   output        cfg_en4026,
   output        cfg_en4027,
   output        cfg_en4028,
   output        cfg_en4029,
   output        cfg_en4030,
   output        cfg_en4031,
   output        cfg_en4032,
   output        cfg_en4033,
   output        cfg_en4034,
   output        cfg_en4035,
   output        cfg_en4036,
   output        cfg_en4037,
   output        cfg_en4038,
   output        cfg_en4039,
   output        cfg_en4040,
   output        cfg_en4041,
   output        cfg_en4042,
   output        cfg_en4043,
   output        cfg_en4044,
   output        cfg_en4045,
   output        cfg_en4046,
   output        cfg_en4047,
   output        cfg_en4048,
   output        cfg_en4049,
   output        cfg_en4050,
   output        cfg_en4051,
   output        cfg_en4052,
   output        cfg_en4053,
   output        cfg_en4054,
   output        cfg_en4055,
   output        cfg_en4056,
   output        cfg_en4057,
   output        cfg_en4058,
   output        cfg_en4059,
   output        cfg_en4060,
   output        cfg_en4061,
   output        cfg_en4062,
   output        cfg_en4063,
   output        cfg_en4064,
   output        cfg_en4065,
   output        cfg_en4066,
   output        cfg_en4067,
   output        cfg_en4068,
   output        cfg_en4069,
   output        cfg_en4070,
   output        cfg_en4071,
   output        cfg_en4072,
   output        cfg_en4073,
   output        cfg_en4074,
   output        cfg_en4075,
   output        cfg_en4076,
   output        cfg_en4077,
   output        cfg_en4078,
   output        cfg_en4079,
   output        cfg_en4080,
   output        cfg_en4081,
   output        cfg_en4082,
   output        cfg_en4083,
   output        cfg_en4084,
   output        cfg_en4085,
   output        cfg_en4086,
   output        cfg_en4087,
   output        cfg_en4088,
   output        cfg_en4089,
   output        cfg_en4090,
   output        cfg_en4091,
   output        cfg_en4092,
   output        cfg_en4093,
   output        cfg_en4094,
   output        cfg_en4095,
   output        cfg_en4096,
   output        cfg_en4097,
   output        cfg_en4098,
   output        cfg_en4099,
   output        cfg_en4100,
   output        cfg_en4101,
   output        cfg_en4102,
   output        cfg_en4103,
   output        cfg_en4104,
   output        cfg_en4105,
   output        cfg_en4106,
   output        cfg_en4107,
   output        cfg_en4108,
   output        cfg_en4109,
   output        cfg_en4110,
   output        cfg_en4111,
   output        cfg_en4112,
   output        cfg_en4113,
   output        cfg_en4114,
   output        cfg_en4115,
   output        cfg_en4116,
   output        cfg_en4117,
   output        cfg_en4118,
   output        cfg_en4119,
   output        cfg_en4120,
   output        cfg_en4121,
   output        cfg_en4122,
   output        cfg_en4123,
   output        cfg_en4124,
   output        cfg_en4125,
   output        cfg_en4126,
   output        cfg_en4127,
   output        cfg_en4128,
   output        cfg_en4129,
   output        cfg_en4130,
   output        cfg_en4131,
   output        cfg_en4132,
   output        cfg_en4133,
   output        cfg_en4134,
   output        cfg_en4135,
   output        cfg_en4136,
   output        cfg_en4137,
   output        cfg_en4138,
   output        cfg_en4139,
   output        cfg_en4140,
   output        cfg_en4141,
   output        cfg_en4142,
   output        cfg_en4143,
   output        cfg_en4144,
   output        cfg_en4145,
   output        cfg_en4146,
   output        cfg_en4147,
   output        cfg_en4148,
   output        cfg_en4149,
   output        cfg_en4150,
   output        cfg_en4151,
   output        cfg_en4152,
   output        cfg_en4153,
   output        cfg_en4154,
   output        cfg_en4155,
   output        cfg_en4156,
   output        cfg_en4157,
   output        cfg_en4158,
   output        cfg_en4159,
   output        cfg_en4160,
   output        cfg_en4161,
   output        cfg_en4162,
   output        cfg_en4163,
   output        cfg_en4164,
   output        cfg_en4165,
   output        cfg_en4166,
   output        cfg_en4167,
   output        cfg_en4168,
   output        cfg_en4169,
   output        cfg_en4170,
   output        cfg_en4171,
   output        cfg_en4172,
   output        cfg_en4173,
   output        cfg_en4174,
   output        cfg_en4175,
   output        cfg_en4176,
   output        cfg_en4177,
   output        cfg_en4178,
   output        cfg_en4179,
   output        cfg_en4180,
   output        cfg_en4181,
   output        cfg_en4182,
   output        cfg_en4183,
   output        cfg_en4184,
   output        cfg_en4185,
   output        cfg_en4186,
   output        cfg_en4187,
   output        cfg_en4188,
   output        cfg_en4189,
   output        cfg_en4190,
   output        cfg_en4191,
   output        cfg_en4192,
   output        cfg_en4193,
   output        cfg_en4194,
   output        cfg_en4195,
   output        cfg_en4196,
   output        cfg_en4197,
   output        cfg_en4198,
   output        cfg_en4199,
   output        cfg_en4200,
   output        cfg_en4201,
   output        cfg_en4202,
   output        cfg_en4203,
   output        cfg_en4204,
   output        cfg_en4205,
   output        cfg_en4206,
   output        cfg_en4207,
   output        cfg_en4208,
   output        cfg_en4209,
   output        cfg_en4210,
   output        cfg_en4211,
   output        cfg_en4212,
   output        cfg_en4213,
   output        cfg_en4214,
   output        cfg_en4215,
   output        cfg_en4216,
   output        cfg_en4217,
   output        cfg_en4218,
   output        cfg_en4219,
   output        cfg_en4220,
   output        cfg_en4221,
   output        cfg_en4222,
   output        cfg_en4223,
   output        cfg_en4224,
   output        cfg_en4225,
   output        cfg_en4226,
   output        cfg_en4227,
   output        cfg_en4228,
   output        cfg_en4229,
   output        cfg_en4230,
   output        cfg_en4231,
   output        cfg_en4232,
   output        cfg_en4233,
   output        cfg_en4234,
   output        cfg_en4235,
   output        cfg_en4236,
   output        cfg_en4237,
   output        cfg_en4238,
   output        cfg_en4239,
   output        cfg_en4240,
   output        cfg_en4241,
   output        cfg_en4242,
   output        cfg_en4243,
   output        cfg_en4244,
   output        cfg_en4245,
   output        cfg_en4246,
   output        cfg_en4247,
   output        cfg_en4248,
   output        cfg_en4249,
   output        cfg_en4250,
   output        cfg_en4251,
   output        cfg_en4252,
   output        cfg_en4253,
   output        cfg_en4254,
   output        cfg_en4255,
   output        cfg_en4256,
   output        cfg_en4257,
   output        cfg_en4258,
   output        cfg_en4259,
   output        cfg_en4260,
   output        cfg_en4261,
   output        cfg_en4262,
   output        cfg_en4263,
   output        cfg_en4264,
   output        cfg_en4265,
   output        cfg_en4266,
   output        cfg_en4267,
   output        cfg_en4268,
   output        cfg_en4269,
   output        cfg_en4270,
   output        cfg_en4271,
   output        cfg_en4272,
   output        cfg_en4273,
   output        cfg_en4274,
   output        cfg_en4275,
   output        cfg_en4276,
   output        cfg_en4277,
   output        cfg_en4278,
   output        cfg_en4279,
   output        cfg_en4280,
   output        cfg_en4281,
   output        cfg_en4282,
   output        cfg_en4283,
   output        cfg_en4284,
   output        cfg_en4285,
   output        cfg_en4286,
   output        cfg_en4287,
   output        cfg_en4288,
   output        cfg_en4289,
   output        cfg_en4290,
   output        cfg_en4291,
   output        cfg_en4292,
   output        cfg_en4293,
   output        cfg_en4294,
   output        cfg_en4295,
   output        cfg_en4296,
   output        cfg_en4297,
   output        cfg_en4298,
   output        cfg_en4299,
   output        cfg_en4300,
   output        cfg_en4301,
   output        cfg_en4302,
   output        cfg_en4303,
   output        cfg_en4304,
   output        cfg_en4305,
   output        cfg_en4306,
   output        cfg_en4307,
   output        cfg_en4308,
   output        cfg_en4309,
   output        cfg_en4310,
   output        cfg_en4311,
   output        cfg_en4312,
   output        cfg_en4313,
   output        cfg_en4314,
   output        cfg_en4315,
   output        cfg_en4316,
   output        cfg_en4317,
   output        cfg_en4318,
   output        cfg_en4319,
   output        cfg_en4320,
   output        cfg_en4321,
   output        cfg_en4322,
   output        cfg_en4323,
   output        cfg_en4324,
   output        cfg_en4325,
   output        cfg_en4326,
   output        cfg_en4327,
   output        cfg_en4328,
   output        cfg_en4329,
   output        cfg_en4330,
   output        cfg_en4331,
   output        cfg_en4332,
   output        cfg_en4333,
   output        cfg_en4334,
   output        cfg_en4335,
   output        cfg_en4336,
   output        cfg_en4337,
   output        cfg_en4338,
   output        cfg_en4339,
   output        cfg_en4340,
   output        cfg_en4341,
   output        cfg_en4342,
   output        cfg_en4343,
   output        cfg_en4344,
   output        cfg_en4345,
   output        cfg_en4346,
   output        cfg_en4347,
   output        cfg_en4348,
   output        cfg_en4349,
   output        cfg_en4350,
   output        cfg_en4351,
   output        cfg_en4352,
   output        cfg_en4353,
   output        cfg_en4354,
   output        cfg_en4355,
   output        cfg_en4356,
   output        cfg_en4357,
   output        cfg_en4358,
   output        cfg_en4359,
   output        cfg_en4360,
   output        cfg_en4361,
   output        cfg_en4362,
   output        cfg_en4363,
   output        cfg_en4364,
   output        cfg_en4365,
   output        cfg_en4366,
   output        cfg_en4367,
   output        cfg_en4368,
   output        cfg_en4369,
   output        cfg_en4370,
   output        cfg_en4371,
   output        cfg_en4372,
   output        cfg_en4373,
   output        cfg_en4374,
   output        cfg_en4375,
   output        cfg_en4376,
   output        cfg_en4377,
   output        cfg_en4378,
   output        cfg_en4379,
   output        cfg_en4380,
   output        cfg_en4381,
   output        cfg_en4382,
   output        cfg_en4383,
   output        cfg_en4384,
   output        cfg_en4385,
   output        cfg_en4386,
   output        cfg_en4387,
   output        cfg_en4388,
   output        cfg_en4389,
   output        cfg_en4390,
   output        cfg_en4391,
   output        cfg_en4392,
   output        cfg_en4393,
   output        cfg_en4394,
   output        cfg_en4395,
   output        cfg_en4396,
   output        cfg_en4397,
   output        cfg_en4398,
   output        cfg_en4399,
   output        cfg_en4400,
   output        cfg_en4401,
   output        cfg_en4402,
   output        cfg_en4403,
   output        cfg_en4404,
   output        cfg_en4405,
   output        cfg_en4406,
   output        cfg_en4407,
   output        cfg_en4408,
   output        cfg_en4409,
   output        cfg_en4410,
   output        cfg_en4411,
   output        cfg_en4412,
   output        cfg_en4413,
   output        cfg_en4414,
   output        cfg_en4415,
   output        cfg_en4416,
   output        cfg_en4417,
   output        cfg_en4418,
   output        cfg_en4419,
   output        cfg_en4420,
   output        cfg_en4421,
   output        cfg_en4422,
   output        cfg_en4423,
   output        cfg_en4424,
   output        cfg_en4425,
   output        cfg_en4426,
   output        cfg_en4427,
   output        cfg_en4428,
   output        cfg_en4429,
   output        cfg_en4430,
   output        cfg_en4431,
   output        cfg_en4432,
   output        cfg_en4433,
   output        cfg_en4434,
   output        cfg_en4435,
   output        cfg_en4436,
   output        cfg_en4437,
   output        cfg_en4438,
   output        cfg_en4439,
   output        cfg_en4440,
   output        cfg_en4441,
   output        cfg_en4442,
   output        cfg_en4443,
   output        cfg_en4444,
   output        cfg_en4445,
   output        cfg_en4446,
   output        cfg_en4447,
   output        cfg_en4448,
   output        cfg_en4449,
   output        cfg_en4450,
   output        cfg_en4451,
   output        cfg_en4452,
   output        cfg_en4453,
   output        cfg_en4454,
   output        cfg_en4455,
   output        cfg_en4456,
   output        cfg_en4457,
   output        cfg_en4458,
   output        cfg_en4459,
   output        cfg_en4460,
   output        cfg_en4461,
   output        cfg_en4462,
   output        cfg_en4463,
   output        cfg_en4464,
   output        cfg_en4465,
   output        cfg_en4466,
   output        cfg_en4467,
   output        cfg_en4468,
   output        cfg_en4469,
   output        cfg_en4470,
   output        cfg_en4471,
   output        cfg_en4472,
   output        cfg_en4473,
   output        cfg_en4474,
   output        cfg_en4475,
   output        cfg_en4476,
   output        cfg_en4477,
   output        cfg_en4478,
   output        cfg_en4479,
   output        cfg_en4480,
   output        cfg_en4481,
   output        cfg_en4482,
   output        cfg_en4483,
   output        cfg_en4484,
   output        cfg_en4485,
   output        cfg_en4486,
   output        cfg_en4487,
   output        cfg_en4488,
   output        cfg_en4489,
   output        cfg_en4490,
   output        cfg_en4491,
   output        cfg_en4492,
   output        cfg_en4493,
   output        cfg_en4494,
   output        cfg_en4495,
   output        cfg_en4496,
   output        cfg_en4497,
   output        cfg_en4498,
   output        cfg_en4499,
   output        cfg_en4500,
   output        cfg_en4501,
   output        cfg_en4502,
   output        cfg_en4503,
   output        cfg_en4504,
   output        cfg_en4505,
   output        cfg_en4506,
   output        cfg_en4507,
   output        cfg_en4508,
   output        cfg_en4509,
   output        cfg_en4510,
   output        cfg_en4511,
   output        cfg_en4512,
   output        cfg_en4513,
   output        cfg_en4514,
   output        cfg_en4515,
   output        cfg_en4516,
   output        cfg_en4517,
   output        cfg_en4518,
   output        cfg_en4519,
   output        cfg_en4520,
   output        cfg_en4521,
   output        cfg_en4522,
   output        cfg_en4523,
   output        cfg_en4524,
   output        cfg_en4525,
   output        cfg_en4526,
   output        cfg_en4527,
   output        cfg_en4528,
   output        cfg_en4529,
   output        cfg_en4530,
   output        cfg_en4531,
   output        cfg_en4532,
   output        cfg_en4533,
   output        cfg_en4534,
   output        cfg_en4535,
   output        cfg_en4536,
   output        cfg_en4537,
   output        cfg_en4538,
   output        cfg_en4539,
   output        cfg_en4540,
   output        cfg_en4541,
   output        cfg_en4542,
   output        cfg_en4543,
   output        cfg_en4544,
   output        cfg_en4545,
   output        cfg_en4546,
   output        cfg_en4547,
   output        cfg_en4548,
   output        cfg_en4549,
   output        cfg_en4550,
   output        cfg_en4551,
   output        cfg_en4552,
   output        cfg_en4553,
   output        cfg_en4554,
   output        cfg_en4555,
   output        cfg_en4556,
   output        cfg_en4557,
   output        cfg_en4558,
   output        cfg_en4559,
   output        cfg_en4560,
   output        cfg_en4561,
   output        cfg_en4562,
   output        cfg_en4563,
   output        cfg_en4564,
   output        cfg_en4565,
   output        cfg_en4566,
   output        cfg_en4567,
   output        cfg_en4568,
   output        cfg_en4569,
   output        cfg_en4570,
   output        cfg_en4571,
   output        cfg_en4572,
   output        cfg_en4573,
   output        cfg_en4574,
   output        cfg_en4575,
   output        cfg_en4576,
   output        cfg_en4577,
   output        cfg_en4578,
   output        cfg_en4579,
   output        cfg_en4580,
   output        cfg_en4581,
   output        cfg_en4582,
   output        cfg_en4583,
   output        cfg_en4584,
   output        cfg_en4585,
   output        cfg_en4586,
   output        cfg_en4587,
   output        cfg_en4588,
   output        cfg_en4589,
   output        cfg_en4590,
   output        cfg_en4591,
   output        cfg_en4592,
   output        cfg_en4593,
   output        cfg_en4594,
   output        cfg_en4595,
   output        cfg_en4596,
   output        cfg_en4597,
   output        cfg_en4598,
   output        cfg_en4599,
   output        cfg_en4600,
   output        cfg_en4601,
   output        cfg_en4602,
   output        cfg_en4603,
   output        cfg_en4604,
   output        cfg_en4605,
   output        cfg_en4606,
   output        cfg_en4607,
   output        cfg_en4608,
   output        cfg_en4609,
   output        cfg_en4610,
   output        cfg_en4611,
   output        cfg_en4612,
   output        cfg_en4613,
   output        cfg_en4614,
   output        cfg_en4615,
   output        cfg_en4616,
   output        cfg_en4617,
   output        cfg_en4618,
   output        cfg_en4619,
   output        cfg_en4620,
   output        cfg_en4621,
   output        cfg_en4622,
   output        cfg_en4623,
   output        cfg_en4624,
   output        cfg_en4625,
   output        cfg_en4626,
   output        cfg_en4627,
   output        cfg_en4628,
   output        cfg_en4629,
   output        cfg_en4630,
   output        cfg_en4631,
   output        cfg_en4632,
   output        cfg_en4633,
   output        cfg_en4634,
   output        cfg_en4635,
   output        cfg_en4636,
   output        cfg_en4637,
   output        cfg_en4638,
   output        cfg_en4639,
   output        cfg_en4640,
   output        cfg_en4641,
   output        cfg_en4642,
   output        cfg_en4643,
   output        cfg_en4644,
   output        cfg_en4645,
   output        cfg_en4646,
   output        cfg_en4647,
   output        cfg_en4648,
   output        cfg_en4649,
   output        cfg_en4650,
   output        cfg_en4651,
   output        cfg_en4652,
   output        cfg_en4653,
   output        cfg_en4654,
   output        cfg_en4655,
   output        cfg_en4656,
   output        cfg_en4657,
   output        cfg_en4658,
   output        cfg_en4659,
   output        cfg_en4660,
   output        cfg_en4661,
   output        cfg_en4662,
   output        cfg_en4663,
   output        cfg_en4664,
   output        cfg_en4665,
   output        cfg_en4666,
   output        cfg_en4667,
   output        cfg_en4668,
   output        cfg_en4669,
   output        cfg_en4670,
   output        cfg_en4671,
   output        cfg_en4672,
   output        cfg_en4673,
   output        cfg_en4674,
   output        cfg_en4675,
   output        cfg_en4676,
   output        cfg_en4677,
   output        cfg_en4678,
   output        cfg_en4679,
   output        cfg_en4680,
   output        cfg_en4681,
   output        cfg_en4682,
   output        cfg_en4683,
   output        cfg_en4684,
   output        cfg_en4685,
   output        cfg_en4686,
   output        cfg_en4687,
   output        cfg_en4688,
   output        cfg_en4689,
   output        cfg_en4690,
   output        cfg_en4691,
   output        cfg_en4692,
   output        cfg_en4693,
   output        cfg_en4694,
   output        cfg_en4695,
   output        cfg_en4696,
   output        cfg_en4697,
   output        cfg_en4698,
   output        cfg_en4699,
   output        cfg_en4700,
   output        cfg_en4701,
   output        cfg_en4702,
   output        cfg_en4703,
   output        cfg_en4704,
   output        cfg_en4705,
   output        cfg_en4706,
   output        cfg_en4707,
   output        cfg_en4708,
   output        cfg_en4709,
   output        cfg_en4710,
   output        cfg_en4711,
   output        cfg_en4712,
   output        cfg_en4713,
   output        cfg_en4714,
   output        cfg_en4715,
   output        cfg_en4716,
   output        cfg_en4717,
   output        cfg_en4718,
   output        cfg_en4719,
   output        cfg_en4720,
   output        cfg_en4721,
   output        cfg_en4722,
   output        cfg_en4723,
   output        cfg_en4724,
   output        cfg_en4725,
   output        cfg_en4726,
   output        cfg_en4727,
   output        cfg_en4728,
   output        cfg_en4729,
   output        cfg_en4730,
   output        cfg_en4731,
   output        cfg_en4732,
   output        cfg_en4733,
   output        cfg_en4734,
   output        cfg_en4735,
   output        cfg_en4736,
   output        cfg_en4737,
   output        cfg_en4738,
   output        cfg_en4739,
   output        cfg_en4740,
   output        cfg_en4741,
   output        cfg_en4742,
   output        cfg_en4743,
   output        cfg_en4744,
   output        cfg_en4745,
   output        cfg_en4746,
   output        cfg_en4747,
   output        cfg_en4748,
   output        cfg_en4749,
   output        cfg_en4750,
   output        cfg_en4751,
   output        cfg_en4752,
   output        cfg_en4753,
   output        cfg_en4754,
   output        cfg_en4755,
   output        cfg_en4756,
   output        cfg_en4757,
   output        cfg_en4758,
   output        cfg_en4759,
   output        cfg_en4760,
   output        cfg_en4761,
   output        cfg_en4762,
   output        cfg_en4763,
   output        cfg_en4764,
   output        cfg_en4765,
   output        cfg_en4766,
   output        cfg_en4767,
   output        cfg_en4768,
   output        cfg_en4769,
   output        cfg_en4770,
   output        cfg_en4771,
   output        cfg_en4772,
   output        cfg_en4773,
   output        cfg_en4774,
   output        cfg_en4775,
   output        cfg_en4776,
   output        cfg_en4777,
   output        cfg_en4778,
   output        cfg_en4779,
   output        cfg_en4780,
   output        cfg_en4781,
   output        cfg_en4782,
   output        cfg_en4783,
   output        cfg_en4784,
   output        cfg_en4785,
   output        cfg_en4786,
   output        cfg_en4787,
   output        cfg_en4788,
   output        cfg_en4789,
   output        cfg_en4790,
   output        cfg_en4791,
   output        cfg_en4792,
   output        cfg_en4793,
   output        cfg_en4794,
   output        cfg_en4795,
   output        cfg_en4796,
   output        cfg_en4797,
   output        cfg_en4798,
   output        cfg_en4799,
   output        cfg_en4800,
   output        cfg_en4801,
   output        cfg_en4802,
   output        cfg_en4803,
   output        cfg_en4804,
   output        cfg_en4805,
   output        cfg_en4806,
   output        cfg_en4807,
   output        cfg_en4808,
   output        cfg_en4809,
   output        cfg_en4810,
   output        cfg_en4811,
   output        cfg_en4812,
   output        cfg_en4813,
   output        cfg_en4814,
   output        cfg_en4815,
   output        cfg_en4816,
   output        cfg_en4817,
   output        cfg_en4818,
   output        cfg_en4819,
   output        cfg_en4820,
   output        cfg_en4821,
   output        cfg_en4822,
   output        cfg_en4823,
   output        cfg_en4824,
   output        cfg_en4825,
   output        cfg_en4826,
   output        cfg_en4827,
   output        cfg_en4828,
   output        cfg_en4829,
   output        cfg_en4830,
   output        cfg_en4831,
   output        cfg_en4832,
   output        cfg_en4833,
   output        cfg_en4834,
   output        cfg_en4835,
   output        cfg_en4836,
   output        cfg_en4837,
   output        cfg_en4838,
   output        cfg_en4839,
   output        cfg_en4840,
   output        cfg_en4841,
   output        cfg_en4842,
   output        cfg_en4843,
   output        cfg_en4844,
   output        cfg_en4845,
   output        cfg_en4846,
   output        cfg_en4847,
   output        cfg_en4848,
   output        cfg_en4849,
   output        cfg_en4850,
   output        cfg_en4851,
   output        cfg_en4852,
   output        cfg_en4853,
   output        cfg_en4854,
   output        cfg_en4855,
   output        cfg_en4856,
   output        cfg_en4857,
   output        cfg_en4858,
   output        cfg_en4859,
   output        cfg_en4860,
   output        cfg_en4861,
   output        cfg_en4862,
   output        cfg_en4863,
   output        cfg_en4864,
   output        cfg_en4865,
   output        cfg_en4866,
   output        cfg_en4867,
   output        cfg_en4868,
   output        cfg_en4869,
   output        cfg_en4870,
   output        cfg_en4871,
   output        cfg_en4872,
   output        cfg_en4873,
   output        cfg_en4874,
   output        cfg_en4875,
   output        cfg_en4876,
   output        cfg_en4877,
   output        cfg_en4878,
   output        cfg_en4879,
   output        cfg_en4880,
   output        cfg_en4881,
   output        cfg_en4882,
   output        cfg_en4883,
   output        cfg_en4884,
   output        cfg_en4885,
   output        cfg_en4886,
   output        cfg_en4887,
   output        cfg_en4888,
   output        cfg_en4889,
   output        cfg_en4890,
   output        cfg_en4891,
   output        cfg_en4892,
   output        cfg_en4893,
   output        cfg_en4894,
   output        cfg_en4895,
   output        cfg_en4896,
   output        cfg_en4897,
   output        cfg_en4898,
   output        cfg_en4899,
   output        cfg_en4900,
   output        cfg_en4901,
   output        cfg_en4902,
   output        cfg_en4903,
   output        cfg_en4904,
   output        cfg_en4905,
   output        cfg_en4906,
   output        cfg_en4907,
   output        cfg_en4908,
   output        cfg_en4909,
   output        cfg_en4910,
   output        cfg_en4911,
   output        cfg_en4912,
   output        cfg_en4913,
   output        cfg_en4914,
   output        cfg_en4915,
   output        cfg_en4916,
   output        cfg_en4917,
   output        cfg_en4918,
   output        cfg_en4919,
   output        cfg_en4920,
   output        cfg_en4921,
   output        cfg_en4922,
   output        cfg_en4923,
   output        cfg_en4924,
   output        cfg_en4925,
   output        cfg_en4926,
   output        cfg_en4927,
   output        cfg_en4928,
   output        cfg_en4929,
   output        cfg_en4930,
   output        cfg_en4931,
   output        cfg_en4932,
   output        cfg_en4933,
   output        cfg_en4934,
   output        cfg_en4935,
   output        cfg_en4936,
   output        cfg_en4937,
   output        cfg_en4938,
   output        cfg_en4939,
   output        cfg_en4940,
   output        cfg_en4941,
   output        cfg_en4942,
   output        cfg_en4943,
   output        cfg_en4944,
   output        cfg_en4945,
   output        cfg_en4946,
   output        cfg_en4947,
   output        cfg_en4948,
   output        cfg_en4949,
   output        cfg_en4950,
   output        cfg_en4951,
   output        cfg_en4952,
   output        cfg_en4953,
   output        cfg_en4954,
   output        cfg_en4955,
   output        cfg_en4956,
   output        cfg_en4957,
   output        cfg_en4958,
   output        cfg_en4959,
   output        cfg_en4960,
   output        cfg_en4961,
   output        cfg_en4962,
   output        cfg_en4963,
   output        cfg_en4964,
   output        cfg_en4965,
   output        cfg_en4966,
   output        cfg_en4967,
   output        cfg_en4968,
   output        cfg_en4969,
   output        cfg_en4970,
   output        cfg_en4971,
   output        cfg_en4972,
   output        cfg_en4973,
   output        cfg_en4974,
   output        cfg_en4975,
   output        cfg_en4976,
   output        cfg_en4977,
   output        cfg_en4978,
   output        cfg_en4979,
   output        cfg_en4980,
   output        cfg_en4981,
   output        cfg_en4982,
   output        cfg_en4983,
   output        cfg_en4984,
   output        cfg_en4985,
   output        cfg_en4986,
   output        cfg_en4987,
   output        cfg_en4988,
   output        cfg_en4989,
   output        cfg_en4990,
   output        cfg_en4991,
   output        cfg_en4992,
   output        cfg_en4993,
   output        cfg_en4994,
   output        cfg_en4995,
   output        cfg_en4996,
   output        cfg_en4997,
   output        cfg_en4998,
   output        cfg_en4999,
   output        cfg_en5000,
   output        cfg_en5001,
   output        cfg_en5002,
   output        cfg_en5003,
   output        cfg_en5004,
   output        cfg_en5005,
   output        cfg_en5006,
   output        cfg_en5007,
   output        cfg_en5008,
   output        cfg_en5009,
   output        cfg_en5010,
   output        cfg_en5011,
   output        cfg_en5012,
   output        cfg_en5013,
   output        cfg_en5014,
   output        cfg_en5015,
   output        cfg_en5016,
   output        cfg_en5017,
   output        cfg_en5018,
   output        cfg_en5019,
   output        cfg_en5020,
   output        cfg_en5021,
   output        cfg_en5022,
   output        cfg_en5023,
   output        cfg_en5024,
   output        cfg_en5025,
   output        cfg_en5026,
   output        cfg_en5027,
   output        cfg_en5028,
   output        cfg_en5029,
   output        cfg_en5030,
   output        cfg_en5031,
   output        cfg_en5032,
   output        cfg_en5033,
   output        cfg_en5034,
   output        cfg_en5035,
   output        cfg_en5036,
   output        cfg_en5037,
   output        cfg_en5038,
   output        cfg_en5039,
   output        cfg_en5040,
   output        cfg_en5041,
   output        cfg_en5042,
   output        cfg_en5043,
   output        cfg_en5044,
   output        cfg_en5045,
   output        cfg_en5046,
   output        cfg_en5047,
   output        cfg_en5048,
   output        cfg_en5049,
   output        cfg_en5050,
   output        cfg_en5051,
   output        cfg_en5052,
   output        cfg_en5053,
   output        cfg_en5054,
   output        cfg_en5055,
   output        cfg_en5056,
   output        cfg_en5057,
   output        cfg_en5058,
   output        cfg_en5059,
   output        cfg_en5060,
   output        cfg_en5061,
   output        cfg_en5062,
   output        cfg_en5063,
   output        cfg_en5064,
   output        cfg_en5065,
   output        cfg_en5066,
   output        cfg_en5067,
   output        cfg_en5068,
   output        cfg_en5069,
   output        cfg_en5070,
   output        cfg_en5071,
   output        cfg_en5072,
   output        cfg_en5073,
   output        cfg_en5074,
   output        cfg_en5075,
   output        cfg_en5076,
   output        cfg_en5077,
   output        cfg_en5078,
   output        cfg_en5079,
   output        cfg_en5080,
   output        cfg_en5081,
   output        cfg_en5082,
   output        cfg_en5083,
   output        cfg_en5084,
   output        cfg_en5085,
   output        cfg_en5086,
   output        cfg_en5087,
   output        cfg_en5088,
   output        cfg_en5089,
   output        cfg_en5090,
   output        cfg_en5091,
   output        cfg_en5092,
   output        cfg_en5093,
   output        cfg_en5094,
   output        cfg_en5095,
   output        cfg_en5096,
   output        cfg_en5097,
   output        cfg_en5098,
   output        cfg_en5099,
   output        cfg_en5100,
   output        cfg_en5101,
   output        cfg_en5102,
   output        cfg_en5103,
   output        cfg_en5104,
   output        cfg_en5105,
   output        cfg_en5106,
   output        cfg_en5107,
   output        cfg_en5108,
   output        cfg_en5109,
   output        cfg_en5110,
   output        cfg_en5111,
   output        cfg_en5112,
   output        cfg_en5113,
   output        cfg_en5114,
   output        cfg_en5115,
   output        cfg_en5116,
   output        cfg_en5117,
   output        cfg_en5118,
   output        cfg_en5119,
   output        cfg_en5120,
   output        cfg_en5121,
   output        cfg_en5122,
   output        cfg_en5123,
   output        cfg_en5124,
   output        cfg_en5125,
   output        cfg_en5126,
   output        cfg_en5127,
   output        cfg_en5128,
   output        cfg_en5129,
   output        cfg_en5130,
   output        cfg_en5131,
   output        cfg_en5132,
   output        cfg_en5133,
   output        cfg_en5134,
   output        cfg_en5135,
   output        cfg_en5136,
   output        cfg_en5137,
   output        cfg_en5138,
   output        cfg_en5139,
   output        cfg_en5140,
   output        cfg_en5141,
   output        cfg_en5142,
   output        cfg_en5143,
   output        cfg_en5144,
   output        cfg_en5145,
   output        cfg_en5146,
   output        cfg_en5147,
   output        cfg_en5148,
   output        cfg_en5149,
   output        cfg_en5150,
   output        cfg_en5151,
   output        cfg_en5152,
   output        cfg_en5153,
   output        cfg_en5154,
   output        cfg_en5155,
   output        cfg_en5156,
   output        cfg_en5157,
   output        cfg_en5158,
   output        cfg_en5159,
   output        cfg_en5160,
   output        cfg_en5161,
   output        cfg_en5162,
   output        cfg_en5163,
   output        cfg_en5164,
   output        cfg_en5165,
   output        cfg_en5166,
   output        cfg_en5167,
   output        cfg_en5168,
   output        cfg_en5169,
   output        cfg_en5170,
   output        cfg_en5171,
   output        cfg_en5172,
   output        cfg_en5173,
   output        cfg_en5174,
   output        cfg_en5175,
   output        cfg_en5176,
   output        cfg_en5177,
   output        cfg_en5178,
   output        cfg_en5179,
   output        cfg_en5180,
   output        cfg_en5181,
   output        cfg_en5182,
   output        cfg_en5183,
   output        cfg_en5184,
   output        cfg_en5185,
   output        cfg_en5186,
   output        cfg_en5187,
   output        cfg_en5188,
   output        cfg_en5189,
   output        cfg_en5190,
   output        cfg_en5191,
   output        cfg_en5192,
   output        cfg_en5193,
   output        cfg_en5194,
   output        cfg_en5195,
   output        cfg_en5196,
   output        cfg_en5197,
   output        cfg_en5198,
   output        cfg_en5199,
   output        cfg_en5200,
   output        cfg_en5201,
   output        cfg_en5202,
   output        cfg_en5203,
   output        cfg_en5204,
   output        cfg_en5205,
   output        cfg_en5206,
   output        cfg_en5207,
   output        cfg_en5208,
   output        cfg_en5209,
   output        cfg_en5210,
   output        cfg_en5211,
   output        cfg_en5212,
   output        cfg_en5213,
   output        cfg_en5214,
   output        cfg_en5215,
   output        cfg_en5216,
   output        cfg_en5217,
   output        cfg_en5218,
   output        cfg_en5219,
   output        cfg_en5220,
   output        cfg_en5221,
   output        cfg_en5222,
   output        cfg_en5223,
   output        cfg_en5224,
   output        cfg_en5225,
   output        cfg_en5226,
   output        cfg_en5227,
   output        cfg_en5228,
   output        cfg_en5229,
   output        cfg_en5230,
   output        cfg_en5231,
   output        cfg_en5232,
   output        cfg_en5233,
   output        cfg_en5234,
   output        cfg_en5235,
   output        cfg_en5236,
   output        cfg_en5237,
   output        cfg_en5238,
   output        cfg_en5239,
   output        cfg_en5240,
   output        cfg_en5241,
   output        cfg_en5242,
   output        cfg_en5243,
   output        cfg_en5244,
   output        cfg_en5245,
   output        cfg_en5246,
   output        cfg_en5247,
   output        cfg_en5248,
   output        cfg_en5249,
   output        cfg_en5250,
   output        cfg_en5251,
   output        cfg_en5252,
   output        cfg_en5253,
   output        cfg_en5254,
   output        cfg_en5255,
   output        cfg_en5256,
   output        cfg_en5257,
   output        cfg_en5258,
   output        cfg_en5259,
   output        cfg_en5260,
   output        cfg_en5261,
   output        cfg_en5262,
   output        cfg_en5263,
   output        cfg_en5264,
   output        cfg_en5265,
   output        cfg_en5266,
   output        cfg_en5267,
   output        cfg_en5268,
   output        cfg_en5269,
   output        cfg_en5270,
   output        cfg_en5271,
   output        cfg_en5272,
   output        cfg_en5273,
   output        cfg_en5274,
   output        cfg_en5275,
   output        cfg_en5276,
   output        cfg_en5277,
   output        cfg_en5278,
   output        cfg_en5279,
   output        cfg_en5280,
   output        cfg_en5281,
   output        cfg_en5282,
   output        cfg_en5283,
   output        cfg_en5284,
   output        cfg_en5285,
   output        cfg_en5286,
   output        cfg_en5287,
   output        cfg_en5288,
   output        cfg_en5289,
   output        cfg_en5290,
   output        cfg_en5291,
   output        cfg_en5292,
   output        cfg_en5293,
   output        cfg_en5294,
   output        cfg_en5295,
   output        cfg_en5296,
   output        cfg_en5297,
   output        cfg_en5298,
   output        cfg_en5299,
   output        cfg_en5300,
   output        cfg_en5301,
   output        cfg_en5302,
   output        cfg_en5303,
   output        cfg_en5304,
   output        cfg_en5305,
   output        cfg_en5306,
   output        cfg_en5307,
   output        cfg_en5308,
   output        cfg_en5309,
   output        cfg_en5310,
   output        cfg_en5311,
   output        cfg_en5312,
   output        cfg_en5313,
   output        cfg_en5314,
   output        cfg_en5315,
   output        cfg_en5316,
   output        cfg_en5317,
   output        cfg_en5318,
   output        cfg_en5319,
   output        cfg_en5320,
   output        cfg_en5321,
   output        cfg_en5322,
   output        cfg_en5323,
   output        cfg_en5324,
   output        cfg_en5325,
   output        cfg_en5326,
   output        cfg_en5327,
   output        cfg_en5328,
   output        cfg_en5329,
   output        cfg_en5330,
   output        cfg_en5331,
   output        cfg_en5332,
   output        cfg_en5333,
   output        cfg_en5334,
   output        cfg_en5335,
   output        cfg_en5336,
   output        cfg_en5337,
   output        cfg_en5338,
   output        cfg_en5339,
   output        cfg_en5340,
   output        cfg_en5341,
   output        cfg_en5342,
   output        cfg_en5343,
   output        cfg_en5344,
   output        cfg_en5345,
   output        cfg_en5346,
   output        cfg_en5347,
   output        cfg_en5348,
   output        cfg_en5349,
   output        cfg_en5350,
   output        cfg_en5351,
   output        cfg_en5352,
   output        cfg_en5353,
   output        cfg_en5354,
   output        cfg_en5355,
   output        cfg_en5356,
   output        cfg_en5357,
   output        cfg_en5358,
   output        cfg_en5359,
   output        cfg_en5360,
   output        cfg_en5361,
   output        cfg_en5362,
   output        cfg_en5363,
   output        cfg_en5364,
   output        cfg_en5365,
   output        cfg_en5366,
   output        cfg_en5367,
   output        cfg_en5368,
   output        cfg_en5369,
   output        cfg_en5370,
   output        cfg_en5371,
   output        cfg_en5372,
   output        cfg_en5373,
   output        cfg_en5374,
   output        cfg_en5375,
   output        cfg_en5376,
   output        cfg_en5377,
   output        cfg_en5378,
   output        cfg_en5379,
   output        cfg_en5380,
   output        cfg_en5381,
   output        cfg_en5382,
   output        cfg_en5383,
   output        cfg_en5384,
   output        cfg_en5385,
   output        cfg_en5386,
   output        cfg_en5387,
   output        cfg_en5388,
   output        cfg_en5389,
   output        cfg_en5390,
   output        cfg_en5391,
   output        cfg_en5392,
   output        cfg_en5393,
   output        cfg_en5394,
   output        cfg_en5395,
   output        cfg_en5396,
   output        cfg_en5397,
   output        cfg_en5398,
   output        cfg_en5399,
   output        cfg_en5400,
   output        cfg_en5401,
   output        cfg_en5402,
   output        cfg_en5403,
   output        cfg_en5404,
   output        cfg_en5405,
   output        cfg_en5406,
   output        cfg_en5407,
   output        cfg_en5408,
   output        cfg_en5409,
   output        cfg_en5410,
   output        cfg_en5411,
   output        cfg_en5412,
   output        cfg_en5413,
   output        cfg_en5414,
   output        cfg_en5415,
   output        cfg_en5416,
   output        cfg_en5417,
   output        cfg_en5418,
   output        cfg_en5419,
   output        cfg_en5420,
   output        cfg_en5421,
   output        cfg_en5422,
   output        cfg_en5423,
   output        cfg_en5424,
   output        cfg_en5425,
   output        cfg_en5426,
   output        cfg_en5427,
   output        cfg_en5428,
   output        cfg_en5429,
   output        cfg_en5430,
   output        cfg_en5431,
   output        cfg_en5432,
   output        cfg_en5433,
   output        cfg_en5434,
   output        cfg_en5435,
   output        cfg_en5436,
   output        cfg_en5437,
   output        cfg_en5438,
   output        cfg_en5439,
   output        cfg_en5440,
   output        cfg_en5441,
   output        cfg_en5442,
   output        cfg_en5443,
   output        cfg_en5444,
   output        cfg_en5445,
   output        cfg_en5446,
   output        cfg_en5447,
   output        cfg_en5448,
   output        cfg_en5449,
   output        cfg_en5450,
   output        cfg_en5451,
   output        cfg_en5452,
   output        cfg_en5453,
   output        cfg_en5454,
   output        cfg_en5455,
   output        cfg_en5456,
   output        cfg_en5457,
   output        cfg_en5458,
   output        cfg_en5459,
   output        cfg_en5460,
   output        cfg_en5461,
   output        cfg_en5462,
   output        cfg_en5463,
   output        cfg_en5464,
   output        cfg_en5465,
   output        cfg_en5466,
   output        cfg_en5467,
   output        cfg_en5468,
   output        cfg_en5469,
   output        cfg_en5470,
   output        cfg_en5471,
   output        cfg_en5472,
   output        cfg_en5473,
   output        cfg_en5474,
   output        cfg_en5475,
   output        cfg_en5476,
   output        cfg_en5477,
   output        cfg_en5478,
   output        cfg_en5479,
   output        cfg_en5480,
   output        cfg_en5481,
   output        cfg_en5482,
   output        cfg_en5483,
   output        cfg_en5484,
   output        cfg_en5485,
   output        cfg_en5486,
   output        cfg_en5487,
   output        cfg_en5488,
   output        cfg_en5489,
   output        cfg_en5490,
   output        cfg_en5491,
   output        cfg_en5492,
   output        cfg_en5493,
   output        cfg_en5494,
   output        cfg_en5495,
   output        cfg_en5496,
   output        cfg_en5497,
   output        cfg_en5498,
   output        cfg_en5499,
   output        cfg_en5500,
   output        cfg_en5501,
   output        cfg_en5502,
   output        cfg_en5503,
   output        cfg_en5504,
   output        cfg_en5505,
   output        cfg_en5506,
   output        cfg_en5507,
   output        cfg_en5508,
   output        cfg_en5509,
   output        cfg_en5510,
   output        cfg_en5511,
   output        cfg_en5512,
   output        cfg_en5513,
   output        cfg_en5514,
   output        cfg_en5515,
   output        cfg_en5516,
   output        cfg_en5517,
   output        cfg_en5518,
   output        cfg_en5519,
   output        cfg_en5520,
   output        cfg_en5521,
   output        cfg_en5522,
   output        cfg_en5523,
   output        cfg_en5524,
   output        cfg_en5525,
   output        cfg_en5526,
   output        cfg_en5527,
   output        cfg_en5528,
   output        cfg_en5529,
   output        cfg_en5530,
   output        cfg_en5531,
   output        cfg_en5532,
   output        cfg_en5533,
   output        cfg_en5534,
   output        cfg_en5535,
   output        cfg_en5536,
   output        cfg_en5537,
   output        cfg_en5538,
   output        cfg_en5539,
   output        cfg_en5540,
   output        cfg_en5541,
   output        cfg_en5542,
   output        cfg_en5543,
   output        cfg_en5544,
   output        cfg_en5545,
   output        cfg_en5546,
   output        cfg_en5547,
   output        cfg_en5548,
   output        cfg_en5549,
   output        cfg_en5550,
   output        cfg_en5551,
   output        cfg_en5552,
   output        cfg_en5553,
   output        cfg_en5554,
   output        cfg_en5555,
   output        cfg_en5556,
   output        cfg_en5557,
   output        cfg_en5558,
   output        cfg_en5559,
   output        cfg_en5560,
   output        cfg_en5561,
   output        cfg_en5562,
   output        cfg_en5563,
   output        cfg_en5564,
   output        cfg_en5565,
   output        cfg_en5566,
   output        cfg_en5567,
   output        cfg_en5568,
   output        cfg_en5569,
   output        cfg_en5570,
   output        cfg_en5571,
   output        cfg_en5572,
   output        cfg_en5573,
   output        cfg_en5574,
   output        cfg_en5575,
   output        cfg_en5576,
   output        cfg_en5577,
   output        cfg_en5578,
   output        cfg_en5579,
   output        cfg_en5580,
   output        cfg_en5581,
   output        cfg_en5582,
   output        cfg_en5583,
   output        cfg_en5584,
   output        cfg_en5585,
   output        cfg_en5586,
   output        cfg_en5587,
   output        cfg_en5588,
   output        cfg_en5589,
   output        cfg_en5590,
   output        cfg_en5591,
   output        cfg_en5592,
   output        cfg_en5593,
   output        cfg_en5594,
   output        cfg_en5595,
   output        cfg_en5596,
   output        cfg_en5597,
   output        cfg_en5598,
   output        cfg_en5599,
   output        cfg_en5600,
   output        cfg_en5601,
   output        cfg_en5602,
   output        cfg_en5603,
   output        cfg_en5604,
   output        cfg_en5605,
   output        cfg_en5606,
   output        cfg_en5607,
   output        cfg_en5608,
   output        cfg_en5609,
   output        cfg_en5610,
   output        cfg_en5611,
   output        cfg_en5612,
   output        cfg_en5613,
   output        cfg_en5614,
   output        cfg_en5615,
   output        cfg_en5616,
   output        cfg_en5617,
   output        cfg_en5618,
   output        cfg_en5619,
   output        cfg_en5620,
   output        cfg_en5621,
   output        cfg_en5622,
   output        cfg_en5623,
   output        cfg_en5624,
   output        cfg_en5625,
   output        cfg_en5626,
   output        cfg_en5627,
   output        cfg_en5628,
   output        cfg_en5629,
   output        cfg_en5630,
   output        cfg_en5631,
   output        cfg_en5632,
   output        cfg_en5633,
   output        cfg_en5634,
   output        cfg_en5635,
   output        cfg_en5636,
   output        cfg_en5637,
   output        cfg_en5638,
   output        cfg_en5639,
   output        cfg_en5640,
   output        cfg_en5641,
   output        cfg_en5642,
   output        cfg_en5643,
   output        cfg_en5644,
   output        cfg_en5645,
   output        cfg_en5646,
   output        cfg_en5647,
   output        cfg_en5648,
   output        cfg_en5649,
   output        cfg_en5650,
   output        cfg_en5651,
   output        cfg_en5652,
   output        cfg_en5653,
   output        cfg_en5654,
   output        cfg_en5655,
   output        cfg_en5656,
   output        cfg_en5657,
   output        cfg_en5658,
   output        cfg_en5659,
   output        cfg_en5660,
   output        cfg_en5661,
   output        cfg_en5662,
   output        cfg_en5663,
   output        cfg_en5664,
   output        cfg_en5665,
   output        cfg_en5666,
   output        cfg_en5667,
   output        cfg_en5668,
   output        cfg_en5669,
   output        cfg_en5670,
   output        cfg_en5671,
   output        cfg_en5672,
   output        cfg_en5673,
   output        cfg_en5674,
   output        cfg_en5675,
   output        cfg_en5676,
   output        cfg_en5677,
   output        cfg_en5678,
   output        cfg_en5679,
   output        cfg_en5680,
   output        cfg_en5681,
   output        cfg_en5682,
   output        cfg_en5683,
   output        cfg_en5684,
   output        cfg_en5685,
   output        cfg_en5686,
   output        cfg_en5687,
   output        cfg_en5688,
   output        cfg_en5689,
   output        cfg_en5690,
   output        cfg_en5691,
   output        cfg_en5692,
   output        cfg_en5693,
   output        cfg_en5694,
   output        cfg_en5695,
   output        cfg_en5696,
   output        cfg_en5697,
   output        cfg_en5698,
   output        cfg_en5699,
   output        cfg_en5700,
   output        cfg_en5701,
   output        cfg_en5702,
   output        cfg_en5703,
   output        cfg_en5704,
   output        cfg_en5705,
   output        cfg_en5706,
   output        cfg_en5707,
   output        cfg_en5708,
   output        cfg_en5709,
   output        cfg_en5710,
   output        cfg_en5711,
   output        cfg_en5712,
   output        cfg_en5713,
   output        cfg_en5714,
   output        cfg_en5715,
   output        cfg_en5716,
   output        cfg_en5717,
   output        cfg_en5718,
   output        cfg_en5719,
   output        cfg_en5720,
   output        cfg_en5721,
   output        cfg_en5722,
   output        cfg_en5723,
   output        cfg_en5724,
   output        cfg_en5725,
   output        cfg_en5726,
   output        cfg_en5727,
   output        cfg_en5728,
   output        cfg_en5729,
   output        cfg_en5730,
   output        cfg_en5731,
   output        cfg_en5732,
   output        cfg_en5733,
   output        cfg_en5734,
   output        cfg_en5735,
   output        cfg_en5736,
   output        cfg_en5737,
   output        cfg_en5738,
   output        cfg_en5739,
   output        cfg_en5740,
   output        cfg_en5741,
   output        cfg_en5742,
   output        cfg_en5743,
   output        cfg_en5744,
   output        cfg_en5745,
   output        cfg_en5746,
   output        cfg_en5747,
   output        cfg_en5748,
   output        cfg_en5749,
   output        cfg_en5750,
   output        cfg_en5751,
   output        cfg_en5752,
   output        cfg_en5753,
   output        cfg_en5754,
   output        cfg_en5755,
   output        cfg_en5756,
   output        cfg_en5757,
   output        cfg_en5758,
   output        cfg_en5759,
   output        cfg_en5760,
   output        cfg_en5761,
   output        cfg_en5762,
   output        cfg_en5763,
   output        cfg_en5764,
   output        cfg_en5765,
   output        cfg_en5766,
   output        cfg_en5767,
   output        cfg_en5768,
   output        cfg_en5769,
   output        cfg_en5770,
   output        cfg_en5771,
   output        cfg_en5772,
   output        cfg_en5773,
   output        cfg_en5774,
   output        cfg_en5775,
   output        cfg_en5776,
   output        cfg_en5777,
   output        cfg_en5778,
   output        cfg_en5779,
   output        cfg_en5780,
   output        cfg_en5781,
   output        cfg_en5782,
   output        cfg_en5783,
   output        cfg_en5784,
   output        cfg_en5785,
   output        cfg_en5786,
   output        cfg_en5787,
   output        cfg_en5788,
   output        cfg_en5789,
   output        cfg_en5790,
   output        cfg_en5791,
   output        cfg_en5792,
   output        cfg_en5793,
   output        cfg_en5794,
   output        cfg_en5795,
   output        cfg_en5796,
   output        cfg_en5797,
   output        cfg_en5798,
   output        cfg_en5799,
   output        cfg_en5800,
   output        cfg_en5801,
   output        cfg_en5802,
   output        cfg_en5803,
   output        cfg_en5804,
   output        cfg_en5805,
   output        cfg_en5806,
   output        cfg_en5807,
   output        cfg_en5808,
   output        cfg_en5809,
   output        cfg_en5810,
   output        cfg_en5811,
   output        cfg_en5812,
   output        cfg_en5813,
   output        cfg_en5814,
   output        cfg_en5815,
   output        cfg_en5816,
   output        cfg_en5817,
   output        cfg_en5818,
   output        cfg_en5819,
   output        cfg_en5820,
   output        cfg_en5821,
   output        cfg_en5822,
   output        cfg_en5823,
   output        cfg_en5824,
   output        cfg_en5825,
   output        cfg_en5826,
   output        cfg_en5827,
   output        cfg_en5828,
   output        cfg_en5829,
   output        cfg_en5830,
   output        cfg_en5831,
   output        cfg_en5832,
   output        cfg_en5833,
   output        cfg_en5834,
   output        cfg_en5835,
   output        cfg_en5836,
   output        cfg_en5837,
   output        cfg_en5838,
   output        cfg_en5839,
   output        cfg_en5840,
   output        cfg_en5841,
   output        cfg_en5842,
   output        cfg_en5843,
   output        cfg_en5844,
   output        cfg_en5845,
   output        cfg_en5846,
   output        cfg_en5847,
   output        cfg_en5848,
   output        cfg_en5849,
   output        cfg_en5850,
   output        cfg_en5851,
   output        cfg_en5852,
   output        cfg_en5853,
   output        cfg_en5854,
   output        cfg_en5855,
   output        cfg_en5856,
   output        cfg_en5857,
   output        cfg_en5858,
   output        cfg_en5859,
   output        cfg_en5860,
   output        cfg_en5861,
   output        cfg_en5862,
   output        cfg_en5863,
   output        cfg_en5864,
   output        cfg_en5865,
   output        cfg_en5866,
   output        cfg_en5867,
   output        cfg_en5868,
   output        cfg_en5869,
   output        cfg_en5870,
   output        cfg_en5871,
   output        cfg_en5872,
   output        cfg_en5873,
   output        cfg_en5874,
   output        cfg_en5875,
   output        cfg_en5876,
   output        cfg_en5877,
   output        cfg_en5878,
   output        cfg_en5879,
   output        cfg_en5880,
   output        cfg_en5881,
   output        cfg_en5882,
   output        cfg_en5883,
   output        cfg_en5884,
   output        cfg_en5885,
   output        cfg_en5886,
   output        cfg_en5887,
   output        cfg_en5888,
   output        cfg_en5889,
   output        cfg_en5890,
   output        cfg_en5891,
   output        cfg_en5892,
   output        cfg_en5893,
   output        cfg_en5894,
   output        cfg_en5895,
   output        cfg_en5896,
   output        cfg_en5897,
   output        cfg_en5898,
   output        cfg_en5899,
   output        cfg_en5900,
   output        cfg_en5901,
   output        cfg_en5902,
   output        cfg_en5903,
   output        cfg_en5904,
   output        cfg_en5905,
   output        cfg_en5906,
   output        cfg_en5907,
   output        cfg_en5908,
   output        cfg_en5909,
   output        cfg_en5910,
   output        cfg_en5911,
   output        cfg_en5912,
   output        cfg_en5913,
   output        cfg_en5914,
   output        cfg_en5915,
   output        cfg_en5916,
   output        cfg_en5917,
   output        cfg_en5918,
   output        cfg_en5919,
   output        cfg_en5920,
   output        cfg_en5921,
   output        cfg_en5922,
   output        cfg_en5923,
   output        cfg_en5924,
   output        cfg_en5925,
   output        cfg_en5926,
   output        cfg_en5927,
   output        cfg_en5928,
   output        cfg_en5929,
   output        cfg_en5930,
   output        cfg_en5931,
   output        cfg_en5932,
   output        cfg_en5933,
   output        cfg_en5934,
   output        cfg_en5935,
   output        cfg_en5936,
   output        cfg_en5937,
   output        cfg_en5938,
   output        cfg_en5939,
   output        cfg_en5940,
   output        cfg_en5941,
   output        cfg_en5942,
   output        cfg_en5943,
   output        cfg_en5944,
   output        cfg_en5945,
   output        cfg_en5946,
   output        cfg_en5947,
   output        cfg_en5948,
   output        cfg_en5949,
   output        cfg_en5950,
   output        cfg_en5951,
   output        cfg_en5952,
   output        cfg_en5953,
   output        cfg_en5954,
   output        cfg_en5955,
   output        cfg_en5956,
   output        cfg_en5957,
   output        cfg_en5958,
   output        cfg_en5959,
   output        cfg_en5960,
   output        cfg_en5961,
   output        cfg_en5962,
   output        cfg_en5963,
   output        cfg_en5964,
   output        cfg_en5965,
   output        cfg_en5966,
   output        cfg_en5967,
   output        cfg_en5968,
   output        cfg_en5969,
   output        cfg_en5970,
   output        cfg_en5971,
   output        cfg_en5972,
   output        cfg_en5973,
   output        cfg_en5974,
   output        cfg_en5975,
   output        cfg_en5976,
   output        cfg_en5977,
   output        cfg_en5978,
   output        cfg_en5979,
   output        cfg_en5980,
   output        cfg_en5981,
   output        cfg_en5982,
   output        cfg_en5983,
   output        cfg_en5984,
   output        cfg_en5985,
   output        cfg_en5986,
   output        cfg_en5987,
   output        cfg_en5988,
   output        cfg_en5989,
   output        cfg_en5990,
   output        cfg_en5991,
   output        cfg_en5992,
   output        cfg_en5993,
   output        cfg_en5994,
   output        cfg_en5995,
   output        cfg_en5996,
   output        cfg_en5997,
   output        cfg_en5998,
   output        cfg_en5999,
   output        cfg_en6000,
   output        cfg_en6001,
   output        cfg_en6002,
   output        cfg_en6003,
   output        cfg_en6004,
   output        cfg_en6005,
   output        cfg_en6006,
   output        cfg_en6007,
   output        cfg_en6008,
   output        cfg_en6009,
   output        cfg_en6010,
   output        cfg_en6011,
   output        cfg_en6012,
   output        cfg_en6013,
   output        cfg_en6014,
   output        cfg_en6015,
   output        cfg_en6016,
   output        cfg_en6017,
   output        cfg_en6018,
   output        cfg_en6019,
   output        cfg_en6020,
   output        cfg_en6021,
   output        cfg_en6022,
   output        cfg_en6023,
   output        cfg_en6024,
   output        cfg_en6025,
   output        cfg_en6026,
   output        cfg_en6027,
   output        cfg_en6028,
   output        cfg_en6029,
   output        cfg_en6030,
   output        cfg_en6031,
   output        cfg_en6032,
   output        cfg_en6033,
   output        cfg_en6034,
   output        cfg_en6035,
   output        cfg_en6036,
   output        cfg_en6037,
   output        cfg_en6038,
   output        cfg_en6039,
   output        cfg_en6040,
   output        cfg_en6041,
   output        cfg_en6042,
   output        cfg_en6043,
   output        cfg_en6044,
   output        cfg_en6045,
   output        cfg_en6046,
   output        cfg_en6047,
   output        cfg_en6048,
   output        cfg_en6049,
   output        cfg_en6050,
   output        cfg_en6051,
   output        cfg_en6052,
   output        cfg_en6053,
   output        cfg_en6054,
   output        cfg_en6055,
   output        cfg_en6056,
   output        cfg_en6057,
   output        cfg_en6058,
   output        cfg_en6059,
   output        cfg_en6060,
   output        cfg_en6061,
   output        cfg_en6062,
   output        cfg_en6063,
   output        cfg_en6064,
   output        cfg_en6065,
   output        cfg_en6066,
   output        cfg_en6067,
   output        cfg_en6068,
   output        cfg_en6069,
   output        cfg_en6070,
   output        cfg_en6071,
   output        cfg_en6072,
   output        cfg_en6073,
   output        cfg_en6074,
   output        cfg_en6075,
   output        cfg_en6076,
   output        cfg_en6077,
   output        cfg_en6078,
   output        cfg_en6079,
   output        cfg_en6080,
   output        cfg_en6081,
   output        cfg_en6082,
   output        cfg_en6083,
   output        cfg_en6084,
   output        cfg_en6085,
   output        cfg_en6086,
   output        cfg_en6087,
   output        cfg_en6088,
   output        cfg_en6089,
   output        cfg_en6090,
   output        cfg_en6091,
   output        cfg_en6092,
   output        cfg_en6093,
   output        cfg_en6094,
   output        cfg_en6095,
   output        cfg_en6096,
   output        cfg_en6097,
   output        cfg_en6098,
   output        cfg_en6099,
   output        cfg_en6100,
   output        cfg_en6101,
   output        cfg_en6102,
   output        cfg_en6103,
   output        cfg_en6104,
   output        cfg_en6105,
   output        cfg_en6106,
   output        cfg_en6107,
   output        cfg_en6108,
   output        cfg_en6109,
   output        cfg_en6110,
   output        cfg_en6111,
   output        cfg_en6112,
   output        cfg_en6113,
   output        cfg_en6114,
   output        cfg_en6115,
   output        cfg_en6116,
   output        cfg_en6117,
   output        cfg_en6118,
   output        cfg_en6119,
   output        cfg_en6120,
   output        cfg_en6121,
   output        cfg_en6122,
   output        cfg_en6123,
   output        cfg_en6124,
   output        cfg_en6125,
   output        cfg_en6126,
   output        cfg_en6127,
   output        cfg_en6128,
   output        cfg_en6129,
   output        cfg_en6130,
   output        cfg_en6131,
   output        cfg_en6132,
   output        cfg_en6133,
   output        cfg_en6134,
   output        cfg_en6135,
   output        cfg_en6136,
   output        cfg_en6137,
   output        cfg_en6138,
   output        cfg_en6139,
   output        cfg_en6140,
   output        cfg_en6141,
   output        cfg_en6142,
   output        cfg_en6143,
   output        cfg_en6144,
   output        cfg_en6145,
   output        cfg_en6146,
   output        cfg_en6147,
   output        cfg_en6148,
   output        cfg_en6149,
   output        cfg_en6150,
   output        cfg_en6151,
   output        cfg_en6152,
   output        cfg_en6153,
   output        cfg_en6154,
   output        cfg_en6155,
   output        cfg_en6156,
   output        cfg_en6157,
   output        cfg_en6158,
   output        cfg_en6159,
   output        cfg_en6160,
   output        cfg_en6161,
   output        cfg_en6162,
   output        cfg_en6163,
   output        cfg_en6164,
   output        cfg_en6165,
   output        cfg_en6166,
   output        cfg_en6167,
   output        cfg_en6168,
   output        cfg_en6169,
   output        cfg_en6170,
   output        cfg_en6171,
   output        cfg_en6172,
   output        cfg_en6173,
   output        cfg_en6174,
   output        cfg_en6175,
   output        cfg_en6176,
   output        cfg_en6177,
   output        cfg_en6178,
   output        cfg_en6179,
   output        cfg_en6180,
   output        cfg_en6181,
   output        cfg_en6182,
   output        cfg_en6183,
   output        cfg_en6184,
   output        cfg_en6185,
   output        cfg_en6186,
   output        cfg_en6187,
   output        cfg_en6188,
   output        cfg_en6189,
   output        cfg_en6190,
   output        cfg_en6191,
   output        cfg_en6192,
   output        cfg_en6193,
   output        cfg_en6194,
   output        cfg_en6195,
   output        cfg_en6196,
   output        cfg_en6197,
   output        cfg_en6198,
   output        cfg_en6199,
   output        cfg_en6200,
   output        cfg_en6201,
   output        cfg_en6202,
   output        cfg_en6203,
   output        cfg_en6204,
   output        cfg_en6205,
   output        cfg_en6206,
   output        cfg_en6207,
   output        cfg_en6208,
   output        cfg_en6209,
   output        cfg_en6210,
   output        cfg_en6211,
   output        cfg_en6212,
   output        cfg_en6213,
   output        cfg_en6214,
   output        cfg_en6215,
   output        cfg_en6216,
   output        cfg_en6217,
   output        cfg_en6218,
   output        cfg_en6219,
   output        cfg_en6220,
   output        cfg_en6221,
   output        cfg_en6222,
   output        cfg_en6223,
   output        cfg_en6224,
   output        cfg_en6225,
   output        cfg_en6226,
   output        cfg_en6227,
   output        cfg_en6228,
   output        cfg_en6229,
   output        cfg_en6230,
   output        cfg_en6231,
   output        cfg_en6232,
   output        cfg_en6233,
   output        cfg_en6234,
   output        cfg_en6235,
   output        cfg_en6236,
   output        cfg_en6237,
   output        cfg_en6238,
   output        cfg_en6239,
   output        cfg_en6240,
   output        cfg_en6241,
   output        cfg_en6242,
   output        cfg_en6243,
   output        cfg_en6244,
   output        cfg_en6245,
   output        cfg_en6246,
   output        cfg_en6247,
   output        cfg_en6248,
   output        cfg_en6249,
   output        cfg_en6250,
   output        cfg_en6251,
   output        cfg_en6252,
   output        cfg_en6253,
   output        cfg_en6254,
   output        cfg_en6255,
   output        cfg_en6256,
   output        cfg_en6257,
   output        cfg_en6258,
   output        cfg_en6259,
   output        cfg_en6260,
   output        cfg_en6261,
   output        cfg_en6262,
   output        cfg_en6263,
   output        cfg_en6264,
   output        cfg_en6265,
   output        cfg_en6266,
   output        cfg_en6267,
   output        cfg_en6268,
   output        cfg_en6269,
   output        cfg_en6270,
   output        cfg_en6271,
   output        cfg_en6272,
   output        cfg_en6273,
   output        cfg_en6274,
   output        cfg_en6275,
   output        cfg_en6276,
   output        cfg_en6277,
   output        cfg_en6278,
   output        cfg_en6279,
   output        cfg_en6280,
   output        cfg_en6281,
   output        cfg_en6282,
   output        cfg_en6283,
   output        cfg_en6284,
   output        cfg_en6285,
   output        cfg_en6286,
   output        cfg_en6287,
   output        cfg_en6288,
   output        cfg_en6289,
   output        cfg_en6290,
   output        cfg_en6291,
   output        cfg_en6292,
   output        cfg_en6293,
   output        cfg_en6294,
   output        cfg_en6295,
   output        cfg_en6296,
   output        cfg_en6297,
   output        cfg_en6298,
   output        cfg_en6299,
   output        cfg_en6300,
   output        cfg_en6301,
   output        cfg_en6302,
   output        cfg_en6303,
   output        cfg_en6304,
   output        cfg_en6305,
   output        cfg_en6306,
   output        cfg_en6307,
   output        cfg_en6308,
   output        cfg_en6309,
   output        cfg_en6310,
   output        cfg_en6311,
   output        cfg_en6312,
   output        cfg_en6313,
   output        cfg_en6314,
   output        cfg_en6315,
   output        cfg_en6316,
   output        cfg_en6317,
   output        cfg_en6318,
   output        cfg_en6319,
   output        cfg_en6320,
   output        cfg_en6321,
   output        cfg_en6322,
   output        cfg_en6323,
   output        cfg_en6324,
   output        cfg_en6325,
   output        cfg_en6326,
   output        cfg_en6327,
   output        cfg_en6328,
   output        cfg_en6329,
   output        cfg_en6330,
   output        cfg_en6331,
   output        cfg_en6332,
   output        cfg_en6333,
   output        cfg_en6334,
   output        cfg_en6335,
   output        cfg_en6336,
   output        cfg_en6337,
   output        cfg_en6338,
   output        cfg_en6339,
   output        cfg_en6340,
   output        cfg_en6341,
   output        cfg_en6342,
   output        cfg_en6343,
   output        cfg_en6344,
   output        cfg_en6345,
   output        cfg_en6346,
   output        cfg_en6347,
   output        cfg_en6348,
   output        cfg_en6349,
   output        cfg_en6350,
   output        cfg_en6351,
   output        cfg_en6352,
   output        cfg_en6353,
   output        cfg_en6354,
   output        cfg_en6355,
   output        cfg_en6356,
   output        cfg_en6357,
   output        cfg_en6358,
   output        cfg_en6359,
   output        cfg_en6360,
   output        cfg_en6361,
   output        cfg_en6362,
   output        cfg_en6363,
   output        cfg_en6364,
   output        cfg_en6365,
   output        cfg_en6366,
   output        cfg_en6367,
   output        cfg_en6368,
   output        cfg_en6369,
   output        cfg_en6370,
   output        cfg_en6371,
   output        cfg_en6372,
   output        cfg_en6373,
   output        cfg_en6374,
   output        cfg_en6375,
   output        cfg_en6376,
   output        cfg_en6377,
   output        cfg_en6378,
   output        cfg_en6379,
   output        cfg_en6380,
   output        cfg_en6381,
   output        cfg_en6382,
   output        cfg_en6383,
   output        cfg_en6384,
   output        cfg_en6385,
   output        cfg_en6386,
   output        cfg_en6387,
   output        cfg_en6388,
   output        cfg_en6389,
   output        cfg_en6390,
   output        cfg_en6391,
   output        cfg_en6392,
   output        cfg_en6393,
   output        cfg_en6394,
   output        cfg_en6395,
   output        cfg_en6396,
   output        cfg_en6397,
   output        cfg_en6398,
   output        cfg_en6399,
   output        cfg_en6400,
   output        cfg_en6401,
   output        cfg_en6402,
   output        cfg_en6403,
   output        cfg_en6404,
   output        cfg_en6405,
   output        cfg_en6406,
   output        cfg_en6407,
   output        cfg_en6408,
   output        cfg_en6409,
   output        cfg_en6410,
   output        cfg_en6411,
   output        cfg_en6412,
   output        cfg_en6413,
   output        cfg_en6414,
   output        cfg_en6415,
   output        cfg_en6416,
   output        cfg_en6417,
   output        cfg_en6418,
   output        cfg_en6419,
   output        cfg_en6420,
   output        cfg_en6421,
   output        cfg_en6422,
   output        cfg_en6423,
   output        cfg_en6424,
   output        cfg_en6425,
   output        cfg_en6426,
   output        cfg_en6427,
   output        cfg_en6428,
   output        cfg_en6429,
   output        cfg_en6430,
   output        cfg_en6431,
   output        cfg_en6432,
   output        cfg_en6433,
   output        cfg_en6434,
   output        cfg_en6435,
   output        cfg_en6436,
   output        cfg_en6437,
   output        cfg_en6438,
   output        cfg_en6439,
   output        cfg_en6440,
   output        cfg_en6441,
   output        cfg_en6442,
   output        cfg_en6443,
   output        cfg_en6444,
   output        cfg_en6445,
   output        cfg_en6446,
   output        cfg_en6447,
   output        cfg_en6448,
   output        cfg_en6449,
   output        cfg_en6450,
   output        cfg_en6451,
   output        cfg_en6452,
   output        cfg_en6453,
   output        cfg_en6454,
   output        cfg_en6455,
   output        cfg_en6456,
   output        cfg_en6457,
   output        cfg_en6458,
   output        cfg_en6459,
   output        cfg_en6460,
   output        cfg_en6461,
   output        cfg_en6462,
   output        cfg_en6463,
   output        cfg_en6464,
   output        cfg_en6465,
   output        cfg_en6466,
   output        cfg_en6467,
   output        cfg_en6468,
   output        cfg_en6469,
   output        cfg_en6470,
   output        cfg_en6471,
   output        cfg_en6472,
   output        cfg_en6473,
   output        cfg_en6474,
   output        cfg_en6475,
   output        cfg_en6476,
   output        cfg_en6477,
   output        cfg_en6478,
   output        cfg_en6479,
   output        cfg_en6480,
   output        cfg_en6481,
   output        cfg_en6482,
   output        cfg_en6483,
   output        cfg_en6484,
   output        cfg_en6485,
   output        cfg_en6486,
   output        cfg_en6487,
   output        cfg_en6488,
   output        cfg_en6489,
   output        cfg_en6490,
   output        cfg_en6491,
   output        cfg_en6492,
   output        cfg_en6493,
   output        cfg_en6494,
   output        cfg_en6495,
   output        cfg_en6496,
   output        cfg_en6497,
   output        cfg_en6498,
   output        cfg_en6499,
   output        cfg_en6500,
   output        cfg_en6501,
   output        cfg_en6502,
   output        cfg_en6503,
   output        cfg_en6504,
   output        cfg_en6505,
   output        cfg_en6506,
   output        cfg_en6507,
   output        cfg_en6508,
   output        cfg_en6509,
   output        cfg_en6510,
   output        cfg_en6511,
   output        cfg_en6512,
   output        cfg_en6513,
   output        cfg_en6514,
   output        cfg_en6515,
   output        cfg_en6516,
   output        cfg_en6517,
   output        cfg_en6518,
   output        cfg_en6519,
   output        cfg_en6520,
   output        cfg_en6521,
   output        cfg_en6522,
   output        cfg_en6523,
   output        cfg_en6524,
   output        cfg_en6525,
   output        cfg_en6526,
   output        cfg_en6527,
   output        cfg_en6528,
   output        cfg_en6529,
   output        cfg_en6530,
   output        cfg_en6531,
   output        cfg_en6532,
   output        cfg_en6533,
   output        cfg_en6534,
   output        cfg_en6535,
   output        cfg_en6536,
   output        cfg_en6537,
   output        cfg_en6538,
   output        cfg_en6539,
   output        cfg_en6540,
   output        cfg_en6541,
   output        cfg_en6542,
   output        cfg_en6543,
   output        cfg_en6544,
   output        cfg_en6545,
   output        cfg_en6546,
   output        cfg_en6547,
   output        cfg_en6548,
   output        cfg_en6549,
   output        cfg_en6550,
   output        cfg_en6551,
   output        cfg_en6552,
   output        cfg_en6553,
   output        cfg_en6554,
   output        cfg_en6555,
   output        cfg_en6556,
   output        cfg_en6557,
   output        cfg_en6558,
   output        cfg_en6559,
   output        cfg_en6560,
   output        cfg_en6561,
   output        cfg_en6562,
   output        cfg_en6563,
   output        cfg_en6564,
   output        cfg_en6565,
   output        cfg_en6566,
   output        cfg_en6567,
   output        cfg_en6568,
   output        cfg_en6569,
   output        cfg_en6570,
   output        cfg_en6571,
   output        cfg_en6572,
   output        cfg_en6573,
   output        cfg_en6574,
   output        cfg_en6575,
   output        cfg_en6576,
   output        cfg_en6577,
   output        cfg_en6578,
   output        cfg_en6579,
   output        cfg_en6580,
   output        cfg_en6581,
   output        cfg_en6582,
   output        cfg_en6583,
   output        cfg_en6584,
   output        cfg_en6585,
   output        cfg_en6586,
   output        cfg_en6587,
   output        cfg_en6588,
   output        cfg_en6589,
   output        cfg_en6590,
   output        cfg_en6591,
   output        cfg_en6592,
   output        cfg_en6593,
   output        cfg_en6594,
   output        cfg_en6595,
   output        cfg_en6596,
   output        cfg_en6597,
   output        cfg_en6598,
   output        cfg_en6599,
   output        cfg_en6600,
   output        cfg_en6601,
   output        cfg_en6602,
   output        cfg_en6603,
   output        cfg_en6604,
   output        cfg_en6605,
   output        cfg_en6606,
   output        cfg_en6607,
   output        cfg_en6608,
   output        cfg_en6609,
   output        cfg_en6610,
   output        cfg_en6611,
   output        cfg_en6612,
   output        cfg_en6613,
   output        cfg_en6614,
   output        cfg_en6615,
   output        cfg_en6616,
   output        cfg_en6617,
   output        cfg_en6618,
   output        cfg_en6619,
   output        cfg_en6620,
   output        cfg_en6621,
   output        cfg_en6622,
   output        cfg_en6623,
   output        cfg_en6624,
   output        cfg_en6625,
   output        cfg_en6626,
   output        cfg_en6627,
   output        cfg_en6628,
   output        cfg_en6629,
   output        cfg_en6630,
   output        cfg_en6631,
   output        cfg_en6632,
   output        cfg_en6633,
   output        cfg_en6634,
   output        cfg_en6635,
   output        cfg_en6636,
   output        cfg_en6637,
   output        cfg_en6638,
   output        cfg_en6639,
   output        cfg_en6640,
   output        cfg_en6641,
   output        cfg_en6642,
   output        cfg_en6643,
   output        cfg_en6644,
   output        cfg_en6645,
   output        cfg_en6646,
   output        cfg_en6647,
   output        cfg_en6648,
   output        cfg_en6649,
   output        cfg_en6650,
   output        cfg_en6651,
   output        cfg_en6652,
   output        cfg_en6653,
   output        cfg_en6654,
   output        cfg_en6655,
   output        cfg_en6656,
   output        cfg_en6657,
   output        cfg_en6658,
   output        cfg_en6659,
   output        cfg_en6660,
   output        cfg_en6661,
   output        cfg_en6662,
   output        cfg_en6663,
   output        cfg_en6664,
   output        cfg_en6665,
   output        cfg_en6666,
   output        cfg_en6667,
   output        cfg_en6668,
   output        cfg_en6669,
   output        cfg_en6670,
   output        cfg_en6671,
   output        cfg_en6672,
   output        cfg_en6673,
   output        cfg_en6674,
   output        cfg_en6675,
   output        cfg_en6676,
   output        cfg_en6677,
   output        cfg_en6678,
   output        cfg_en6679,
   output        cfg_en6680,
   output        cfg_en6681,
   output        cfg_en6682,
   output        cfg_en6683,
   output        cfg_en6684,
   output        cfg_en6685,
   output        cfg_en6686,
   output        cfg_en6687,
   output        cfg_en6688,
   output        cfg_en6689,
   output        cfg_en6690,
   output        cfg_en6691,
   output        cfg_en6692,
   output        cfg_en6693,
   output        cfg_en6694,
   output        cfg_en6695,
   output        cfg_en6696,
   output        cfg_en6697,
   output        cfg_en6698,
   output        cfg_en6699,
   output        cfg_en6700,
   output        cfg_en6701,
   output        cfg_en6702,
   output        cfg_en6703,
   output        cfg_en6704,
   output        cfg_en6705,
   output        cfg_en6706,
   output        cfg_en6707,
   output        cfg_en6708,
   output        cfg_en6709,
   output        cfg_en6710,
   output        cfg_en6711,
   output        cfg_en6712,
   output        cfg_en6713,
   output        cfg_en6714,
   output        cfg_en6715,
   output        cfg_en6716,
   output        cfg_en6717,
   output        cfg_en6718,
   output        cfg_en6719,
   output        cfg_en6720,
   output        cfg_en6721,
   output        cfg_en6722,
   output        cfg_en6723,
   output        cfg_en6724,
   output        cfg_en6725,
   output        cfg_en6726,
   output        cfg_en6727,
   output        cfg_en6728,
   output        cfg_en6729,
   output        cfg_en6730,
   output        cfg_en6731,
   output        cfg_en6732,
   output        cfg_en6733,
   output        cfg_en6734,
   output        cfg_en6735,
   output        cfg_en6736,
   output        cfg_en6737,
   output        cfg_en6738,
   output        cfg_en6739,
   output        cfg_en6740,
   output        cfg_en6741,
   output        cfg_en6742,
   output        cfg_en6743,
   output        cfg_en6744,
   output        cfg_en6745,
   output        cfg_en6746,
   output        cfg_en6747,
   output        cfg_en6748,
   output        cfg_en6749,
   output        cfg_en6750,
   output        cfg_en6751,
   output        cfg_en6752,
   output        cfg_en6753,
   output        cfg_en6754,
   output        cfg_en6755,
   output        cfg_en6756,
   output        cfg_en6757,
   output        cfg_en6758,
   output        cfg_en6759,
   output        cfg_en6760,
   output        cfg_en6761,
   output        cfg_en6762,
   output        cfg_en6763,
   output        cfg_en6764,
   output        cfg_en6765,
   output        cfg_en6766,
   output        cfg_en6767,
   output        cfg_en6768,
   output        cfg_en6769,
   output        cfg_en6770,
   output        cfg_en6771,
   output        cfg_en6772,
   output        cfg_en6773,
   output        cfg_en6774,
   output        cfg_en6775,
   output        cfg_en6776,
   output        cfg_en6777,
   output        cfg_en6778,
   output        cfg_en6779,
   output        cfg_en6780,
   output        cfg_en6781,
   output        cfg_en6782,
   output        cfg_en6783,
   output        cfg_en6784,
   output        cfg_en6785,
   output        cfg_en6786,
   output        cfg_en6787,
   output        cfg_en6788,
   output        cfg_en6789,
   output        cfg_en6790,
   output        cfg_en6791,
   output        cfg_en6792,
   output        cfg_en6793,
   output        cfg_en6794,
   output        cfg_en6795,
   output        cfg_en6796,
   output        cfg_en6797,
   output        cfg_en6798,
   output        cfg_en6799,
   output        cfg_en6800,
   output        cfg_en6801,
   output        cfg_en6802,
   output        cfg_en6803,
   output        cfg_en6804,
   output        cfg_en6805,
   output        cfg_en6806,
   output        cfg_en6807,
   output        cfg_en6808,
   output        cfg_en6809,
   output        cfg_en6810,
   output        cfg_en6811,
   output        cfg_en6812,
   output        cfg_en6813,
   output        cfg_en6814,
   output        cfg_en6815,
   output        cfg_en6816,
   output        cfg_en6817,
   output        cfg_en6818,
   output        cfg_en6819,
   output        cfg_en6820,
   output        cfg_en6821,
   output        cfg_en6822,
   output        cfg_en6823,
   output        cfg_en6824,
   output        cfg_en6825,
   output        cfg_en6826,
   output        cfg_en6827,
   output        cfg_en6828,
   output        cfg_en6829,
   output        cfg_en6830,
   output        cfg_en6831,
   output        cfg_en6832,
   output        cfg_en6833,
   output        cfg_en6834,
   output        cfg_en6835,
   output        cfg_en6836,
   output        cfg_en6837,
   output        cfg_en6838,
   output        cfg_en6839,
   output        cfg_en6840,
   output        cfg_en6841,
   output        cfg_en6842,
   output        cfg_en6843,
   output        cfg_en6844,
   output        cfg_en6845,
   output        cfg_en6846,
   output        cfg_en6847,
   output        cfg_en6848,
   output        cfg_en6849,
   output        cfg_en6850,
   output        cfg_en6851,
   output        cfg_en6852,
   output        cfg_en6853,
   output        cfg_en6854,
   output        cfg_en6855,
   output        cfg_en6856,
   output        cfg_en6857,
   output        cfg_en6858,
   output        cfg_en6859,
   output        cfg_en6860,
   output        cfg_en6861,
   output        cfg_en6862,
   output        cfg_en6863,
   output        cfg_en6864,
   output        cfg_en6865,
   output        cfg_en6866,
   output        cfg_en6867,
   output        cfg_en6868,
   output        cfg_en6869,
   output        cfg_en6870,
   output        cfg_en6871,
   output        cfg_en6872,
   output        cfg_en6873,
   output        cfg_en6874,
   output        cfg_en6875,
   output        cfg_en6876,
   output        cfg_en6877,
   output        cfg_en6878,
   output        cfg_en6879,
   output        cfg_en6880,
   output        cfg_en6881,
   output        cfg_en6882,
   output        cfg_en6883,
   output        cfg_en6884,
   output        cfg_en6885,
   output        cfg_en6886,
   output        cfg_en6887,
   output        cfg_en6888,
   output        cfg_en6889,
   output        cfg_en6890,
   output        cfg_en6891,
   output        cfg_en6892,
   output        cfg_en6893,
   output        cfg_en6894,
   output        cfg_en6895,
   output        cfg_en6896,
   output        cfg_en6897,
   output        cfg_en6898,
   output        cfg_en6899,
   output        cfg_en6900,
   output        cfg_en6901,
   output        cfg_en6902,
   output        cfg_en6903,
   output        cfg_en6904,
   output        cfg_en6905,
   output        cfg_en6906,
   output        cfg_en6907,
   output        cfg_en6908,
   output        cfg_en6909,
   output        cfg_en6910,
   output        cfg_en6911,
   output        cfg_en6912,
   output        cfg_en6913,
   output        cfg_en6914,
   output        cfg_en6915,
   output        cfg_en6916,
   output        cfg_en6917,
   output        cfg_en6918,
   output        cfg_en6919,
   output        cfg_en6920,
   output        cfg_en6921,
   output        cfg_en6922,
   output        cfg_en6923,
   output        cfg_en6924,
   output        cfg_en6925,
   output        cfg_en6926,
   output        cfg_en6927,
   output        cfg_en6928,
   output        cfg_en6929,
   output        cfg_en6930,
   output        cfg_en6931,
   output        cfg_en6932,
   output        cfg_en6933,
   output        cfg_en6934,
   output        cfg_en6935,
   output        cfg_en6936,
   output        cfg_en6937,
   output        cfg_en6938,
   output        cfg_en6939,
   output        cfg_en6940,
   output        cfg_en6941,
   output        cfg_en6942,
   output        cfg_en6943,
   output        cfg_en6944,
   output        cfg_en6945,
   output        cfg_en6946,
   output        cfg_en6947,
   output        cfg_en6948,
   output        cfg_en6949,
   output        cfg_en6950,
   output        cfg_en6951,
   output        cfg_en6952,
   output        cfg_en6953,
   output        cfg_en6954,
   output        cfg_en6955,
   output        cfg_en6956,
   output        cfg_en6957,
   output        cfg_en6958,
   output        cfg_en6959,
   output        cfg_en6960,
   output        cfg_en6961,
   output        cfg_en6962,
   output        cfg_en6963,
   output        cfg_en6964,
   output        cfg_en6965,
   output        cfg_en6966,
   output        cfg_en6967,
   output        cfg_en6968,
   output        cfg_en6969,
   output        cfg_en6970,
   output        cfg_en6971,
   output        cfg_en6972,
   output        cfg_en6973,
   output        cfg_en6974,
   output        cfg_en6975,
   output        cfg_en6976,
   output        cfg_en6977,
   output        cfg_en6978,
   output        cfg_en6979,
   output        cfg_en6980,
   output        cfg_en6981,
   output        cfg_en6982,
   output        cfg_en6983,
   output        cfg_en6984,
   output        cfg_en6985,
   output        cfg_en6986,
   output        cfg_en6987,
   output        cfg_en6988,
   output        cfg_en6989,
   output        cfg_en6990,
   output        cfg_en6991,
   output        cfg_en6992,
   output        cfg_en6993,
   output        cfg_en6994,
   output        cfg_en6995,
   output        cfg_en6996,
   output        cfg_en6997,
   output        cfg_en6998,
   output        cfg_en6999,
   output        cfg_en7000,
   output        cfg_en7001,
   output        cfg_en7002,
   output        cfg_en7003,
   output        cfg_en7004,
   output        cfg_en7005,
   output        cfg_en7006,
   output        cfg_en7007,
   output        cfg_en7008,
   output        cfg_en7009,
   output        cfg_en7010,
   output        cfg_en7011,
   output        cfg_en7012,
   output        cfg_en7013,
   output        cfg_en7014,
   output        cfg_en7015,
   output        cfg_en7016,
   output        cfg_en7017,
   output        cfg_en7018,
   output        cfg_en7019,
   output        cfg_en7020,
   output        cfg_en7021,
   output        cfg_en7022,
   output        cfg_en7023,
   output        cfg_en7024,
   output        cfg_en7025,
   output        cfg_en7026,
   output        cfg_en7027,
   output        cfg_en7028,
   output        cfg_en7029,
   output        cfg_en7030,
   output        cfg_en7031,
   output        cfg_en7032,
   output        cfg_en7033,
   output        cfg_en7034,
   output        cfg_en7035,
   output        cfg_en7036,
   output        cfg_en7037,
   output        cfg_en7038,
   output        cfg_en7039,
   output        cfg_en7040,
   output        cfg_en7041,
   output        cfg_en7042,
   output        cfg_en7043,
   output        cfg_en7044,
   output        cfg_en7045,
   output        cfg_en7046,
   output        cfg_en7047,
   output        cfg_en7048,
   output        cfg_en7049,
   output        cfg_en7050,
   output        cfg_en7051,
   output        cfg_en7052,
   output        cfg_en7053,
   output        cfg_en7054,
   output        cfg_en7055,
   output        cfg_en7056,
   output        cfg_en7057,
   output        cfg_en7058,
   output        cfg_en7059,
   output        cfg_en7060,
   output        cfg_en7061,
   output        cfg_en7062,
   output        cfg_en7063,
   output        cfg_en7064,
   output        cfg_en7065,
   output        cfg_en7066,
   output        cfg_en7067,
   output        cfg_en7068,
   output        cfg_en7069,
   output        cfg_en7070,
   output        cfg_en7071,
   output        cfg_en7072,
   output        cfg_en7073,
   output        cfg_en7074,
   output        cfg_en7075,
   output        cfg_en7076,
   output        cfg_en7077,
   output        cfg_en7078,
   output        cfg_en7079,
   output        cfg_en7080,
   output        cfg_en7081,
   output        cfg_en7082,
   output        cfg_en7083,
   output        cfg_en7084,
   output        cfg_en7085,
   output        cfg_en7086,
   output        cfg_en7087,
   output        cfg_en7088,
   output        cfg_en7089,
   output        cfg_en7090,
   output        cfg_en7091,
   output        cfg_en7092,
   output        cfg_en7093,
   output        cfg_en7094,
   output        cfg_en7095,
   output        cfg_en7096,
   output        cfg_en7097,
   output        cfg_en7098,
   output        cfg_en7099,
   output        cfg_en7100,
   output        cfg_en7101,
   output        cfg_en7102,
   output        cfg_en7103,
   output        cfg_en7104,
   output        cfg_en7105,
   output        cfg_en7106,
   output        cfg_en7107,
   output        cfg_en7108,
   output        cfg_en7109,
   output        cfg_en7110,
   output        cfg_en7111,
   output        cfg_en7112,
   output        cfg_en7113,
   output        cfg_en7114,
   output        cfg_en7115,
   output        cfg_en7116,
   output        cfg_en7117,
   output        cfg_en7118,
   output        cfg_en7119,
   output        cfg_en7120,
   output        cfg_en7121,
   output        cfg_en7122,
   output        cfg_en7123,
   output        cfg_en7124,
   output        cfg_en7125,
   output        cfg_en7126,
   output        cfg_en7127,
   output        cfg_en7128,
   output        cfg_en7129,
   output        cfg_en7130,
   output        cfg_en7131,
   output        cfg_en7132,
   output        cfg_en7133,
   output        cfg_en7134,
   output        cfg_en7135,
   output        cfg_en7136,
   output        cfg_en7137,
   output        cfg_en7138,
   output        cfg_en7139,
   output        cfg_en7140,
   output        cfg_en7141,
   output        cfg_en7142,
   output        cfg_en7143,
   output        cfg_en7144,
   output        cfg_en7145,
   output        cfg_en7146,
   output        cfg_en7147,
   output        cfg_en7148,
   output        cfg_en7149,
   output        cfg_en7150,
   output        cfg_en7151,
   output        cfg_en7152,
   output        cfg_en7153,
   output        cfg_en7154,
   output        cfg_en7155,
   output        cfg_en7156,
   output        cfg_en7157,
   output        cfg_en7158,
   output        cfg_en7159,
   output        cfg_en7160,
   output        cfg_en7161,
   output        cfg_en7162,
   output        cfg_en7163,
   output        cfg_en7164,
   output        cfg_en7165,
   output        cfg_en7166,
   output        cfg_en7167,
   output        cfg_en7168,
   output        cfg_en7169,
   output        cfg_en7170,
   output        cfg_en7171,
   output        cfg_en7172,
   output        cfg_en7173,
   output        cfg_en7174,
   output        cfg_en7175,
   output        cfg_en7176,
   output        cfg_en7177,
   output        cfg_en7178,
   output        cfg_en7179,
   output        cfg_en7180,
   output        cfg_en7181,
   output        cfg_en7182,
   output        cfg_en7183,
   output        cfg_en7184,
   output        cfg_en7185,
   output        cfg_en7186,
   output        cfg_en7187,
   output        cfg_en7188,
   output        cfg_en7189,
   output        cfg_en7190,
   output        cfg_en7191,
   output        cfg_en7192,
   output        cfg_en7193,
   output        cfg_en7194,
   output        cfg_en7195,
   output        cfg_en7196,
   output        cfg_en7197,
   output        cfg_en7198,
   output        cfg_en7199,
   output        cfg_en7200,
   output        cfg_en7201,
   output        cfg_en7202,
   output        cfg_en7203,
   output        cfg_en7204,
   output        cfg_en7205,
   output        cfg_en7206,
   output        cfg_en7207,
   output        cfg_en7208,
   output        cfg_en7209,
   output        cfg_en7210,
   output        cfg_en7211,
   output        cfg_en7212,
   output        cfg_en7213,
   output        cfg_en7214,
   output        cfg_en7215,
   output        cfg_en7216,
   output        cfg_en7217,
   output        cfg_en7218,
   output        cfg_en7219,
   output        cfg_en7220,
   output        cfg_en7221,
   output        cfg_en7222,
   output        cfg_en7223,
   output        cfg_en7224,
   output        cfg_en7225,
   output        cfg_en7226,
   output        cfg_en7227,
   output        cfg_en7228,
   output        cfg_en7229,
   output        cfg_en7230,
   output        cfg_en7231,
   output        cfg_en7232,
   output        cfg_en7233,
   output        cfg_en7234,
   output        cfg_en7235,
   output        cfg_en7236,
   output        cfg_en7237,
   output        cfg_en7238,
   output        cfg_en7239,
   output        cfg_en7240,
   output        cfg_en7241,
   output        cfg_en7242,
   output        cfg_en7243,
   output        cfg_en7244,
   output        cfg_en7245,
   output        cfg_en7246,
   output        cfg_en7247,
   output        cfg_en7248,
   output        cfg_en7249,
   output        cfg_en7250,
   output        cfg_en7251,
   output        cfg_en7252,
   output        cfg_en7253,
   output        cfg_en7254,
   output        cfg_en7255,
   output        cfg_en7256,
   output        cfg_en7257,
   output        cfg_en7258,
   output        cfg_en7259,
   output        cfg_en7260,
   output        cfg_en7261,
   output        cfg_en7262,
   output        cfg_en7263,
   output        cfg_en7264,
   output        cfg_en7265,
   output        cfg_en7266,
   output        cfg_en7267,
   output        cfg_en7268,
   output        cfg_en7269,
   output        cfg_en7270,
   output        cfg_en7271,
   output        cfg_en7272,
   output        cfg_en7273,
   output        cfg_en7274,
   output        cfg_en7275,
   output        cfg_en7276,
   output        cfg_en7277,
   output        cfg_en7278,
   output        cfg_en7279,
   output        cfg_en7280,
   output        cfg_en7281,
   output        cfg_en7282,
   output        cfg_en7283,
   output        cfg_en7284,
   output        cfg_en7285,
   output        cfg_en7286,
   output        cfg_en7287,
   output        cfg_en7288,
   output        cfg_en7289,
   output        cfg_en7290,
   output        cfg_en7291,
   output        cfg_en7292,
   output        cfg_en7293,
   output        cfg_en7294,
   output        cfg_en7295,
   output        cfg_en7296,
   output        cfg_en7297,
   output        cfg_en7298,
   output        cfg_en7299,
   output        cfg_en7300,
   output        cfg_en7301,
   output        cfg_en7302,
   output        cfg_en7303,
   output        cfg_en7304,
   output        cfg_en7305,
   output        cfg_en7306,
   output        cfg_en7307,
   output        cfg_en7308,
   output        cfg_en7309,
   output        cfg_en7310,
   output        cfg_en7311,
   output        cfg_en7312,
   output        cfg_en7313,
   output        cfg_en7314,
   output        cfg_en7315,
   output        cfg_en7316,
   output        cfg_en7317,
   output        cfg_en7318,
   output        cfg_en7319,
   output        cfg_en7320,
   output        cfg_en7321,
   output        cfg_en7322,
   output        cfg_en7323,
   output        cfg_en7324,
   output        cfg_en7325,
   output        cfg_en7326,
   output        cfg_en7327,
   output        cfg_en7328,
   output        cfg_en7329,
   output        cfg_en7330,
   output        cfg_en7331,
   output        cfg_en7332,
   output        cfg_en7333,
   output        cfg_en7334,
   output        cfg_en7335,
   output        cfg_en7336,
   output        cfg_en7337,
   output        cfg_en7338,
   output        cfg_en7339,
   output        cfg_en7340,
   output        cfg_en7341,
   output        cfg_en7342,
   output        cfg_en7343,
   output        cfg_en7344,
   output        cfg_en7345,
   output        cfg_en7346,
   output        cfg_en7347,
   output        cfg_en7348,
   output        cfg_en7349,
   output        cfg_en7350,
   output        cfg_en7351,
   output        cfg_en7352,
   output        cfg_en7353,
   output        cfg_en7354,
   output        cfg_en7355,
   output        cfg_en7356,
   output        cfg_en7357,
   output        cfg_en7358,
   output        cfg_en7359,
   output        cfg_en7360,
   output        cfg_en7361,
   output        cfg_en7362,
   output        cfg_en7363,
   output        cfg_en7364,
   output        cfg_en7365,
   output        cfg_en7366,
   output        cfg_en7367,
   output        cfg_en7368,
   output        cfg_en7369,
   output        cfg_en7370,
   output        cfg_en7371,
   output        cfg_en7372,
   output        cfg_en7373,
   output        cfg_en7374,
   output        cfg_en7375,
   output        cfg_en7376,
   output        cfg_en7377,
   output        cfg_en7378,
   output        cfg_en7379,
   output        cfg_en7380,
   output        cfg_en7381,
   output        cfg_en7382,
   output        cfg_en7383,
   output        cfg_en7384,
   output        cfg_en7385,
   output        cfg_en7386,
   output        cfg_en7387,
   output        cfg_en7388,
   output        cfg_en7389,
   output        cfg_en7390,
   output        cfg_en7391,
   output        cfg_en7392,
   output        cfg_en7393,
   output        cfg_en7394,
   output        cfg_en7395,
   output        cfg_en7396,
   output        cfg_en7397,
   output        cfg_en7398,
   output        cfg_en7399,
   output        cfg_en7400,
   output        cfg_en7401,
   output        cfg_en7402,
   output        cfg_en7403,
   output        cfg_en7404,
   output        cfg_en7405,
   output        cfg_en7406,
   output        cfg_en7407,
   output        cfg_en7408,
   output        cfg_en7409,
   output        cfg_en7410,
   output        cfg_en7411,
   output        cfg_en7412,
   output        cfg_en7413,
   output        cfg_en7414,
   output        cfg_en7415,
   output        cfg_en7416,
   output        cfg_en7417,
   output        cfg_en7418,
   output        cfg_en7419,
   output        cfg_en7420,
   output        cfg_en7421,
   output        cfg_en7422,
   output        cfg_en7423,
   output        cfg_en7424,
   output        cfg_en7425,
   output        cfg_en7426,
   output        cfg_en7427,
   output        cfg_en7428,
   output        cfg_en7429,
   output        cfg_en7430,
   output        cfg_en7431,
   output        cfg_en7432,
   output        cfg_en7433,
   output        cfg_en7434,
   output        cfg_en7435,
   output        cfg_en7436,
   output        cfg_en7437,
   output        cfg_en7438,
   output        cfg_en7439,
   output        cfg_en7440,
   output        cfg_en7441,
   output        cfg_en7442,
   output        cfg_en7443,
   output        cfg_en7444,
   output        cfg_en7445,
   output        cfg_en7446,
   output        cfg_en7447,
   output        cfg_en7448,
   output        cfg_en7449,
   output        cfg_en7450,
   output        cfg_en7451,
   output        cfg_en7452,
   output        cfg_en7453,
   output        cfg_en7454,
   output        cfg_en7455,
   output        cfg_en7456,
   output        cfg_en7457,
   output        cfg_en7458,
   output        cfg_en7459,
   output        cfg_en7460,
   output        cfg_en7461,
   output        cfg_en7462,
   output        cfg_en7463,
   output        cfg_en7464,
   output        cfg_en7465,
   output        cfg_en7466,
   output        cfg_en7467,
   output        cfg_en7468,
   output        cfg_en7469,
   output        cfg_en7470,
   output        cfg_en7471,
   output        cfg_en7472,
   output        cfg_en7473,
   output        cfg_en7474,
   output        cfg_en7475,
   output        cfg_en7476,
   output        cfg_en7477,
   output        cfg_en7478,
   output        cfg_en7479,
   output        cfg_en7480,
   output        cfg_en7481,
   output        cfg_en7482,
   output        cfg_en7483,
   output        cfg_en7484,
   output        cfg_en7485,
   output        cfg_en7486,
   output        cfg_en7487,
   output        cfg_en7488,
   output        cfg_en7489,
   output        cfg_en7490,
   output        cfg_en7491,
   output        cfg_en7492,
   output        cfg_en7493,
   output        cfg_en7494,
   output        cfg_en7495,
   output        cfg_en7496,
   output        cfg_en7497,
   output        cfg_en7498,
   output        cfg_en7499,
   output        cfg_en7500,
   output        cfg_en7501,
   output        cfg_en7502,
   output        cfg_en7503,
   output        cfg_en7504,
   output        cfg_en7505,
   output        cfg_en7506,
   output        cfg_en7507,
   output        cfg_en7508,
   output        cfg_en7509,
   output        cfg_en7510,
   output        cfg_en7511,
   output        cfg_en7512,
   output        cfg_en7513,
   output        cfg_en7514,
   output        cfg_en7515,
   output        cfg_en7516,
   output        cfg_en7517,
   output        cfg_en7518,
   output        cfg_en7519,
   output        cfg_en7520,
   output        cfg_en7521,
   output        cfg_en7522,
   output        cfg_en7523,
   output        cfg_en7524,
   output        cfg_en7525,
   output        cfg_en7526,
   output        cfg_en7527,
   output        cfg_en7528,
   output        cfg_en7529,
   output        cfg_en7530,
   output        cfg_en7531,
   output        cfg_en7532,
   output        cfg_en7533,
   output        cfg_en7534,
   output        cfg_en7535,
   output        cfg_en7536,
   output        cfg_en7537,
   output        cfg_en7538,
   output        cfg_en7539,
   output        cfg_en7540,
   output        cfg_en7541,
   output        cfg_en7542,
   output        cfg_en7543,
   output        cfg_en7544,
   output        cfg_en7545,
   output        cfg_en7546,
   output        cfg_en7547,
   output        cfg_en7548,
   output        cfg_en7549,
   output        cfg_en7550,
   output        cfg_en7551,
   output        cfg_en7552,
   output        cfg_en7553,
   output        cfg_en7554,
   output        cfg_en7555,
   output        cfg_en7556,
   output        cfg_en7557,
   output        cfg_en7558,
   output        cfg_en7559,
   output        cfg_en7560,
   output        cfg_en7561,
   output        cfg_en7562,
   output        cfg_en7563,
   output        cfg_en7564,
   output        cfg_en7565,
   output        cfg_en7566,
   output        cfg_en7567,
   output        cfg_en7568,
   output        cfg_en7569,
   output        cfg_en7570,
   output        cfg_en7571,
   output        cfg_en7572,
   output        cfg_en7573,
   output        cfg_en7574,
   output        cfg_en7575,
   output        cfg_en7576,
   output        cfg_en7577,
   output        cfg_en7578,
   output        cfg_en7579,
   output        cfg_en7580,
   output        cfg_en7581,
   output        cfg_en7582,
   output        cfg_en7583,
   output        cfg_en7584,
   output        cfg_en7585,
   output        cfg_en7586,
   output        cfg_en7587,
   output        cfg_en7588,
   output        cfg_en7589,
   output        cfg_en7590,
   output        cfg_en7591,
   output        cfg_en7592,
   output        cfg_en7593,
   output        cfg_en7594,
   output        cfg_en7595,
   output        cfg_en7596,
   output        cfg_en7597,
   output        cfg_en7598,
   output        cfg_en7599,
   output        cfg_en7600,
   output        cfg_en7601,
   output        cfg_en7602,
   output        cfg_en7603,
   output        cfg_en7604,
   output        cfg_en7605,
   output        cfg_en7606,
   output        cfg_en7607,
   output        cfg_en7608,
   output        cfg_en7609,
   output        cfg_en7610,
   output        cfg_en7611,
   output        cfg_en7612,
   output        cfg_en7613,
   output        cfg_en7614,
   output        cfg_en7615,
   output        cfg_en7616,
   output        cfg_en7617,
   output        cfg_en7618,
   output        cfg_en7619,
   output        cfg_en7620,
   output        cfg_en7621,
   output        cfg_en7622,
   output        cfg_en7623,
   output        cfg_en7624,
   output        cfg_en7625,
   output        cfg_en7626,
   output        cfg_en7627,
   output        cfg_en7628,
   output        cfg_en7629,
   output        cfg_en7630,
   output        cfg_en7631,
   output        cfg_en7632,
   output        cfg_en7633,
   output        cfg_en7634,
   output        cfg_en7635,
   output        cfg_en7636,
   output        cfg_en7637,
   output        cfg_en7638,
   output        cfg_en7639,
   output        cfg_en7640,
   output        cfg_en7641,
   output        cfg_en7642,
   output        cfg_en7643,
   output        cfg_en7644,
   output        cfg_en7645,
   output        cfg_en7646,
   output        cfg_en7647,
   output        cfg_en7648,
   output        cfg_en7649,
   output        cfg_en7650,
   output        cfg_en7651,
   output        cfg_en7652,
   output        cfg_en7653,
   output        cfg_en7654,
   output        cfg_en7655,
   output        cfg_en7656,
   output        cfg_en7657,
   output        cfg_en7658,
   output        cfg_en7659,
   output        cfg_en7660,
   output        cfg_en7661,
   output        cfg_en7662,
   output        cfg_en7663,
   output        cfg_en7664,
   output        cfg_en7665,
   output        cfg_en7666,
   output        cfg_en7667,
   output        cfg_en7668,
   output        cfg_en7669,
   output        cfg_en7670,
   output        cfg_en7671,
   output        cfg_en7672,
   output        cfg_en7673,
   output        cfg_en7674,
   output        cfg_en7675,
   output        cfg_en7676,
   output        cfg_en7677,
   output        cfg_en7678,
   output        cfg_en7679,
   output        cfg_en7680,
   output        cfg_en7681,
   output        cfg_en7682,
   output        cfg_en7683,
   output        cfg_en7684,
   output        cfg_en7685,
   output        cfg_en7686,
   output        cfg_en7687,
   output        cfg_en7688,
   output        cfg_en7689,
   output        cfg_en7690,
   output        cfg_en7691,
   output        cfg_en7692,
   output        cfg_en7693,
   output        cfg_en7694,
   output        cfg_en7695,
   output        cfg_en7696,
   output        cfg_en7697,
   output        cfg_en7698,
   output        cfg_en7699,
   output        cfg_en7700,
   output        cfg_en7701,
   output        cfg_en7702,
   output        cfg_en7703,
   output        cfg_en7704,
   output        cfg_en7705,
   output        cfg_en7706,
   output        cfg_en7707,
   output        cfg_en7708,
   output        cfg_en7709,
   output        cfg_en7710,
   output        cfg_en7711,
   output        cfg_en7712,
   output        cfg_en7713,
   output        cfg_en7714,
   output        cfg_en7715,
   output        cfg_en7716,
   output        cfg_en7717,
   output        cfg_en7718,
   output        cfg_en7719,
   output        cfg_en7720,
   output        cfg_en7721,
   output        cfg_en7722,
   output        cfg_en7723,
   output        cfg_en7724,
   output        cfg_en7725,
   output        cfg_en7726,
   output        cfg_en7727,
   output        cfg_en7728,
   output        cfg_en7729,
   output        cfg_en7730,
   output        cfg_en7731,
   output        cfg_en7732,
   output        cfg_en7733,
   output        cfg_en7734,
   output        cfg_en7735,
   output        cfg_en7736,
   output        cfg_en7737,
   output        cfg_en7738,
   output        cfg_en7739,
   output        cfg_en7740,
   output        cfg_en7741,
   output        cfg_en7742,
   output        cfg_en7743,
   output        cfg_en7744,
   output        cfg_en7745,
   output        cfg_en7746,
   output        cfg_en7747,
   output        cfg_en7748,
   output        cfg_en7749,
   output        cfg_en7750,
   output        cfg_en7751,
   output        cfg_en7752,
   output        cfg_en7753,
   output        cfg_en7754,
   output        cfg_en7755,
   output        cfg_en7756,
   output        cfg_en7757,
   output        cfg_en7758,
   output        cfg_en7759,
   output        cfg_en7760,
   output        cfg_en7761,
   output        cfg_en7762,
   output        cfg_en7763,
   output        cfg_en7764,
   output        cfg_en7765,
   output        cfg_en7766,
   output        cfg_en7767,
   output        cfg_en7768,
   output        cfg_en7769,
   output        cfg_en7770,
   output        cfg_en7771,
   output        cfg_en7772,
   output        cfg_en7773,
   output        cfg_en7774,
   output        cfg_en7775,
   output        cfg_en7776,
   output        cfg_en7777,
   output        cfg_en7778,
   output        cfg_en7779,
   output        cfg_en7780,
   output        cfg_en7781,
   output        cfg_en7782,
   output        cfg_en7783,
   output        cfg_en7784,
   output        cfg_en7785,
   output        cfg_en7786,
   output        cfg_en7787,
   output        cfg_en7788,
   output        cfg_en7789,
   output        cfg_en7790,
   output        cfg_en7791,
   output        cfg_en7792,
   output        cfg_en7793,
   output        cfg_en7794,
   output        cfg_en7795,
   output        cfg_en7796,
   output        cfg_en7797,
   output        cfg_en7798,
   output        cfg_en7799,
   output        cfg_en7800,
   output        cfg_en7801,
   output        cfg_en7802,
   output        cfg_en7803,
   output        cfg_en7804,
   output        cfg_en7805,
   output        cfg_en7806,
   output        cfg_en7807,
   output        cfg_en7808,
   output        cfg_en7809,
   output        cfg_en7810,
   output        cfg_en7811,
   output        cfg_en7812,
   output        cfg_en7813,
   output        cfg_en7814,
   output        cfg_en7815,
   output        cfg_en7816,
   output        cfg_en7817,
   output        cfg_en7818,
   output        cfg_en7819,
   output        cfg_en7820,
   output        cfg_en7821,
   output        cfg_en7822,
   output        cfg_en7823,
   output        cfg_en7824,
   output        cfg_en7825,
   output        cfg_en7826,
   output        cfg_en7827,
   output        cfg_en7828,
   output        cfg_en7829,
   output        cfg_en7830,
   output        cfg_en7831,
   output        cfg_en7832,
   output        cfg_en7833,
   output        cfg_en7834,
   output        cfg_en7835,
   output        cfg_en7836,
   output        cfg_en7837,
   output        cfg_en7838,
   output        cfg_en7839,
   output        cfg_en7840,
   output        cfg_en7841,
   output        cfg_en7842,
   output        cfg_en7843,
   output        cfg_en7844,
   output        cfg_en7845,
   output        cfg_en7846,
   output        cfg_en7847,
   output        cfg_en7848,
   output        cfg_en7849,
   output        cfg_en7850,
   output        cfg_en7851,
   output        cfg_en7852,
   output        cfg_en7853,
   output        cfg_en7854,
   output        cfg_en7855,
   output        cfg_en7856,
   output        cfg_en7857,
   output        cfg_en7858,
   output        cfg_en7859,
   output        cfg_en7860,
   output        cfg_en7861,
   output        cfg_en7862,
   output        cfg_en7863,
   output        cfg_en7864,
   output        cfg_en7865,
   output        cfg_en7866,
   output        cfg_en7867,
   output        cfg_en7868,
   output        cfg_en7869,
   output        cfg_en7870,
   output        cfg_en7871,
   output        cfg_en7872,
   output        cfg_en7873,
   output        cfg_en7874,
   output        cfg_en7875,
   output        cfg_en7876,
   output        cfg_en7877,
   output        cfg_en7878,
   output        cfg_en7879,
   output        cfg_en7880,
   output        cfg_en7881,
   output        cfg_en7882,
   output        cfg_en7883,
   output        cfg_en7884,
   output        cfg_en7885,
   output        cfg_en7886,
   output        cfg_en7887,
   output        cfg_en7888,
   output        cfg_en7889,
   output        cfg_en7890,
   output        cfg_en7891,
   output        cfg_en7892,
   output        cfg_en7893,
   output        cfg_en7894,
   output        cfg_en7895,
   output        cfg_en7896,
   output        cfg_en7897,
   output        cfg_en7898,
   output        cfg_en7899,
   output        cfg_en7900,
   output        cfg_en7901,
   output        cfg_en7902,
   output        cfg_en7903,
   output        cfg_en7904,
   output        cfg_en7905,
   output        cfg_en7906,
   output        cfg_en7907,
   output        cfg_en7908,
   output        cfg_en7909,
   output        cfg_en7910,
   output        cfg_en7911,
   output        cfg_en7912,
   output        cfg_en7913,
   output        cfg_en7914,
   output        cfg_en7915,
   output        cfg_en7916,
   output        cfg_en7917,
   output        cfg_en7918,
   output        cfg_en7919,
   output        cfg_en7920,
   output        cfg_en7921,
   output        cfg_en7922,
   output        cfg_en7923,
   output        cfg_en7924,
   output        cfg_en7925,
   output        cfg_en7926,
   output        cfg_en7927,
   output        cfg_en7928,
   output        cfg_en7929,
   output        cfg_en7930,
   output        cfg_en7931,
   output        cfg_en7932,
   output        cfg_en7933,
   output        cfg_en7934,
   output        cfg_en7935,
   output        cfg_en7936,
   output        cfg_en7937,
   output        cfg_en7938,
   output        cfg_en7939,
   output        cfg_en7940,
   output        cfg_en7941,
   output        cfg_en7942,
   output        cfg_en7943,
   output        cfg_en7944,
   output        cfg_en7945,
   output        cfg_en7946,
   output        cfg_en7947,
   output        cfg_en7948,
   output        cfg_en7949,
   output        cfg_en7950,
   output        cfg_en7951,
   output        cfg_en7952,
   output        cfg_en7953,
   output        cfg_en7954,
   output        cfg_en7955,
   output        cfg_en7956,
   output        cfg_en7957,
   output        cfg_en7958,
   output        cfg_en7959,
   output        cfg_en7960,
   output        cfg_en7961,
   output        cfg_en7962,
   output        cfg_en7963,
   output        cfg_en7964,
   output        cfg_en7965,
   output        cfg_en7966,
   output        cfg_en7967,
   output        cfg_en7968,
   output        cfg_en7969,
   output        cfg_en7970,
   output        cfg_en7971,
   output        cfg_en7972,
   output        cfg_en7973,
   output        cfg_en7974,
   output        cfg_en7975,
   output        cfg_en7976,
   output        cfg_en7977,
   output        cfg_en7978,
   output        cfg_en7979,
   output        cfg_en7980,
   output        cfg_en7981,
   output        cfg_en7982,
   output        cfg_en7983,
   output        cfg_en7984,
   output        cfg_en7985,
   output        cfg_en7986,
   output        cfg_en7987,
   output        cfg_en7988,
   output        cfg_en7989,
   output        cfg_en7990,
   output        cfg_en7991,
   output        cfg_en7992,
   output        cfg_en7993,
   output        cfg_en7994,
   output        cfg_en7995,
   output        cfg_en7996,
   output        cfg_en7997,
   output        cfg_en7998,
   output        cfg_en7999,
   output        cfg_en8000,
   output        cfg_en8001,
   output        cfg_en8002,
   output        cfg_en8003,
   output        cfg_en8004,
   output        cfg_en8005,
   output        cfg_en8006,
   output        cfg_en8007,
   output        cfg_en8008,
   output        cfg_en8009,
   output        cfg_en8010,
   output        cfg_en8011,
   output        cfg_en8012,
   output        cfg_en8013,
   output        cfg_en8014,
   output        cfg_en8015,
   output        cfg_en8016,
   output        cfg_en8017,
   output        cfg_en8018,
   output        cfg_en8019,
   output        cfg_en8020,
   output        cfg_en8021,
   output        cfg_en8022,
   output        cfg_en8023,
   output        cfg_en8024,
   output        cfg_en8025,
   output        cfg_en8026,
   output        cfg_en8027,
   output        cfg_en8028,
   output        cfg_en8029,
   output        cfg_en8030,
   output        cfg_en8031,
   output        cfg_en8032,
   output        cfg_en8033,
   output        cfg_en8034,
   output        cfg_en8035,
   output        cfg_en8036,
   output        cfg_en8037,
   output        cfg_en8038,
   output        cfg_en8039,
   output        cfg_en8040,
   output        cfg_en8041,
   output        cfg_en8042,
   output        cfg_en8043,
   output        cfg_en8044,
   output        cfg_en8045,
   output        cfg_en8046,
   output        cfg_en8047,
   output        cfg_en8048,
   output        cfg_en8049,
   output        cfg_en8050,
   output        cfg_en8051,
   output        cfg_en8052,
   output        cfg_en8053,
   output        cfg_en8054,
   output        cfg_en8055,
   output        cfg_en8056,
   output        cfg_en8057,
   output        cfg_en8058,
   output        cfg_en8059,
   output        cfg_en8060,
   output        cfg_en8061,
   output        cfg_en8062,
   output        cfg_en8063,
   output        cfg_en8064,
   output        cfg_en8065,
   output        cfg_en8066,
   output        cfg_en8067,
   output        cfg_en8068,
   output        cfg_en8069,
   output        cfg_en8070,
   output        cfg_en8071,
   output        cfg_en8072,
   output        cfg_en8073,
   output        cfg_en8074,
   output        cfg_en8075,
   output        cfg_en8076,
   output        cfg_en8077,
   output        cfg_en8078,
   output        cfg_en8079,
   output        cfg_en8080,
   output        cfg_en8081,
   output        cfg_en8082,
   output        cfg_en8083,
   output        cfg_en8084,
   output        cfg_en8085,
   output        cfg_en8086,
   output        cfg_en8087,
   output        cfg_en8088,
   output        cfg_en8089,
   output        cfg_en8090,
   output        cfg_en8091,
   output        cfg_en8092,
   output        cfg_en8093,
   output        cfg_en8094,
   output        cfg_en8095,
   output        cfg_en8096,
   output        cfg_en8097,
   output        cfg_en8098,
   output        cfg_en8099,
   output        cfg_en8100,
   output        cfg_en8101,
   output        cfg_en8102,
   output        cfg_en8103,
   output        cfg_en8104,
   output        cfg_en8105,
   output        cfg_en8106,
   output        cfg_en8107,
   output        cfg_en8108,
   output        cfg_en8109,
   output        cfg_en8110,
   output        cfg_en8111,
   output        cfg_en8112,
   output        cfg_en8113,
   output        cfg_en8114,
   output        cfg_en8115,
   output        cfg_en8116,
   output        cfg_en8117,
   output        cfg_en8118,
   output        cfg_en8119,
   output        cfg_en8120,
   output        cfg_en8121,
   output        cfg_en8122,
   output        cfg_en8123,
   output        cfg_en8124,
   output        cfg_en8125,
   output        cfg_en8126,
   output        cfg_en8127,
   output        cfg_en8128,
   output        cfg_en8129,
   output        cfg_en8130,
   output        cfg_en8131,
   output        cfg_en8132,
   output        cfg_en8133,
   output        cfg_en8134,
   output        cfg_en8135,
   output        cfg_en8136,
   output        cfg_en8137,
   output        cfg_en8138,
   output        cfg_en8139,
   output        cfg_en8140,
   output        cfg_en8141,
   output        cfg_en8142,
   output        cfg_en8143,
   output        cfg_en8144,
   output        cfg_en8145,
   output        cfg_en8146,
   output        cfg_en8147,
   output        cfg_en8148,
   output        cfg_en8149,
   output        cfg_en8150,
   output        cfg_en8151,
   output        cfg_en8152,
   output        cfg_en8153,
   output        cfg_en8154,
   output        cfg_en8155,
   output        cfg_en8156,
   output        cfg_en8157,
   output        cfg_en8158,
   output        cfg_en8159,
   output        cfg_en8160,
   output        cfg_en8161,
   output        cfg_en8162,
   output        cfg_en8163,
   output        cfg_en8164,
   output        cfg_en8165,
   output        cfg_en8166,
   output        cfg_en8167,
   output        cfg_en8168,
   output        cfg_en8169,
   output        cfg_en8170,
   output        cfg_en8171,
   output        cfg_en8172,
   output        cfg_en8173,
   output        cfg_en8174,
   output        cfg_en8175,
   output        cfg_en8176,
   output        cfg_en8177,
   output        cfg_en8178,
   output        cfg_en8179,
   output        cfg_en8180,
   output        cfg_en8181,
   output        cfg_en8182,
   output        cfg_en8183,
   output        cfg_en8184,
   output        cfg_en8185,
   output        cfg_en8186,
   output        cfg_en8187,
   output        cfg_en8188,
   output        cfg_en8189,
   output        cfg_en8190,
   output        cfg_en8191,
   output        tc_cfg_en,
   output        cc_cfg_en0,
   output        cc_cfg_en1,
   output        cc_cfg_en2,
   output        cc_cfg_en3,
   output        cfg_din0,
   output        cfg_din1,
   output        cfg_din2,
   output        cfg_din3,
   output        cfg_din4,
   output        cfg_din5,
   output        cfg_din6,
   output        cfg_din7,
   output        cfg_din8,
   output        cfg_din9,
   output        cfg_din10,
   output        cfg_din11,
   output        cfg_din12,
   output        cfg_din13,
   output        cfg_din14,
   output        cfg_din15,
   output        cfg_din16,
   output        cfg_din17,
   output        cfg_din18,
   output        cfg_din19,
   output        cfg_din20,
   output        cfg_din21,
   output        cfg_din22,
   output        cfg_din23,
   output        cfg_din24,
   output        cfg_din25,
   output        cfg_din26,
   output        cfg_din27,
   output        cfg_din28,
   output        cfg_din29,
   output        cfg_din30,
   output        cfg_din31,
   output        cfg_din32,
   output        cfg_din33,
   output        cfg_din34,
   output        cfg_din35,
   output        cfg_din36,
   output        cfg_din37,
   output        cfg_din38,
   output        cfg_din39,
   output        cfg_din40,
   output        cfg_din41,
   output        cfg_din42,
   output        cfg_din43,
   output        cfg_din44,
   output        cfg_din45,
   output        cfg_din46,
   output        cfg_din47,
   output        cfg_din48,
   output        cfg_din49,
   output        cfg_din50,
   output        cfg_din51,
   output        cfg_din52,
   output        cfg_din53,
   output        cfg_din54,
   output        cfg_din55,
   output        cfg_din56,
   output        cfg_din57,
   output        cfg_din58,
   output        cfg_din59,
   output        cfg_din60,
   output        cfg_din61,
   output        cfg_din62,
   output        cfg_din63,
   output        cfg_din64,
   output        cfg_din65,
   output        cfg_din66,
   output        cfg_din67,
   output        cfg_din68,
   output        cfg_din69,
   output        cfg_din70,
   output        cfg_din71,
   output        cfg_din72,
   output        cfg_din73,
   output        cfg_din74,
   output        cfg_din75,
   output        cfg_din76,
   output        cfg_din77,
   output        cfg_din78,
   output        cfg_din79,
   output        cfg_din80,
   output        cfg_din81,
   output        cfg_din82,
   output        cfg_din83,
   output        cfg_din84,
   output        cfg_din85,
   output        cfg_din86,
   output        cfg_din87,
   output        cfg_din88,
   output        cfg_din89,
   output        cfg_din90,
   output        cfg_din91,
   output        cfg_din92,
   output        cfg_din93,
   output        cfg_din94,
   output        cfg_din95,
   output        cfg_din96,
   output        cfg_din97,
   output        cfg_din98,
   output        cfg_din99,
   output        cfg_din100,
   output        cfg_din101,
   output        cfg_din102,
   output        cfg_din103,
   output        cfg_din104,
   output        cfg_din105,
   output        cfg_din106,
   output        cfg_din107,
   output        cfg_din108,
   output        cfg_din109,
   output        cfg_din110,
   output        cfg_din111,
   output        cfg_din112,
   output        cfg_din113,
   output        cfg_din114,
   output        cfg_din115,
   output        cfg_din116,
   output        cfg_din117,
   output        cfg_din118,
   output        cfg_din119,
   output        cfg_din120,
   output        cfg_din121,
   output        cfg_din122,
   output        cfg_din123,
   output        cfg_din124,
   output        cfg_din125,
   output        cfg_din126,
   output        cfg_din127,
   output        cfg_din128,
   output        cfg_din129,
   output        cfg_din130,
   output        cfg_din131,
   output        cfg_din132,
   output        cfg_din133,
   output        cfg_din134,
   output        cfg_din135,
   output        cfg_din136,
   output        cfg_din137,
   output        cfg_din138,
   output        cfg_din139,
   output        cfg_din140,
   output        cfg_din141,
   output        cfg_din142,
   output        cfg_din143,
   output        cfg_din144,
   output        cfg_din145,
   output        cfg_din146,
   output        cfg_din147,
   output        cfg_din148,
   output        cfg_din149,
   output        cfg_din150,
   output        cfg_din151,
   output        cfg_din152,
   output        cfg_din153,
   output        cfg_din154,
   output        cfg_din155,
   output        cfg_din156,
   output        cfg_din157,
   output        cfg_din158,
   output        cfg_din159,
   output        cfg_din160,
   output        cfg_din161,
   output        cfg_din162,
   output        cfg_din163,
   output        cfg_din164,
   output        cfg_din165,
   output        cfg_din166,
   output        cfg_din167,
   output        cfg_din168,
   output        cfg_din169,
   output        cfg_din170,
   output        cfg_din171,
   output        cfg_din172,
   output        cfg_din173,
   output        cfg_din174,
   output        cfg_din175,
   output        cfg_din176,
   output        cfg_din177,
   output        cfg_din178,
   output        cfg_din179,
   output        cfg_din180,
   output        cfg_din181,
   output        cfg_din182,
   output        cfg_din183,
   output        cfg_din184,
   output        cfg_din185,
   output        cfg_din186,
   output        cfg_din187,
   output        cfg_din188,
   output        cfg_din189,
   output        cfg_din190,
   output        cfg_din191,
   output        cfg_din192,
   output        cfg_din193,
   output        cfg_din194,
   output        cfg_din195,
   output        cfg_din196,
   output        cfg_din197,
   output        cfg_din198,
   output        cfg_din199,
   output        cfg_din200,
   output        cfg_din201,
   output        cfg_din202,
   output        cfg_din203,
   output        cfg_din204,
   output        cfg_din205,
   output        cfg_din206,
   output        cfg_din207,
   output        cfg_din208,
   output        cfg_din209,
   output        cfg_din210,
   output        cfg_din211,
   output        cfg_din212,
   output        cfg_din213,
   output        cfg_din214,
   output        cfg_din215,
   output        cfg_din216,
   output        cfg_din217,
   output        cfg_din218,
   output        cfg_din219,
   output        cfg_din220,
   output        cfg_din221,
   output        cfg_din222,
   output        cfg_din223,
   output        cfg_din224,
   output        cfg_din225,
   output        cfg_din226,
   output        cfg_din227,
   output        cfg_din228,
   output        cfg_din229,
   output        cfg_din230,
   output        cfg_din231,
   output        cfg_din232,
   output        cfg_din233,
   output        cfg_din234,
   output        cfg_din235,
   output        cfg_din236,
   output        cfg_din237,
   output        cfg_din238,
   output        cfg_din239,
   output        cfg_din240,
   output        cfg_din241,
   output        cfg_din242,
   output        cfg_din243,
   output        cfg_din244,
   output        cfg_din245,
   output        cfg_din246,
   output        cfg_din247,
   output        cfg_din248,
   output        cfg_din249,
   output        cfg_din250,
   output        cfg_din251,
   output        cfg_din252,
   output        cfg_din253,
   output        cfg_din254,
   output        cfg_din255,
   output        cfg_din256,
   output        cfg_din257,
   output        cfg_din258,
   output        cfg_din259,
   output        cfg_din260,
   output        cfg_din261,
   output        cfg_din262,
   output        cfg_din263,
   output        cfg_din264,
   output        cfg_din265,
   output        cfg_din266,
   output        cfg_din267,
   output        cfg_din268,
   output        cfg_din269,
   output        cfg_din270,
   output        cfg_din271,
   output        cfg_din272,
   output        cfg_din273,
   output        cfg_din274,
   output        cfg_din275,
   output        cfg_din276,
   output        cfg_din277,
   output        cfg_din278,
   output        cfg_din279,
   output        cfg_din280,
   output        cfg_din281,
   output        cfg_din282,
   output        cfg_din283,
   output        cfg_din284,
   output        cfg_din285,
   output        cfg_din286,
   output        cfg_din287,
   output        cfg_din288,
   output        cfg_din289,
   output        cfg_din290,
   output        cfg_din291,
   output        cfg_din292,
   output        cfg_din293,
   output        cfg_din294,
   output        cfg_din295,
   output        cfg_din296,
   output        cfg_din297,
   output        cfg_din298,
   output        cfg_din299,
   output        cfg_din300,
   output        cfg_din301,
   output        cfg_din302,
   output        cfg_din303,
   output        cfg_din304,
   output        cfg_din305,
   output        cfg_din306,
   output        cfg_din307,
   output        cfg_din308,
   output        cfg_din309,
   output        cfg_din310,
   output        cfg_din311,
   output        cfg_din312,
   output        cfg_din313,
   output        cfg_din314,
   output        cfg_din315,
   output        cfg_din316,
   output        cfg_din317,
   output        cfg_din318,
   output        cfg_din319,
   output        cfg_din320,
   output        cfg_din321,
   output        cfg_din322,
   output        cfg_din323,
   output        cfg_din324,
   output        cfg_din325,
   output        cfg_din326,
   output        cfg_din327,
   output        cfg_din328,
   output        cfg_din329,
   output        cfg_din330,
   output        cfg_din331,
   output        cfg_din332,
   output        cfg_din333,
   output        cfg_din334,
   output        cfg_din335,
   output        cfg_din336,
   output        cfg_din337,
   output        cfg_din338,
   output        cfg_din339,
   output        cfg_din340,
   output        cfg_din341,
   output        cfg_din342,
   output        cfg_din343,
   output        cfg_din344,
   output        cfg_din345,
   output        cfg_din346,
   output        cfg_din347,
   output        cfg_din348,
   output        cfg_din349,
   output        cfg_din350,
   output        cfg_din351,
   output        cfg_din352,
   output        cfg_din353,
   output        cfg_din354,
   output        cfg_din355,
   output        cfg_din356,
   output        cfg_din357,
   output        cfg_din358,
   output        cfg_din359,
   output        cfg_din360,
   output        cfg_din361,
   output        cfg_din362,
   output        cfg_din363,
   output        cfg_din364,
   output        cfg_din365,
   output        cfg_din366,
   output        cfg_din367,
   output        cfg_din368,
   output        cfg_din369,
   output        cfg_din370,
   output        cfg_din371,
   output        cfg_din372,
   output        cfg_din373,
   output        cfg_din374,
   output        cfg_din375,
   output        cfg_din376,
   output        cfg_din377,
   output        cfg_din378,
   output        cfg_din379,
   output        cfg_din380,
   output        cfg_din381,
   output        cfg_din382,
   output        cfg_din383,
   output        cfg_din384,
   output        cfg_din385,
   output        cfg_din386,
   output        cfg_din387,
   output        cfg_din388,
   output        cfg_din389,
   output        cfg_din390,
   output        cfg_din391,
   output        cfg_din392,
   output        cfg_din393,
   output        cfg_din394,
   output        cfg_din395,
   output        cfg_din396,
   output        cfg_din397,
   output        cfg_din398,
   output        cfg_din399,
   output        cfg_din400,
   output        cfg_din401,
   output        cfg_din402,
   output        cfg_din403,
   output        cfg_din404,
   output        cfg_din405,
   output        cfg_din406,
   output        cfg_din407,
   output        cfg_din408,
   output        cfg_din409,
   output        cfg_din410,
   output        cfg_din411,
   output        cfg_din412,
   output        cfg_din413,
   output        cfg_din414,
   output        cfg_din415,
   output        cfg_din416,
   output        cfg_din417,
   output        cfg_din418,
   output        cfg_din419,
   output        cfg_din420,
   output        cfg_din421,
   output        cfg_din422,
   output        cfg_din423,
   output        cfg_din424,
   output        cfg_din425,
   output        cfg_din426,
   output        cfg_din427,
   output        cfg_din428,
   output        cfg_din429,
   output        cfg_din430,
   output        cfg_din431,
   output        cfg_din432,
   output        cfg_din433,
   output        cfg_din434,
   output        cfg_din435,
   output        cfg_din436,
   output        cfg_din437,
   output        cfg_din438,
   output        cfg_din439,
   output        cfg_din440,
   output        cfg_din441,
   output        cfg_din442,
   output        cfg_din443,
   output        cfg_din444,
   output        cfg_din445,
   output        cfg_din446,
   output        cfg_din447,
   output        cfg_din448,
   output        cfg_din449,
   output        cfg_din450,
   output        cfg_din451,
   output        cfg_din452,
   output        cfg_din453,
   output        cfg_din454,
   output        cfg_din455,
   output        cfg_din456,
   output        cfg_din457,
   output        cfg_din458,
   output        cfg_din459,
   output        cfg_din460,
   output        cfg_din461,
   output        cfg_din462,
   output        cfg_din463,
   output        cfg_din464,
   output        cfg_din465,
   output        cfg_din466,
   output        cfg_din467,
   output        cfg_din468,
   output        cfg_din469,
   output        cfg_din470,
   output        cfg_din471,
   output        cfg_din472,
   output        cfg_din473,
   output        cfg_din474,
   output        cfg_din475,
   output        cfg_din476,
   output        cfg_din477,
   output        cfg_din478,
   output        cfg_din479,
   output        cfg_din480,
   output        cfg_din481,
   output        cfg_din482,
   output        cfg_din483,
   output        cfg_din484,
   output        cfg_din485,
   output        cfg_din486,
   output        cfg_din487,
   output        cfg_din488,
   output        cfg_din489,
   output        cfg_din490,
   output        cfg_din491,
   output        cfg_din492,
   output        cfg_din493,
   output        cfg_din494,
   output        cfg_din495,
   output        cfg_din496,
   output        cfg_din497,
   output        cfg_din498,
   output        cfg_din499,
   output        cfg_din500,
   output        cfg_din501,
   output        cfg_din502,
   output        cfg_din503,
   output        cfg_din504,
   output        cfg_din505,
   output        cfg_din506,
   output        cfg_din507,
   output        cfg_din508,
   output        cfg_din509,
   output        cfg_din510,
   output        cfg_din511,
   output        cfg_din512,
   output        cfg_din513,
   output        cfg_din514,
   output        cfg_din515,
   output        cfg_din516,
   output        cfg_din517,
   output        cfg_din518,
   output        cfg_din519,
   output        cfg_din520,
   output        cfg_din521,
   output        cfg_din522,
   output        cfg_din523,
   output        cfg_din524,
   output        cfg_din525,
   output        cfg_din526,
   output        cfg_din527,
   output        cfg_din528,
   output        cfg_din529,
   output        cfg_din530,
   output        cfg_din531,
   output        cfg_din532,
   output        cfg_din533,
   output        cfg_din534,
   output        cfg_din535,
   output        cfg_din536,
   output        cfg_din537,
   output        cfg_din538,
   output        cfg_din539,
   output        cfg_din540,
   output        cfg_din541,
   output        cfg_din542,
   output        cfg_din543,
   output        cfg_din544,
   output        cfg_din545,
   output        cfg_din546,
   output        cfg_din547,
   output        cfg_din548,
   output        cfg_din549,
   output        cfg_din550,
   output        cfg_din551,
   output        cfg_din552,
   output        cfg_din553,
   output        cfg_din554,
   output        cfg_din555,
   output        cfg_din556,
   output        cfg_din557,
   output        cfg_din558,
   output        cfg_din559,
   output        cfg_din560,
   output        cfg_din561,
   output        cfg_din562,
   output        cfg_din563,
   output        cfg_din564,
   output        cfg_din565,
   output        cfg_din566,
   output        cfg_din567,
   output        cfg_din568,
   output        cfg_din569,
   output        cfg_din570,
   output        cfg_din571,
   output        cfg_din572,
   output        cfg_din573,
   output        cfg_din574,
   output        cfg_din575,
   output        cfg_din576,
   output        cfg_din577,
   output        cfg_din578,
   output        cfg_din579,
   output        cfg_din580,
   output        cfg_din581,
   output        cfg_din582,
   output        cfg_din583,
   output        cfg_din584,
   output        cfg_din585,
   output        cfg_din586,
   output        cfg_din587,
   output        cfg_din588,
   output        cfg_din589,
   output        cfg_din590,
   output        cfg_din591,
   output        cfg_din592,
   output        cfg_din593,
   output        cfg_din594,
   output        cfg_din595,
   output        cfg_din596,
   output        cfg_din597,
   output        cfg_din598,
   output        cfg_din599,
   output        cfg_din600,
   output        cfg_din601,
   output        cfg_din602,
   output        cfg_din603,
   output        cfg_din604,
   output        cfg_din605,
   output        cfg_din606,
   output        cfg_din607,
   output        cfg_din608,
   output        cfg_din609,
   output        cfg_din610,
   output        cfg_din611,
   output        cfg_din612,
   output        cfg_din613,
   output        cfg_din614,
   output        cfg_din615,
   output        cfg_din616,
   output        cfg_din617,
   output        cfg_din618,
   output        cfg_din619,
   output        cfg_din620,
   output        cfg_din621,
   output        cfg_din622,
   output        cfg_din623,
   output        cfg_din624,
   output        cfg_din625,
   output        cfg_din626,
   output        cfg_din627,
   output        cfg_din628,
   output        cfg_din629,
   output        cfg_din630,
   output        cfg_din631,
   output        cfg_din632,
   output        cfg_din633,
   output        cfg_din634,
   output        cfg_din635,
   output        cfg_din636,
   output        cfg_din637,
   output        cfg_din638,
   output        cfg_din639,
   output        cfg_din640,
   output        cfg_din641,
   output        cfg_din642,
   output        cfg_din643,
   output        cfg_din644,
   output        cfg_din645,
   output        cfg_din646,
   output        cfg_din647,
   output        cfg_din648,
   output        cfg_din649,
   output        cfg_din650,
   output        cfg_din651,
   output        cfg_din652,
   output        cfg_din653,
   output        cfg_din654,
   output        cfg_din655,
   output        cfg_din656,
   output        cfg_din657,
   output        cfg_din658,
   output        cfg_din659,
   output        cfg_din660,
   output        cfg_din661,
   output        cfg_din662,
   output        cfg_din663,
   output        cfg_din664,
   output        cfg_din665,
   output        cfg_din666,
   output        cfg_din667,
   output        cfg_din668,
   output        cfg_din669,
   output        cfg_din670,
   output        cfg_din671,
   output        cfg_din672,
   output        cfg_din673,
   output        cfg_din674,
   output        cfg_din675,
   output        cfg_din676,
   output        cfg_din677,
   output        cfg_din678,
   output        cfg_din679,
   output        cfg_din680,
   output        cfg_din681,
   output        cfg_din682,
   output        cfg_din683,
   output        cfg_din684,
   output        cfg_din685,
   output        cfg_din686,
   output        cfg_din687,
   output        cfg_din688,
   output        cfg_din689,
   output        cfg_din690,
   output        cfg_din691,
   output        cfg_din692,
   output        cfg_din693,
   output        cfg_din694,
   output        cfg_din695,
   output        cfg_din696,
   output        cfg_din697,
   output        cfg_din698,
   output        cfg_din699,
   output        cfg_din700,
   output        cfg_din701,
   output        cfg_din702,
   output        cfg_din703,
   output        cfg_din704,
   output        cfg_din705,
   output        cfg_din706,
   output        cfg_din707,
   output        cfg_din708,
   output        cfg_din709,
   output        cfg_din710,
   output        cfg_din711,
   output        cfg_din712,
   output        cfg_din713,
   output        cfg_din714,
   output        cfg_din715,
   output        cfg_din716,
   output        cfg_din717,
   output        cfg_din718,
   output        cfg_din719,
   output        cfg_din720,
   output        cfg_din721,
   output        cfg_din722,
   output        cfg_din723,
   output        cfg_din724,
   output        cfg_din725,
   output        cfg_din726,
   output        cfg_din727,
   output        cfg_din728,
   output        cfg_din729,
   output        cfg_din730,
   output        cfg_din731,
   output        cfg_din732,
   output        cfg_din733,
   output        cfg_din734,
   output        cfg_din735,
   output        cfg_din736,
   output        cfg_din737,
   output        cfg_din738,
   output        cfg_din739,
   output        cfg_din740,
   output        cfg_din741,
   output        cfg_din742,
   output        cfg_din743,
   output        cfg_din744,
   output        cfg_din745,
   output        cfg_din746,
   output        cfg_din747,
   output        cfg_din748,
   output        cfg_din749,
   output        cfg_din750,
   output        cfg_din751,
   output        cfg_din752,
   output        cfg_din753,
   output        cfg_din754,
   output        cfg_din755,
   output        cfg_din756,
   output        cfg_din757,
   output        cfg_din758,
   output        cfg_din759,
   output        cfg_din760,
   output        cfg_din761,
   output        cfg_din762,
   output        cfg_din763,
   output        cfg_din764,
   output        cfg_din765,
   output        cfg_din766,
   output        cfg_din767,
   output        cfg_din768,
   output        cfg_din769,
   output        cfg_din770,
   output        cfg_din771,
   output        cfg_din772,
   output        cfg_din773,
   output        cfg_din774,
   output        cfg_din775,
   output        cfg_din776,
   output        cfg_din777,
   output        cfg_din778,
   output        cfg_din779,
   output        cfg_din780,
   output        cfg_din781,
   output        cfg_din782,
   output        cfg_din783,
   output        cfg_din784,
   output        cfg_din785,
   output        cfg_din786,
   output        cfg_din787,
   output        cfg_din788,
   output        cfg_din789,
   output        cfg_din790,
   output        cfg_din791,
   output        cfg_din792,
   output        cfg_din793,
   output        cfg_din794,
   output        cfg_din795,
   output        cfg_din796,
   output        cfg_din797,
   output        cfg_din798,
   output        cfg_din799,
   output        cfg_din800,
   output        cfg_din801,
   output        cfg_din802,
   output        cfg_din803,
   output        cfg_din804,
   output        cfg_din805,
   output        cfg_din806,
   output        cfg_din807,
   output        cfg_din808,
   output        cfg_din809,
   output        cfg_din810,
   output        cfg_din811,
   output        cfg_din812,
   output        cfg_din813,
   output        cfg_din814,
   output        cfg_din815,
   output        cfg_din816,
   output        cfg_din817,
   output        cfg_din818,
   output        cfg_din819,
   output        cfg_din820,
   output        cfg_din821,
   output        cfg_din822,
   output        cfg_din823,
   output        cfg_din824,
   output        cfg_din825,
   output        cfg_din826,
   output        cfg_din827,
   output        cfg_din828,
   output        cfg_din829,
   output        cfg_din830,
   output        cfg_din831,
   output        cfg_din832,
   output        cfg_din833,
   output        cfg_din834,
   output        cfg_din835,
   output        cfg_din836,
   output        cfg_din837,
   output        cfg_din838,
   output        cfg_din839,
   output        cfg_din840,
   output        cfg_din841,
   output        cfg_din842,
   output        cfg_din843,
   output        cfg_din844,
   output        cfg_din845,
   output        cfg_din846,
   output        cfg_din847,
   output        cfg_din848,
   output        cfg_din849,
   output        cfg_din850,
   output        cfg_din851,
   output        cfg_din852,
   output        cfg_din853,
   output        cfg_din854,
   output        cfg_din855,
   output        cfg_din856,
   output        cfg_din857,
   output        cfg_din858,
   output        cfg_din859,
   output        cfg_din860,
   output        cfg_din861,
   output        cfg_din862,
   output        cfg_din863,
   output        cfg_din864,
   output        cfg_din865,
   output        cfg_din866,
   output        cfg_din867,
   output        cfg_din868,
   output        cfg_din869,
   output        cfg_din870,
   output        cfg_din871,
   output        cfg_din872,
   output        cfg_din873,
   output        cfg_din874,
   output        cfg_din875,
   output        cfg_din876,
   output        cfg_din877,
   output        cfg_din878,
   output        cfg_din879,
   output        cfg_din880,
   output        cfg_din881,
   output        cfg_din882,
   output        cfg_din883,
   output        cfg_din884,
   output        cfg_din885,
   output        cfg_din886,
   output        cfg_din887,
   output        cfg_din888,
   output        cfg_din889,
   output        cfg_din890,
   output        cfg_din891,
   output        cfg_din892,
   output        cfg_din893,
   output        cfg_din894,
   output        cfg_din895,
   output        cfg_din896,
   output        cfg_din897,
   output        cfg_din898,
   output        cfg_din899,
   output        cfg_din900,
   output        cfg_din901,
   output        cfg_din902,
   output        cfg_din903,
   output        cfg_din904,
   output        cfg_din905,
   output        cfg_din906,
   output        cfg_din907,
   output        cfg_din908,
   output        cfg_din909,
   output        cfg_din910,
   output        cfg_din911,
   output        cfg_din912,
   output        cfg_din913,
   output        cfg_din914,
   output        cfg_din915,
   output        cfg_din916,
   output        cfg_din917,
   output        cfg_din918,
   output        cfg_din919,
   output        cfg_din920,
   output        cfg_din921,
   output        cfg_din922,
   output        cfg_din923,
   output        cfg_din924,
   output        cfg_din925,
   output        cfg_din926,
   output        cfg_din927,
   output        cfg_din928,
   output        cfg_din929,
   output        cfg_din930,
   output        cfg_din931,
   output        cfg_din932,
   output        cfg_din933,
   output        cfg_din934,
   output        cfg_din935,
   output        cfg_din936,
   output        cfg_din937,
   output        cfg_din938,
   output        cfg_din939,
   output        cfg_din940,
   output        cfg_din941,
   output        cfg_din942,
   output        cfg_din943,
   output        cfg_din944,
   output        cfg_din945,
   output        cfg_din946,
   output        cfg_din947,
   output        cfg_din948,
   output        cfg_din949,
   output        cfg_din950,
   output        cfg_din951,
   output        cfg_din952,
   output        cfg_din953,
   output        cfg_din954,
   output        cfg_din955,
   output        cfg_din956,
   output        cfg_din957,
   output        cfg_din958,
   output        cfg_din959,
   output        cfg_din960,
   output        cfg_din961,
   output        cfg_din962,
   output        cfg_din963,
   output        cfg_din964,
   output        cfg_din965,
   output        cfg_din966,
   output        cfg_din967,
   output        cfg_din968,
   output        cfg_din969,
   output        cfg_din970,
   output        cfg_din971,
   output        cfg_din972,
   output        cfg_din973,
   output        cfg_din974,
   output        cfg_din975,
   output        cfg_din976,
   output        cfg_din977,
   output        cfg_din978,
   output        cfg_din979,
   output        cfg_din980,
   output        cfg_din981,
   output        cfg_din982,
   output        cfg_din983,
   output        cfg_din984,
   output        cfg_din985,
   output        cfg_din986,
   output        cfg_din987,
   output        cfg_din988,
   output        cfg_din989,
   output        cfg_din990,
   output        cfg_din991,
   output        cfg_din992,
   output        cfg_din993,
   output        cfg_din994,
   output        cfg_din995,
   output        cfg_din996,
   output        cfg_din997,
   output        cfg_din998,
   output        cfg_din999,
   output        cfg_din1000,
   output        cfg_din1001,
   output        cfg_din1002,
   output        cfg_din1003,
   output        cfg_din1004,
   output        cfg_din1005,
   output        cfg_din1006,
   output        cfg_din1007,
   output        cfg_din1008,
   output        cfg_din1009,
   output        cfg_din1010,
   output        cfg_din1011,
   output        cfg_din1012,
   output        cfg_din1013,
   output        cfg_din1014,
   output        cfg_din1015,
   output        cfg_din1016,
   output        cfg_din1017,
   output        cfg_din1018,
   output        cfg_din1019,
   output        cfg_din1020,
   output        cfg_din1021,
   output        cfg_din1022,
   output        cfg_din1023,
   output        cfg_din1024,
   output        cfg_din1025,
   output        cfg_din1026,
   output        cfg_din1027,
   output        cfg_din1028,
   output        cfg_din1029,
   output        cfg_din1030,
   output        cfg_din1031,
   output        cfg_din1032,
   output        cfg_din1033,
   output        cfg_din1034,
   output        cfg_din1035,
   output        cfg_din1036,
   output        cfg_din1037,
   output        cfg_din1038,
   output        cfg_din1039,
   output        cfg_din1040,
   output        cfg_din1041,
   output        cfg_din1042,
   output        cfg_din1043,
   output        cfg_din1044,
   output        cfg_din1045,
   output        cfg_din1046,
   output        cfg_din1047,
   output        cfg_din1048,
   output        cfg_din1049,
   output        cfg_din1050,
   output        cfg_din1051,
   output        cfg_din1052,
   output        cfg_din1053,
   output        cfg_din1054,
   output        cfg_din1055,
   output        cfg_din1056,
   output        cfg_din1057,
   output        cfg_din1058,
   output        cfg_din1059,
   output        cfg_din1060,
   output        cfg_din1061,
   output        cfg_din1062,
   output        cfg_din1063,
   output        cfg_din1064,
   output        cfg_din1065,
   output        cfg_din1066,
   output        cfg_din1067,
   output        cfg_din1068,
   output        cfg_din1069,
   output        cfg_din1070,
   output        cfg_din1071,
   output        cfg_din1072,
   output        cfg_din1073,
   output        cfg_din1074,
   output        cfg_din1075,
   output        cfg_din1076,
   output        cfg_din1077,
   output        cfg_din1078,
   output        cfg_din1079,
   output        cfg_din1080,
   output        cfg_din1081,
   output        cfg_din1082,
   output        cfg_din1083,
   output        cfg_din1084,
   output        cfg_din1085,
   output        cfg_din1086,
   output        cfg_din1087,
   output        cfg_din1088,
   output        cfg_din1089,
   output        cfg_din1090,
   output        cfg_din1091,
   output        cfg_din1092,
   output        cfg_din1093,
   output        cfg_din1094,
   output        cfg_din1095,
   output        cfg_din1096,
   output        cfg_din1097,
   output        cfg_din1098,
   output        cfg_din1099,
   output        cfg_din1100,
   output        cfg_din1101,
   output        cfg_din1102,
   output        cfg_din1103,
   output        cfg_din1104,
   output        cfg_din1105,
   output        cfg_din1106,
   output        cfg_din1107,
   output        cfg_din1108,
   output        cfg_din1109,
   output        cfg_din1110,
   output        cfg_din1111,
   output        cfg_din1112,
   output        cfg_din1113,
   output        cfg_din1114,
   output        cfg_din1115,
   output        cfg_din1116,
   output        cfg_din1117,
   output        cfg_din1118,
   output        cfg_din1119,
   output        cfg_din1120,
   output        cfg_din1121,
   output        cfg_din1122,
   output        cfg_din1123,
   output        cfg_din1124,
   output        cfg_din1125,
   output        cfg_din1126,
   output        cfg_din1127,
   output        cfg_din1128,
   output        cfg_din1129,
   output        cfg_din1130,
   output        cfg_din1131,
   output        cfg_din1132,
   output        cfg_din1133,
   output        cfg_din1134,
   output        cfg_din1135,
   output        cfg_din1136,
   output        cfg_din1137,
   output        cfg_din1138,
   output        cfg_din1139,
   output        cfg_din1140,
   output        cfg_din1141,
   output        cfg_din1142,
   output        cfg_din1143,
   output        cfg_din1144,
   output        cfg_din1145,
   output        cfg_din1146,
   output        cfg_din1147,
   output        cfg_din1148,
   output        cfg_din1149,
   output        cfg_din1150,
   output        cfg_din1151,
   output        cfg_din1152,
   output        cfg_din1153,
   output        cfg_din1154,
   output        cfg_din1155,
   output        cfg_din1156,
   output        cfg_din1157,
   output        cfg_din1158,
   output        cfg_din1159,
   output        cfg_din1160,
   output        cfg_din1161,
   output        cfg_din1162,
   output        cfg_din1163,
   output        cfg_din1164,
   output        cfg_din1165,
   output        cfg_din1166,
   output        cfg_din1167,
   output        cfg_din1168,
   output        cfg_din1169,
   output        cfg_din1170,
   output        cfg_din1171,
   output        cfg_din1172,
   output        cfg_din1173,
   output        cfg_din1174,
   output        cfg_din1175,
   output        cfg_din1176,
   output        cfg_din1177,
   output        cfg_din1178,
   output        cfg_din1179,
   output        cfg_din1180,
   output        cfg_din1181,
   output        cfg_din1182,
   output        cfg_din1183,
   output        cfg_din1184,
   output        cfg_din1185,
   output        cfg_din1186,
   output        cfg_din1187,
   output        cfg_din1188,
   output        cfg_din1189,
   output        cfg_din1190,
   output        cfg_din1191,
   output        cfg_din1192,
   output        cfg_din1193,
   output        cfg_din1194,
   output        cfg_din1195,
   output        cfg_din1196,
   output        cfg_din1197,
   output        cfg_din1198,
   output        cfg_din1199,
   output        cfg_din1200,
   output        cfg_din1201,
   output        cfg_din1202,
   output        cfg_din1203,
   output        cfg_din1204,
   output        cfg_din1205,
   output        cfg_din1206,
   output        cfg_din1207,
   output        cfg_din1208,
   output        cfg_din1209,
   output        cfg_din1210,
   output        cfg_din1211,
   output        cfg_din1212,
   output        cfg_din1213,
   output        cfg_din1214,
   output        cfg_din1215,
   output        cfg_din1216,
   output        cfg_din1217,
   output        cfg_din1218,
   output        cfg_din1219,
   output        cfg_din1220,
   output        cfg_din1221,
   output        cfg_din1222,
   output        cfg_din1223,
   output        cfg_din1224,
   output        cfg_din1225,
   output        cfg_din1226,
   output        cfg_din1227,
   output        cfg_din1228,
   output        cfg_din1229,
   output        cfg_din1230,
   output        cfg_din1231,
   output        cfg_din1232,
   output        cfg_din1233,
   output        cfg_din1234,
   output        cfg_din1235,
   output        cfg_din1236,
   output        cfg_din1237,
   output        cfg_din1238,
   output        cfg_din1239,
   output        cfg_din1240,
   output        cfg_din1241,
   output        cfg_din1242,
   output        cfg_din1243,
   output        cfg_din1244,
   output        cfg_din1245,
   output        cfg_din1246,
   output        cfg_din1247,
   output        cfg_din1248,
   output        cfg_din1249,
   output        cfg_din1250,
   output        cfg_din1251,
   output        cfg_din1252,
   output        cfg_din1253,
   output        cfg_din1254,
   output        cfg_din1255,
   output        cfg_din1256,
   output        cfg_din1257,
   output        cfg_din1258,
   output        cfg_din1259,
   output        cfg_din1260,
   output        cfg_din1261,
   output        cfg_din1262,
   output        cfg_din1263,
   output        cfg_din1264,
   output        cfg_din1265,
   output        cfg_din1266,
   output        cfg_din1267,
   output        cfg_din1268,
   output        cfg_din1269,
   output        cfg_din1270,
   output        cfg_din1271,
   output        cfg_din1272,
   output        cfg_din1273,
   output        cfg_din1274,
   output        cfg_din1275,
   output        cfg_din1276,
   output        cfg_din1277,
   output        cfg_din1278,
   output        cfg_din1279,
   output        cfg_din1280,
   output        cfg_din1281,
   output        cfg_din1282,
   output        cfg_din1283,
   output        cfg_din1284,
   output        cfg_din1285,
   output        cfg_din1286,
   output        cfg_din1287,
   output        cfg_din1288,
   output        cfg_din1289,
   output        cfg_din1290,
   output        cfg_din1291,
   output        cfg_din1292,
   output        cfg_din1293,
   output        cfg_din1294,
   output        cfg_din1295,
   output        cfg_din1296,
   output        cfg_din1297,
   output        cfg_din1298,
   output        cfg_din1299,
   output        cfg_din1300,
   output        cfg_din1301,
   output        cfg_din1302,
   output        cfg_din1303,
   output        cfg_din1304,
   output        cfg_din1305,
   output        cfg_din1306,
   output        cfg_din1307,
   output        cfg_din1308,
   output        cfg_din1309,
   output        cfg_din1310,
   output        cfg_din1311,
   output        cfg_din1312,
   output        cfg_din1313,
   output        cfg_din1314,
   output        cfg_din1315,
   output        cfg_din1316,
   output        cfg_din1317,
   output        cfg_din1318,
   output        cfg_din1319,
   output        cfg_din1320,
   output        cfg_din1321,
   output        cfg_din1322,
   output        cfg_din1323,
   output        cfg_din1324,
   output        cfg_din1325,
   output        cfg_din1326,
   output        cfg_din1327,
   output        cfg_din1328,
   output        cfg_din1329,
   output        cfg_din1330,
   output        cfg_din1331,
   output        cfg_din1332,
   output        cfg_din1333,
   output        cfg_din1334,
   output        cfg_din1335,
   output        cfg_din1336,
   output        cfg_din1337,
   output        cfg_din1338,
   output        cfg_din1339,
   output        cfg_din1340,
   output        cfg_din1341,
   output        cfg_din1342,
   output        cfg_din1343,
   output        cfg_din1344,
   output        cfg_din1345,
   output        cfg_din1346,
   output        cfg_din1347,
   output        cfg_din1348,
   output        cfg_din1349,
   output        cfg_din1350,
   output        cfg_din1351,
   output        cfg_din1352,
   output        cfg_din1353,
   output        cfg_din1354,
   output        cfg_din1355,
   output        cfg_din1356,
   output        cfg_din1357,
   output        cfg_din1358,
   output        cfg_din1359,
   output        cfg_din1360,
   output        cfg_din1361,
   output        cfg_din1362,
   output        cfg_din1363,
   output        cfg_din1364,
   output        cfg_din1365,
   output        cfg_din1366,
   output        cfg_din1367,
   output        cfg_din1368,
   output        cfg_din1369,
   output        cfg_din1370,
   output        cfg_din1371,
   output        cfg_din1372,
   output        cfg_din1373,
   output        cfg_din1374,
   output        cfg_din1375,
   output        cfg_din1376,
   output        cfg_din1377,
   output        cfg_din1378,
   output        cfg_din1379,
   output        cfg_din1380,
   output        cfg_din1381,
   output        cfg_din1382,
   output        cfg_din1383,
   output        cfg_din1384,
   output        cfg_din1385,
   output        cfg_din1386,
   output        cfg_din1387,
   output        cfg_din1388,
   output        cfg_din1389,
   output        cfg_din1390,
   output        cfg_din1391,
   output        cfg_din1392,
   output        cfg_din1393,
   output        cfg_din1394,
   output        cfg_din1395,
   output        cfg_din1396,
   output        cfg_din1397,
   output        cfg_din1398,
   output        cfg_din1399,
   output        cfg_din1400,
   output        cfg_din1401,
   output        cfg_din1402,
   output        cfg_din1403,
   output        cfg_din1404,
   output        cfg_din1405,
   output        cfg_din1406,
   output        cfg_din1407,
   output        cfg_din1408,
   output        cfg_din1409,
   output        cfg_din1410,
   output        cfg_din1411,
   output        cfg_din1412,
   output        cfg_din1413,
   output        cfg_din1414,
   output        cfg_din1415,
   output        cfg_din1416,
   output        cfg_din1417,
   output        cfg_din1418,
   output        cfg_din1419,
   output        cfg_din1420,
   output        cfg_din1421,
   output        cfg_din1422,
   output        cfg_din1423,
   output        cfg_din1424,
   output        cfg_din1425,
   output        cfg_din1426,
   output        cfg_din1427,
   output        cfg_din1428,
   output        cfg_din1429,
   output        cfg_din1430,
   output        cfg_din1431,
   output        cfg_din1432,
   output        cfg_din1433,
   output        cfg_din1434,
   output        cfg_din1435,
   output        cfg_din1436,
   output        cfg_din1437,
   output        cfg_din1438,
   output        cfg_din1439,
   output        cfg_din1440,
   output        cfg_din1441,
   output        cfg_din1442,
   output        cfg_din1443,
   output        cfg_din1444,
   output        cfg_din1445,
   output        cfg_din1446,
   output        cfg_din1447,
   output        cfg_din1448,
   output        cfg_din1449,
   output        cfg_din1450,
   output        cfg_din1451,
   output        cfg_din1452,
   output        cfg_din1453,
   output        cfg_din1454,
   output        cfg_din1455,
   output        cfg_din1456,
   output        cfg_din1457,
   output        cfg_din1458,
   output        cfg_din1459,
   output        cfg_din1460,
   output        cfg_din1461,
   output        cfg_din1462,
   output        cfg_din1463,
   output        cfg_din1464,
   output        cfg_din1465,
   output        cfg_din1466,
   output        cfg_din1467,
   output        cfg_din1468,
   output        cfg_din1469,
   output        cfg_din1470,
   output        cfg_din1471,
   output        cfg_din1472,
   output        cfg_din1473,
   output        cfg_din1474,
   output        cfg_din1475,
   output        cfg_din1476,
   output        cfg_din1477,
   output        cfg_din1478,
   output        cfg_din1479,
   output        cfg_din1480,
   output        cfg_din1481,
   output        cfg_din1482,
   output        cfg_din1483,
   output        cfg_din1484,
   output        cfg_din1485,
   output        cfg_din1486,
   output        cfg_din1487,
   output        cfg_din1488,
   output        cfg_din1489,
   output        cfg_din1490,
   output        cfg_din1491,
   output        cfg_din1492,
   output        cfg_din1493,
   output        cfg_din1494,
   output        cfg_din1495,
   output        cfg_din1496,
   output        cfg_din1497,
   output        cfg_din1498,
   output        cfg_din1499,
   output        cfg_din1500,
   output        cfg_din1501,
   output        cfg_din1502,
   output        cfg_din1503,
   output        cfg_din1504,
   output        cfg_din1505,
   output        cfg_din1506,
   output        cfg_din1507,
   output        cfg_din1508,
   output        cfg_din1509,
   output        cfg_din1510,
   output        cfg_din1511,
   output        cfg_din1512,
   output        cfg_din1513,
   output        cfg_din1514,
   output        cfg_din1515,
   output        cfg_din1516,
   output        cfg_din1517,
   output        cfg_din1518,
   output        cfg_din1519,
   output        cfg_din1520,
   output        cfg_din1521,
   output        cfg_din1522,
   output        cfg_din1523,
   output        cfg_din1524,
   output        cfg_din1525,
   output        cfg_din1526,
   output        cfg_din1527,
   output        cfg_din1528,
   output        cfg_din1529,
   output        cfg_din1530,
   output        cfg_din1531,
   output        cfg_din1532,
   output        cfg_din1533,
   output        cfg_din1534,
   output        cfg_din1535,
   output        cfg_din1536,
   output        cfg_din1537,
   output        cfg_din1538,
   output        cfg_din1539,
   output        cfg_din1540,
   output        cfg_din1541,
   output        cfg_din1542,
   output        cfg_din1543,
   output        cfg_din1544,
   output        cfg_din1545,
   output        cfg_din1546,
   output        cfg_din1547,
   output        cfg_din1548,
   output        cfg_din1549,
   output        cfg_din1550,
   output        cfg_din1551,
   output        cfg_din1552,
   output        cfg_din1553,
   output        cfg_din1554,
   output        cfg_din1555,
   output        cfg_din1556,
   output        cfg_din1557,
   output        cfg_din1558,
   output        cfg_din1559,
   output        cfg_din1560,
   output        cfg_din1561,
   output        cfg_din1562,
   output        cfg_din1563,
   output        cfg_din1564,
   output        cfg_din1565,
   output        cfg_din1566,
   output        cfg_din1567,
   output        cfg_din1568,
   output        cfg_din1569,
   output        cfg_din1570,
   output        cfg_din1571,
   output        cfg_din1572,
   output        cfg_din1573,
   output        cfg_din1574,
   output        cfg_din1575,
   output        cfg_din1576,
   output        cfg_din1577,
   output        cfg_din1578,
   output        cfg_din1579,
   output        cfg_din1580,
   output        cfg_din1581,
   output        cfg_din1582,
   output        cfg_din1583,
   output        cfg_din1584,
   output        cfg_din1585,
   output        cfg_din1586,
   output        cfg_din1587,
   output        cfg_din1588,
   output        cfg_din1589,
   output        cfg_din1590,
   output        cfg_din1591,
   output        cfg_din1592,
   output        cfg_din1593,
   output        cfg_din1594,
   output        cfg_din1595,
   output        cfg_din1596,
   output        cfg_din1597,
   output        cfg_din1598,
   output        cfg_din1599,
   output        cfg_din1600,
   output        cfg_din1601,
   output        cfg_din1602,
   output        cfg_din1603,
   output        cfg_din1604,
   output        cfg_din1605,
   output        cfg_din1606,
   output        cfg_din1607,
   output        cfg_din1608,
   output        cfg_din1609,
   output        cfg_din1610,
   output        cfg_din1611,
   output        cfg_din1612,
   output        cfg_din1613,
   output        cfg_din1614,
   output        cfg_din1615,
   output        cfg_din1616,
   output        cfg_din1617,
   output        cfg_din1618,
   output        cfg_din1619,
   output        cfg_din1620,
   output        cfg_din1621,
   output        cfg_din1622,
   output        cfg_din1623,
   output        cfg_din1624,
   output        cfg_din1625,
   output        cfg_din1626,
   output        cfg_din1627,
   output        cfg_din1628,
   output        cfg_din1629,
   output        cfg_din1630,
   output        cfg_din1631,
   output        cfg_din1632,
   output        cfg_din1633,
   output        cfg_din1634,
   output        cfg_din1635,
   output        cfg_din1636,
   output        cfg_din1637,
   output        cfg_din1638,
   output        cfg_din1639,
   output        cfg_din1640,
   output        cfg_din1641,
   output        cfg_din1642,
   output        cfg_din1643,
   output        cfg_din1644,
   output        cfg_din1645,
   output        cfg_din1646,
   output        cfg_din1647,
   output        cfg_din1648,
   output        cfg_din1649,
   output        cfg_din1650,
   output        cfg_din1651,
   output        cfg_din1652,
   output        cfg_din1653,
   output        cfg_din1654,
   output        cfg_din1655,
   output        cfg_din1656,
   output        cfg_din1657,
   output        cfg_din1658,
   output        cfg_din1659,
   output        cfg_din1660,
   output        cfg_din1661,
   output        cfg_din1662,
   output        cfg_din1663,
   output        cfg_din1664,
   output        cfg_din1665,
   output        cfg_din1666,
   output        cfg_din1667,
   output        cfg_din1668,
   output        cfg_din1669,
   output        cfg_din1670,
   output        cfg_din1671,
   output        cfg_din1672,
   output        cfg_din1673,
   output        cfg_din1674,
   output        cfg_din1675,
   output        cfg_din1676,
   output        cfg_din1677,
   output        cfg_din1678,
   output        cfg_din1679,
   output        cfg_din1680,
   output        cfg_din1681,
   output        cfg_din1682,
   output        cfg_din1683,
   output        cfg_din1684,
   output        cfg_din1685,
   output        cfg_din1686,
   output        cfg_din1687,
   output        cfg_din1688,
   output        cfg_din1689,
   output        cfg_din1690,
   output        cfg_din1691,
   output        cfg_din1692,
   output        cfg_din1693,
   output        cfg_din1694,
   output        cfg_din1695,
   output        cfg_din1696,
   output        cfg_din1697,
   output        cfg_din1698,
   output        cfg_din1699,
   output        cfg_din1700,
   output        cfg_din1701,
   output        cfg_din1702,
   output        cfg_din1703,
   output        cfg_din1704,
   output        cfg_din1705,
   output        cfg_din1706,
   output        cfg_din1707,
   output        cfg_din1708,
   output        cfg_din1709,
   output        cfg_din1710,
   output        cfg_din1711,
   output        cfg_din1712,
   output        cfg_din1713,
   output        cfg_din1714,
   output        cfg_din1715,
   output        cfg_din1716,
   output        cfg_din1717,
   output        cfg_din1718,
   output        cfg_din1719,
   output        cfg_din1720,
   output        cfg_din1721,
   output        cfg_din1722,
   output        cfg_din1723,
   output        cfg_din1724,
   output        cfg_din1725,
   output        cfg_din1726,
   output        cfg_din1727,
   output        cfg_din1728,
   output        cfg_din1729,
   output        cfg_din1730,
   output        cfg_din1731,
   output        cfg_din1732,
   output        cfg_din1733,
   output        cfg_din1734,
   output        cfg_din1735,
   output        cfg_din1736,
   output        cfg_din1737,
   output        cfg_din1738,
   output        cfg_din1739,
   output        cfg_din1740,
   output        cfg_din1741,
   output        cfg_din1742,
   output        cfg_din1743,
   output        cfg_din1744,
   output        cfg_din1745,
   output        cfg_din1746,
   output        cfg_din1747,
   output        cfg_din1748,
   output        cfg_din1749,
   output        cfg_din1750,
   output        cfg_din1751,
   output        cfg_din1752,
   output        cfg_din1753,
   output        cfg_din1754,
   output        cfg_din1755,
   output        cfg_din1756,
   output        cfg_din1757,
   output        cfg_din1758,
   output        cfg_din1759,
   output        cfg_din1760,
   output        cfg_din1761,
   output        cfg_din1762,
   output        cfg_din1763,
   output        cfg_din1764,
   output        cfg_din1765,
   output        cfg_din1766,
   output        cfg_din1767,
   output        cfg_din1768,
   output        cfg_din1769,
   output        cfg_din1770,
   output        cfg_din1771,
   output        cfg_din1772,
   output        cfg_din1773,
   output        cfg_din1774,
   output        cfg_din1775,
   output        cfg_din1776,
   output        cfg_din1777,
   output        cfg_din1778,
   output        cfg_din1779,
   output        cfg_din1780,
   output        cfg_din1781,
   output        cfg_din1782,
   output        cfg_din1783,
   output        cfg_din1784,
   output        cfg_din1785,
   output        cfg_din1786,
   output        cfg_din1787,
   output        cfg_din1788,
   output        cfg_din1789,
   output        cfg_din1790,
   output        cfg_din1791,
   output        cfg_din1792,
   output        cfg_din1793,
   output        cfg_din1794,
   output        cfg_din1795,
   output        cfg_din1796,
   output        cfg_din1797,
   output        cfg_din1798,
   output        cfg_din1799,
   output        cfg_din1800,
   output        cfg_din1801,
   output        cfg_din1802,
   output        cfg_din1803,
   output        cfg_din1804,
   output        cfg_din1805,
   output        cfg_din1806,
   output        cfg_din1807,
   output        cfg_din1808,
   output        cfg_din1809,
   output        cfg_din1810,
   output        cfg_din1811,
   output        cfg_din1812,
   output        cfg_din1813,
   output        cfg_din1814,
   output        cfg_din1815,
   output        cfg_din1816,
   output        cfg_din1817,
   output        cfg_din1818,
   output        cfg_din1819,
   output        cfg_din1820,
   output        cfg_din1821,
   output        cfg_din1822,
   output        cfg_din1823,
   output        cfg_din1824,
   output        cfg_din1825,
   output        cfg_din1826,
   output        cfg_din1827,
   output        cfg_din1828,
   output        cfg_din1829,
   output        cfg_din1830,
   output        cfg_din1831,
   output        cfg_din1832,
   output        cfg_din1833,
   output        cfg_din1834,
   output        cfg_din1835,
   output        cfg_din1836,
   output        cfg_din1837,
   output        cfg_din1838,
   output        cfg_din1839,
   output        cfg_din1840,
   output        cfg_din1841,
   output        cfg_din1842,
   output        cfg_din1843,
   output        cfg_din1844,
   output        cfg_din1845,
   output        cfg_din1846,
   output        cfg_din1847,
   output        cfg_din1848,
   output        cfg_din1849,
   output        cfg_din1850,
   output        cfg_din1851,
   output        cfg_din1852,
   output        cfg_din1853,
   output        cfg_din1854,
   output        cfg_din1855,
   output        cfg_din1856,
   output        cfg_din1857,
   output        cfg_din1858,
   output        cfg_din1859,
   output        cfg_din1860,
   output        cfg_din1861,
   output        cfg_din1862,
   output        cfg_din1863,
   output        cfg_din1864,
   output        cfg_din1865,
   output        cfg_din1866,
   output        cfg_din1867,
   output        cfg_din1868,
   output        cfg_din1869,
   output        cfg_din1870,
   output        cfg_din1871,
   output        cfg_din1872,
   output        cfg_din1873,
   output        cfg_din1874,
   output        cfg_din1875,
   output        cfg_din1876,
   output        cfg_din1877,
   output        cfg_din1878,
   output        cfg_din1879,
   output        cfg_din1880,
   output        cfg_din1881,
   output        cfg_din1882,
   output        cfg_din1883,
   output        cfg_din1884,
   output        cfg_din1885,
   output        cfg_din1886,
   output        cfg_din1887,
   output        cfg_din1888,
   output        cfg_din1889,
   output        cfg_din1890,
   output        cfg_din1891,
   output        cfg_din1892,
   output        cfg_din1893,
   output        cfg_din1894,
   output        cfg_din1895,
   output        cfg_din1896,
   output        cfg_din1897,
   output        cfg_din1898,
   output        cfg_din1899,
   output        cfg_din1900,
   output        cfg_din1901,
   output        cfg_din1902,
   output        cfg_din1903,
   output        cfg_din1904,
   output        cfg_din1905,
   output        cfg_din1906,
   output        cfg_din1907,
   output        cfg_din1908,
   output        cfg_din1909,
   output        cfg_din1910,
   output        cfg_din1911,
   output        cfg_din1912,
   output        cfg_din1913,
   output        cfg_din1914,
   output        cfg_din1915,
   output        cfg_din1916,
   output        cfg_din1917,
   output        cfg_din1918,
   output        cfg_din1919,
   output        cfg_din1920,
   output        cfg_din1921,
   output        cfg_din1922,
   output        cfg_din1923,
   output        cfg_din1924,
   output        cfg_din1925,
   output        cfg_din1926,
   output        cfg_din1927,
   output        cfg_din1928,
   output        cfg_din1929,
   output        cfg_din1930,
   output        cfg_din1931,
   output        cfg_din1932,
   output        cfg_din1933,
   output        cfg_din1934,
   output        cfg_din1935,
   output        cfg_din1936,
   output        cfg_din1937,
   output        cfg_din1938,
   output        cfg_din1939,
   output        cfg_din1940,
   output        cfg_din1941,
   output        cfg_din1942,
   output        cfg_din1943,
   output        cfg_din1944,
   output        cfg_din1945,
   output        cfg_din1946,
   output        cfg_din1947,
   output        cfg_din1948,
   output        cfg_din1949,
   output        cfg_din1950,
   output        cfg_din1951,
   output        cfg_din1952,
   output        cfg_din1953,
   output        cfg_din1954,
   output        cfg_din1955,
   output        cfg_din1956,
   output        cfg_din1957,
   output        cfg_din1958,
   output        cfg_din1959,
   output        cfg_din1960,
   output        cfg_din1961,
   output        cfg_din1962,
   output        cfg_din1963,
   output        cfg_din1964,
   output        cfg_din1965,
   output        cfg_din1966,
   output        cfg_din1967,
   output        cfg_din1968,
   output        cfg_din1969,
   output        cfg_din1970,
   output        cfg_din1971,
   output        cfg_din1972,
   output        cfg_din1973,
   output        cfg_din1974,
   output        cfg_din1975,
   output        cfg_din1976,
   output        cfg_din1977,
   output        cfg_din1978,
   output        cfg_din1979,
   output        cfg_din1980,
   output        cfg_din1981,
   output        cfg_din1982,
   output        cfg_din1983,
   output        cfg_din1984,
   output        cfg_din1985,
   output        cfg_din1986,
   output        cfg_din1987,
   output        cfg_din1988,
   output        cfg_din1989,
   output        cfg_din1990,
   output        cfg_din1991,
   output        cfg_din1992,
   output        cfg_din1993,
   output        cfg_din1994,
   output        cfg_din1995,
   output        cfg_din1996,
   output        cfg_din1997,
   output        cfg_din1998,
   output        cfg_din1999,
   output        cfg_din2000,
   output        cfg_din2001,
   output        cfg_din2002,
   output        cfg_din2003,
   output        cfg_din2004,
   output        cfg_din2005,
   output        cfg_din2006,
   output        cfg_din2007,
   output        cfg_din2008,
   output        cfg_din2009,
   output        cfg_din2010,
   output        cfg_din2011,
   output        cfg_din2012,
   output        cfg_din2013,
   output        cfg_din2014,
   output        cfg_din2015,
   output        cfg_din2016,
   output        cfg_din2017,
   output        cfg_din2018,
   output        cfg_din2019,
   output        cfg_din2020,
   output        cfg_din2021,
   output        cfg_din2022,
   output        cfg_din2023,
   output        cfg_din2024,
   output        cfg_din2025,
   output        cfg_din2026,
   output        cfg_din2027,
   output        cfg_din2028,
   output        cfg_din2029,
   output        cfg_din2030,
   output        cfg_din2031,
   output        cfg_din2032,
   output        cfg_din2033,
   output        cfg_din2034,
   output        cfg_din2035,
   output        cfg_din2036,
   output        cfg_din2037,
   output        cfg_din2038,
   output        cfg_din2039,
   output        cfg_din2040,
   output        cfg_din2041,
   output        cfg_din2042,
   output        cfg_din2043,
   output        cfg_din2044,
   output        cfg_din2045,
   output        cfg_din2046,
   output        cfg_din2047,
   output        cfg_din2048,
   output        cfg_din2049,
   output        cfg_din2050,
   output        cfg_din2051,
   output        cfg_din2052,
   output        cfg_din2053,
   output        cfg_din2054,
   output        cfg_din2055,
   output        cfg_din2056,
   output        cfg_din2057,
   output        cfg_din2058,
   output        cfg_din2059,
   output        cfg_din2060,
   output        cfg_din2061,
   output        cfg_din2062,
   output        cfg_din2063,
   output        cfg_din2064,
   output        cfg_din2065,
   output        cfg_din2066,
   output        cfg_din2067,
   output        cfg_din2068,
   output        cfg_din2069,
   output        cfg_din2070,
   output        cfg_din2071,
   output        cfg_din2072,
   output        cfg_din2073,
   output        cfg_din2074,
   output        cfg_din2075,
   output        cfg_din2076,
   output        cfg_din2077,
   output        cfg_din2078,
   output        cfg_din2079,
   output        cfg_din2080,
   output        cfg_din2081,
   output        cfg_din2082,
   output        cfg_din2083,
   output        cfg_din2084,
   output        cfg_din2085,
   output        cfg_din2086,
   output        cfg_din2087,
   output        cfg_din2088,
   output        cfg_din2089,
   output        cfg_din2090,
   output        cfg_din2091,
   output        cfg_din2092,
   output        cfg_din2093,
   output        cfg_din2094,
   output        cfg_din2095,
   output        cfg_din2096,
   output        cfg_din2097,
   output        cfg_din2098,
   output        cfg_din2099,
   output        cfg_din2100,
   output        cfg_din2101,
   output        cfg_din2102,
   output        cfg_din2103,
   output        cfg_din2104,
   output        cfg_din2105,
   output        cfg_din2106,
   output        cfg_din2107,
   output        cfg_din2108,
   output        cfg_din2109,
   output        cfg_din2110,
   output        cfg_din2111,
   output        cfg_din2112,
   output        cfg_din2113,
   output        cfg_din2114,
   output        cfg_din2115,
   output        cfg_din2116,
   output        cfg_din2117,
   output        cfg_din2118,
   output        cfg_din2119,
   output        cfg_din2120,
   output        cfg_din2121,
   output        cfg_din2122,
   output        cfg_din2123,
   output        cfg_din2124,
   output        cfg_din2125,
   output        cfg_din2126,
   output        cfg_din2127,
   output        cfg_din2128,
   output        cfg_din2129,
   output        cfg_din2130,
   output        cfg_din2131,
   output        cfg_din2132,
   output        cfg_din2133,
   output        cfg_din2134,
   output        cfg_din2135,
   output        cfg_din2136,
   output        cfg_din2137,
   output        cfg_din2138,
   output        cfg_din2139,
   output        cfg_din2140,
   output        cfg_din2141,
   output        cfg_din2142,
   output        cfg_din2143,
   output        cfg_din2144,
   output        cfg_din2145,
   output        cfg_din2146,
   output        cfg_din2147,
   output        cfg_din2148,
   output        cfg_din2149,
   output        cfg_din2150,
   output        cfg_din2151,
   output        cfg_din2152,
   output        cfg_din2153,
   output        cfg_din2154,
   output        cfg_din2155,
   output        cfg_din2156,
   output        cfg_din2157,
   output        cfg_din2158,
   output        cfg_din2159,
   output        cfg_din2160,
   output        cfg_din2161,
   output        cfg_din2162,
   output        cfg_din2163,
   output        cfg_din2164,
   output        cfg_din2165,
   output        cfg_din2166,
   output        cfg_din2167,
   output        cfg_din2168,
   output        cfg_din2169,
   output        cfg_din2170,
   output        cfg_din2171,
   output        cfg_din2172,
   output        cfg_din2173,
   output        cfg_din2174,
   output        cfg_din2175,
   output        cfg_din2176,
   output        cfg_din2177,
   output        cfg_din2178,
   output        cfg_din2179,
   output        cfg_din2180,
   output        cfg_din2181,
   output        cfg_din2182,
   output        cfg_din2183,
   output        cfg_din2184,
   output        cfg_din2185,
   output        cfg_din2186,
   output        cfg_din2187,
   output        cfg_din2188,
   output        cfg_din2189,
   output        cfg_din2190,
   output        cfg_din2191,
   output        cfg_din2192,
   output        cfg_din2193,
   output        cfg_din2194,
   output        cfg_din2195,
   output        cfg_din2196,
   output        cfg_din2197,
   output        cfg_din2198,
   output        cfg_din2199,
   output        cfg_din2200,
   output        cfg_din2201,
   output        cfg_din2202,
   output        cfg_din2203,
   output        cfg_din2204,
   output        cfg_din2205,
   output        cfg_din2206,
   output        cfg_din2207,
   output        cfg_din2208,
   output        cfg_din2209,
   output        cfg_din2210,
   output        cfg_din2211,
   output        cfg_din2212,
   output        cfg_din2213,
   output        cfg_din2214,
   output        cfg_din2215,
   output        cfg_din2216,
   output        cfg_din2217,
   output        cfg_din2218,
   output        cfg_din2219,
   output        cfg_din2220,
   output        cfg_din2221,
   output        cfg_din2222,
   output        cfg_din2223,
   output        cfg_din2224,
   output        cfg_din2225,
   output        cfg_din2226,
   output        cfg_din2227,
   output        cfg_din2228,
   output        cfg_din2229,
   output        cfg_din2230,
   output        cfg_din2231,
   output        cfg_din2232,
   output        cfg_din2233,
   output        cfg_din2234,
   output        cfg_din2235,
   output        cfg_din2236,
   output        cfg_din2237,
   output        cfg_din2238,
   output        cfg_din2239,
   output        cfg_din2240,
   output        cfg_din2241,
   output        cfg_din2242,
   output        cfg_din2243,
   output        cfg_din2244,
   output        cfg_din2245,
   output        cfg_din2246,
   output        cfg_din2247,
   output        cfg_din2248,
   output        cfg_din2249,
   output        cfg_din2250,
   output        cfg_din2251,
   output        cfg_din2252,
   output        cfg_din2253,
   output        cfg_din2254,
   output        cfg_din2255,
   output        cfg_din2256,
   output        cfg_din2257,
   output        cfg_din2258,
   output        cfg_din2259,
   output        cfg_din2260,
   output        cfg_din2261,
   output        cfg_din2262,
   output        cfg_din2263,
   output        cfg_din2264,
   output        cfg_din2265,
   output        cfg_din2266,
   output        cfg_din2267,
   output        cfg_din2268,
   output        cfg_din2269,
   output        cfg_din2270,
   output        cfg_din2271,
   output        cfg_din2272,
   output        cfg_din2273,
   output        cfg_din2274,
   output        cfg_din2275,
   output        cfg_din2276,
   output        cfg_din2277,
   output        cfg_din2278,
   output        cfg_din2279,
   output        cfg_din2280,
   output        cfg_din2281,
   output        cfg_din2282,
   output        cfg_din2283,
   output        cfg_din2284,
   output        cfg_din2285,
   output        cfg_din2286,
   output        cfg_din2287,
   output        cfg_din2288,
   output        cfg_din2289,
   output        cfg_din2290,
   output        cfg_din2291,
   output        cfg_din2292,
   output        cfg_din2293,
   output        cfg_din2294,
   output        cfg_din2295,
   output        cfg_din2296,
   output        cfg_din2297,
   output        cfg_din2298,
   output        cfg_din2299,
   output        cfg_din2300,
   output        cfg_din2301,
   output        cfg_din2302,
   output        cfg_din2303,
   output        cfg_din2304,
   output        cfg_din2305,
   output        cfg_din2306,
   output        cfg_din2307,
   output        cfg_din2308,
   output        cfg_din2309,
   output        cfg_din2310,
   output        cfg_din2311,
   output        cfg_din2312,
   output        cfg_din2313,
   output        cfg_din2314,
   output        cfg_din2315,
   output        cfg_din2316,
   output        cfg_din2317,
   output        cfg_din2318,
   output        cfg_din2319,
   output        cfg_din2320,
   output        cfg_din2321,
   output        cfg_din2322,
   output        cfg_din2323,
   output        cfg_din2324,
   output        cfg_din2325,
   output        cfg_din2326,
   output        cfg_din2327,
   output        cfg_din2328,
   output        cfg_din2329,
   output        cfg_din2330,
   output        cfg_din2331,
   output        cfg_din2332,
   output        cfg_din2333,
   output        cfg_din2334,
   output        cfg_din2335,
   output        cfg_din2336,
   output        cfg_din2337,
   output        cfg_din2338,
   output        cfg_din2339,
   output        cfg_din2340,
   output        cfg_din2341,
   output        cfg_din2342,
   output        cfg_din2343,
   output        cfg_din2344,
   output        cfg_din2345,
   output        cfg_din2346,
   output        cfg_din2347,
   output        cfg_din2348,
   output        cfg_din2349,
   output        cfg_din2350,
   output        cfg_din2351,
   output        cfg_din2352,
   output        cfg_din2353,
   output        cfg_din2354,
   output        cfg_din2355,
   output        cfg_din2356,
   output        cfg_din2357,
   output        cfg_din2358,
   output        cfg_din2359,
   output        cfg_din2360,
   output        cfg_din2361,
   output        cfg_din2362,
   output        cfg_din2363,
   output        cfg_din2364,
   output        cfg_din2365,
   output        cfg_din2366,
   output        cfg_din2367,
   output        cfg_din2368,
   output        cfg_din2369,
   output        cfg_din2370,
   output        cfg_din2371,
   output        cfg_din2372,
   output        cfg_din2373,
   output        cfg_din2374,
   output        cfg_din2375,
   output        cfg_din2376,
   output        cfg_din2377,
   output        cfg_din2378,
   output        cfg_din2379,
   output        cfg_din2380,
   output        cfg_din2381,
   output        cfg_din2382,
   output        cfg_din2383,
   output        cfg_din2384,
   output        cfg_din2385,
   output        cfg_din2386,
   output        cfg_din2387,
   output        cfg_din2388,
   output        cfg_din2389,
   output        cfg_din2390,
   output        cfg_din2391,
   output        cfg_din2392,
   output        cfg_din2393,
   output        cfg_din2394,
   output        cfg_din2395,
   output        cfg_din2396,
   output        cfg_din2397,
   output        cfg_din2398,
   output        cfg_din2399,
   output        cfg_din2400,
   output        cfg_din2401,
   output        cfg_din2402,
   output        cfg_din2403,
   output        cfg_din2404,
   output        cfg_din2405,
   output        cfg_din2406,
   output        cfg_din2407,
   output        cfg_din2408,
   output        cfg_din2409,
   output        cfg_din2410,
   output        cfg_din2411,
   output        cfg_din2412,
   output        cfg_din2413,
   output        cfg_din2414,
   output        cfg_din2415,
   output        cfg_din2416,
   output        cfg_din2417,
   output        cfg_din2418,
   output        cfg_din2419,
   output        cfg_din2420,
   output        cfg_din2421,
   output        cfg_din2422,
   output        cfg_din2423,
   output        cfg_din2424,
   output        cfg_din2425,
   output        cfg_din2426,
   output        cfg_din2427,
   output        cfg_din2428,
   output        cfg_din2429,
   output        cfg_din2430,
   output        cfg_din2431,
   output        cfg_din2432,
   output        cfg_din2433,
   output        cfg_din2434,
   output        cfg_din2435,
   output        cfg_din2436,
   output        cfg_din2437,
   output        cfg_din2438,
   output        cfg_din2439,
   output        cfg_din2440,
   output        cfg_din2441,
   output        cfg_din2442,
   output        cfg_din2443,
   output        cfg_din2444,
   output        cfg_din2445,
   output        cfg_din2446,
   output        cfg_din2447,
   output        cfg_din2448,
   output        cfg_din2449,
   output        cfg_din2450,
   output        cfg_din2451,
   output        cfg_din2452,
   output        cfg_din2453,
   output        cfg_din2454,
   output        cfg_din2455,
   output        cfg_din2456,
   output        cfg_din2457,
   output        cfg_din2458,
   output        cfg_din2459,
   output        cfg_din2460,
   output        cfg_din2461,
   output        cfg_din2462,
   output        cfg_din2463,
   output        cfg_din2464,
   output        cfg_din2465,
   output        cfg_din2466,
   output        cfg_din2467,
   output        cfg_din2468,
   output        cfg_din2469,
   output        cfg_din2470,
   output        cfg_din2471,
   output        cfg_din2472,
   output        cfg_din2473,
   output        cfg_din2474,
   output        cfg_din2475,
   output        cfg_din2476,
   output        cfg_din2477,
   output        cfg_din2478,
   output        cfg_din2479,
   output        cfg_din2480,
   output        cfg_din2481,
   output        cfg_din2482,
   output        cfg_din2483,
   output        cfg_din2484,
   output        cfg_din2485,
   output        cfg_din2486,
   output        cfg_din2487,
   output        cfg_din2488,
   output        cfg_din2489,
   output        cfg_din2490,
   output        cfg_din2491,
   output        cfg_din2492,
   output        cfg_din2493,
   output        cfg_din2494,
   output        cfg_din2495,
   output        cfg_din2496,
   output        cfg_din2497,
   output        cfg_din2498,
   output        cfg_din2499,
   output        cfg_din2500,
   output        cfg_din2501,
   output        cfg_din2502,
   output        cfg_din2503,
   output        cfg_din2504,
   output        cfg_din2505,
   output        cfg_din2506,
   output        cfg_din2507,
   output        cfg_din2508,
   output        cfg_din2509,
   output        cfg_din2510,
   output        cfg_din2511,
   output        cfg_din2512,
   output        cfg_din2513,
   output        cfg_din2514,
   output        cfg_din2515,
   output        cfg_din2516,
   output        cfg_din2517,
   output        cfg_din2518,
   output        cfg_din2519,
   output        cfg_din2520,
   output        cfg_din2521,
   output        cfg_din2522,
   output        cfg_din2523,
   output        cfg_din2524,
   output        cfg_din2525,
   output        cfg_din2526,
   output        cfg_din2527,
   output        cfg_din2528,
   output        cfg_din2529,
   output        cfg_din2530,
   output        cfg_din2531,
   output        cfg_din2532,
   output        cfg_din2533,
   output        cfg_din2534,
   output        cfg_din2535,
   output        cfg_din2536,
   output        cfg_din2537,
   output        cfg_din2538,
   output        cfg_din2539,
   output        cfg_din2540,
   output        cfg_din2541,
   output        cfg_din2542,
   output        cfg_din2543,
   output        cfg_din2544,
   output        cfg_din2545,
   output        cfg_din2546,
   output        cfg_din2547,
   output        cfg_din2548,
   output        cfg_din2549,
   output        cfg_din2550,
   output        cfg_din2551,
   output        cfg_din2552,
   output        cfg_din2553,
   output        cfg_din2554,
   output        cfg_din2555,
   output        cfg_din2556,
   output        cfg_din2557,
   output        cfg_din2558,
   output        cfg_din2559,
   output        cfg_din2560,
   output        cfg_din2561,
   output        cfg_din2562,
   output        cfg_din2563,
   output        cfg_din2564,
   output        cfg_din2565,
   output        cfg_din2566,
   output        cfg_din2567,
   output        cfg_din2568,
   output        cfg_din2569,
   output        cfg_din2570,
   output        cfg_din2571,
   output        cfg_din2572,
   output        cfg_din2573,
   output        cfg_din2574,
   output        cfg_din2575,
   output        cfg_din2576,
   output        cfg_din2577,
   output        cfg_din2578,
   output        cfg_din2579,
   output        cfg_din2580,
   output        cfg_din2581,
   output        cfg_din2582,
   output        cfg_din2583,
   output        cfg_din2584,
   output        cfg_din2585,
   output        cfg_din2586,
   output        cfg_din2587,
   output        cfg_din2588,
   output        cfg_din2589,
   output        cfg_din2590,
   output        cfg_din2591,
   output        cfg_din2592,
   output        cfg_din2593,
   output        cfg_din2594,
   output        cfg_din2595,
   output        cfg_din2596,
   output        cfg_din2597,
   output        cfg_din2598,
   output        cfg_din2599,
   output        cfg_din2600,
   output        cfg_din2601,
   output        cfg_din2602,
   output        cfg_din2603,
   output        cfg_din2604,
   output        cfg_din2605,
   output        cfg_din2606,
   output        cfg_din2607,
   output        cfg_din2608,
   output        cfg_din2609,
   output        cfg_din2610,
   output        cfg_din2611,
   output        cfg_din2612,
   output        cfg_din2613,
   output        cfg_din2614,
   output        cfg_din2615,
   output        cfg_din2616,
   output        cfg_din2617,
   output        cfg_din2618,
   output        cfg_din2619,
   output        cfg_din2620,
   output        cfg_din2621,
   output        cfg_din2622,
   output        cfg_din2623,
   output        cfg_din2624,
   output        cfg_din2625,
   output        cfg_din2626,
   output        cfg_din2627,
   output        cfg_din2628,
   output        cfg_din2629,
   output        cfg_din2630,
   output        cfg_din2631,
   output        cfg_din2632,
   output        cfg_din2633,
   output        cfg_din2634,
   output        cfg_din2635,
   output        cfg_din2636,
   output        cfg_din2637,
   output        cfg_din2638,
   output        cfg_din2639,
   output        cfg_din2640,
   output        cfg_din2641,
   output        cfg_din2642,
   output        cfg_din2643,
   output        cfg_din2644,
   output        cfg_din2645,
   output        cfg_din2646,
   output        cfg_din2647,
   output        cfg_din2648,
   output        cfg_din2649,
   output        cfg_din2650,
   output        cfg_din2651,
   output        cfg_din2652,
   output        cfg_din2653,
   output        cfg_din2654,
   output        cfg_din2655,
   output        cfg_din2656,
   output        cfg_din2657,
   output        cfg_din2658,
   output        cfg_din2659,
   output        cfg_din2660,
   output        cfg_din2661,
   output        cfg_din2662,
   output        cfg_din2663,
   output        cfg_din2664,
   output        cfg_din2665,
   output        cfg_din2666,
   output        cfg_din2667,
   output        cfg_din2668,
   output        cfg_din2669,
   output        cfg_din2670,
   output        cfg_din2671,
   output        cfg_din2672,
   output        cfg_din2673,
   output        cfg_din2674,
   output        cfg_din2675,
   output        cfg_din2676,
   output        cfg_din2677,
   output        cfg_din2678,
   output        cfg_din2679,
   output        cfg_din2680,
   output        cfg_din2681,
   output        cfg_din2682,
   output        cfg_din2683,
   output        cfg_din2684,
   output        cfg_din2685,
   output        cfg_din2686,
   output        cfg_din2687,
   output        cfg_din2688,
   output        cfg_din2689,
   output        cfg_din2690,
   output        cfg_din2691,
   output        cfg_din2692,
   output        cfg_din2693,
   output        cfg_din2694,
   output        cfg_din2695,
   output        cfg_din2696,
   output        cfg_din2697,
   output        cfg_din2698,
   output        cfg_din2699,
   output        cfg_din2700,
   output        cfg_din2701,
   output        cfg_din2702,
   output        cfg_din2703,
   output        cfg_din2704,
   output        cfg_din2705,
   output        cfg_din2706,
   output        cfg_din2707,
   output        cfg_din2708,
   output        cfg_din2709,
   output        cfg_din2710,
   output        cfg_din2711,
   output        cfg_din2712,
   output        cfg_din2713,
   output        cfg_din2714,
   output        cfg_din2715,
   output        cfg_din2716,
   output        cfg_din2717,
   output        cfg_din2718,
   output        cfg_din2719,
   output        cfg_din2720,
   output        cfg_din2721,
   output        cfg_din2722,
   output        cfg_din2723,
   output        cfg_din2724,
   output        cfg_din2725,
   output        cfg_din2726,
   output        cfg_din2727,
   output        cfg_din2728,
   output        cfg_din2729,
   output        cfg_din2730,
   output        cfg_din2731,
   output        cfg_din2732,
   output        cfg_din2733,
   output        cfg_din2734,
   output        cfg_din2735,
   output        cfg_din2736,
   output        cfg_din2737,
   output        cfg_din2738,
   output        cfg_din2739,
   output        cfg_din2740,
   output        cfg_din2741,
   output        cfg_din2742,
   output        cfg_din2743,
   output        cfg_din2744,
   output        cfg_din2745,
   output        cfg_din2746,
   output        cfg_din2747,
   output        cfg_din2748,
   output        cfg_din2749,
   output        cfg_din2750,
   output        cfg_din2751,
   output        cfg_din2752,
   output        cfg_din2753,
   output        cfg_din2754,
   output        cfg_din2755,
   output        cfg_din2756,
   output        cfg_din2757,
   output        cfg_din2758,
   output        cfg_din2759,
   output        cfg_din2760,
   output        cfg_din2761,
   output        cfg_din2762,
   output        cfg_din2763,
   output        cfg_din2764,
   output        cfg_din2765,
   output        cfg_din2766,
   output        cfg_din2767,
   output        cfg_din2768,
   output        cfg_din2769,
   output        cfg_din2770,
   output        cfg_din2771,
   output        cfg_din2772,
   output        cfg_din2773,
   output        cfg_din2774,
   output        cfg_din2775,
   output        cfg_din2776,
   output        cfg_din2777,
   output        cfg_din2778,
   output        cfg_din2779,
   output        cfg_din2780,
   output        cfg_din2781,
   output        cfg_din2782,
   output        cfg_din2783,
   output        cfg_din2784,
   output        cfg_din2785,
   output        cfg_din2786,
   output        cfg_din2787,
   output        cfg_din2788,
   output        cfg_din2789,
   output        cfg_din2790,
   output        cfg_din2791,
   output        cfg_din2792,
   output        cfg_din2793,
   output        cfg_din2794,
   output        cfg_din2795,
   output        cfg_din2796,
   output        cfg_din2797,
   output        cfg_din2798,
   output        cfg_din2799,
   output        cfg_din2800,
   output        cfg_din2801,
   output        cfg_din2802,
   output        cfg_din2803,
   output        cfg_din2804,
   output        cfg_din2805,
   output        cfg_din2806,
   output        cfg_din2807,
   output        cfg_din2808,
   output        cfg_din2809,
   output        cfg_din2810,
   output        cfg_din2811,
   output        cfg_din2812,
   output        cfg_din2813,
   output        cfg_din2814,
   output        cfg_din2815,
   output        cfg_din2816,
   output        cfg_din2817,
   output        cfg_din2818,
   output        cfg_din2819,
   output        cfg_din2820,
   output        cfg_din2821,
   output        cfg_din2822,
   output        cfg_din2823,
   output        cfg_din2824,
   output        cfg_din2825,
   output        cfg_din2826,
   output        cfg_din2827,
   output        cfg_din2828,
   output        cfg_din2829,
   output        cfg_din2830,
   output        cfg_din2831,
   output        cfg_din2832,
   output        cfg_din2833,
   output        cfg_din2834,
   output        cfg_din2835,
   output        cfg_din2836,
   output        cfg_din2837,
   output        cfg_din2838,
   output        cfg_din2839,
   output        cfg_din2840,
   output        cfg_din2841,
   output        cfg_din2842,
   output        cfg_din2843,
   output        cfg_din2844,
   output        cfg_din2845,
   output        cfg_din2846,
   output        cfg_din2847,
   output        cfg_din2848,
   output        cfg_din2849,
   output        cfg_din2850,
   output        cfg_din2851,
   output        cfg_din2852,
   output        cfg_din2853,
   output        cfg_din2854,
   output        cfg_din2855,
   output        cfg_din2856,
   output        cfg_din2857,
   output        cfg_din2858,
   output        cfg_din2859,
   output        cfg_din2860,
   output        cfg_din2861,
   output        cfg_din2862,
   output        cfg_din2863,
   output        cfg_din2864,
   output        cfg_din2865,
   output        cfg_din2866,
   output        cfg_din2867,
   output        cfg_din2868,
   output        cfg_din2869,
   output        cfg_din2870,
   output        cfg_din2871,
   output        cfg_din2872,
   output        cfg_din2873,
   output        cfg_din2874,
   output        cfg_din2875,
   output        cfg_din2876,
   output        cfg_din2877,
   output        cfg_din2878,
   output        cfg_din2879,
   output        cfg_din2880,
   output        cfg_din2881,
   output        cfg_din2882,
   output        cfg_din2883,
   output        cfg_din2884,
   output        cfg_din2885,
   output        cfg_din2886,
   output        cfg_din2887,
   output        cfg_din2888,
   output        cfg_din2889,
   output        cfg_din2890,
   output        cfg_din2891,
   output        cfg_din2892,
   output        cfg_din2893,
   output        cfg_din2894,
   output        cfg_din2895,
   output        cfg_din2896,
   output        cfg_din2897,
   output        cfg_din2898,
   output        cfg_din2899,
   output        cfg_din2900,
   output        cfg_din2901,
   output        cfg_din2902,
   output        cfg_din2903,
   output        cfg_din2904,
   output        cfg_din2905,
   output        cfg_din2906,
   output        cfg_din2907,
   output        cfg_din2908,
   output        cfg_din2909,
   output        cfg_din2910,
   output        cfg_din2911,
   output        cfg_din2912,
   output        cfg_din2913,
   output        cfg_din2914,
   output        cfg_din2915,
   output        cfg_din2916,
   output        cfg_din2917,
   output        cfg_din2918,
   output        cfg_din2919,
   output        cfg_din2920,
   output        cfg_din2921,
   output        cfg_din2922,
   output        cfg_din2923,
   output        cfg_din2924,
   output        cfg_din2925,
   output        cfg_din2926,
   output        cfg_din2927,
   output        cfg_din2928,
   output        cfg_din2929,
   output        cfg_din2930,
   output        cfg_din2931,
   output        cfg_din2932,
   output        cfg_din2933,
   output        cfg_din2934,
   output        cfg_din2935,
   output        cfg_din2936,
   output        cfg_din2937,
   output        cfg_din2938,
   output        cfg_din2939,
   output        cfg_din2940,
   output        cfg_din2941,
   output        cfg_din2942,
   output        cfg_din2943,
   output        cfg_din2944,
   output        cfg_din2945,
   output        cfg_din2946,
   output        cfg_din2947,
   output        cfg_din2948,
   output        cfg_din2949,
   output        cfg_din2950,
   output        cfg_din2951,
   output        cfg_din2952,
   output        cfg_din2953,
   output        cfg_din2954,
   output        cfg_din2955,
   output        cfg_din2956,
   output        cfg_din2957,
   output        cfg_din2958,
   output        cfg_din2959,
   output        cfg_din2960,
   output        cfg_din2961,
   output        cfg_din2962,
   output        cfg_din2963,
   output        cfg_din2964,
   output        cfg_din2965,
   output        cfg_din2966,
   output        cfg_din2967,
   output        cfg_din2968,
   output        cfg_din2969,
   output        cfg_din2970,
   output        cfg_din2971,
   output        cfg_din2972,
   output        cfg_din2973,
   output        cfg_din2974,
   output        cfg_din2975,
   output        cfg_din2976,
   output        cfg_din2977,
   output        cfg_din2978,
   output        cfg_din2979,
   output        cfg_din2980,
   output        cfg_din2981,
   output        cfg_din2982,
   output        cfg_din2983,
   output        cfg_din2984,
   output        cfg_din2985,
   output        cfg_din2986,
   output        cfg_din2987,
   output        cfg_din2988,
   output        cfg_din2989,
   output        cfg_din2990,
   output        cfg_din2991,
   output        cfg_din2992,
   output        cfg_din2993,
   output        cfg_din2994,
   output        cfg_din2995,
   output        cfg_din2996,
   output        cfg_din2997,
   output        cfg_din2998,
   output        cfg_din2999,
   output        cfg_din3000,
   output        cfg_din3001,
   output        cfg_din3002,
   output        cfg_din3003,
   output        cfg_din3004,
   output        cfg_din3005,
   output        cfg_din3006,
   output        cfg_din3007,
   output        cfg_din3008,
   output        cfg_din3009,
   output        cfg_din3010,
   output        cfg_din3011,
   output        cfg_din3012,
   output        cfg_din3013,
   output        cfg_din3014,
   output        cfg_din3015,
   output        cfg_din3016,
   output        cfg_din3017,
   output        cfg_din3018,
   output        cfg_din3019,
   output        cfg_din3020,
   output        cfg_din3021,
   output        cfg_din3022,
   output        cfg_din3023,
   output        cfg_din3024,
   output        cfg_din3025,
   output        cfg_din3026,
   output        cfg_din3027,
   output        cfg_din3028,
   output        cfg_din3029,
   output        cfg_din3030,
   output        cfg_din3031,
   output        cfg_din3032,
   output        cfg_din3033,
   output        cfg_din3034,
   output        cfg_din3035,
   output        cfg_din3036,
   output        cfg_din3037,
   output        cfg_din3038,
   output        cfg_din3039,
   output        cfg_din3040,
   output        cfg_din3041,
   output        cfg_din3042,
   output        cfg_din3043,
   output        cfg_din3044,
   output        cfg_din3045,
   output        cfg_din3046,
   output        cfg_din3047,
   output        cfg_din3048,
   output        cfg_din3049,
   output        cfg_din3050,
   output        cfg_din3051,
   output        cfg_din3052,
   output        cfg_din3053,
   output        cfg_din3054,
   output        cfg_din3055,
   output        cfg_din3056,
   output        cfg_din3057,
   output        cfg_din3058,
   output        cfg_din3059,
   output        cfg_din3060,
   output        cfg_din3061,
   output        cfg_din3062,
   output        cfg_din3063,
   output        cfg_din3064,
   output        cfg_din3065,
   output        cfg_din3066,
   output        cfg_din3067,
   output        cfg_din3068,
   output        cfg_din3069,
   output        cfg_din3070,
   output        cfg_din3071,
   output        cfg_din3072,
   output        cfg_din3073,
   output        cfg_din3074,
   output        cfg_din3075,
   output        cfg_din3076,
   output        cfg_din3077,
   output        cfg_din3078,
   output        cfg_din3079,
   output        cfg_din3080,
   output        cfg_din3081,
   output        cfg_din3082,
   output        cfg_din3083,
   output        cfg_din3084,
   output        cfg_din3085,
   output        cfg_din3086,
   output        cfg_din3087,
   output        cfg_din3088,
   output        cfg_din3089,
   output        cfg_din3090,
   output        cfg_din3091,
   output        cfg_din3092,
   output        cfg_din3093,
   output        cfg_din3094,
   output        cfg_din3095,
   output        cfg_din3096,
   output        cfg_din3097,
   output        cfg_din3098,
   output        cfg_din3099,
   output        cfg_din3100,
   output        cfg_din3101,
   output        cfg_din3102,
   output        cfg_din3103,
   output        cfg_din3104,
   output        cfg_din3105,
   output        cfg_din3106,
   output        cfg_din3107,
   output        cfg_din3108,
   output        cfg_din3109,
   output        cfg_din3110,
   output        cfg_din3111,
   output        cfg_din3112,
   output        cfg_din3113,
   output        cfg_din3114,
   output        cfg_din3115,
   output        cfg_din3116,
   output        cfg_din3117,
   output        cfg_din3118,
   output        cfg_din3119,
   output        cfg_din3120,
   output        cfg_din3121,
   output        cfg_din3122,
   output        cfg_din3123,
   output        cfg_din3124,
   output        cfg_din3125,
   output        cfg_din3126,
   output        cfg_din3127,
   output        cfg_din3128,
   output        cfg_din3129,
   output        cfg_din3130,
   output        cfg_din3131,
   output        cfg_din3132,
   output        cfg_din3133,
   output        cfg_din3134,
   output        cfg_din3135,
   output        cfg_din3136,
   output        cfg_din3137,
   output        cfg_din3138,
   output        cfg_din3139,
   output        cfg_din3140,
   output        cfg_din3141,
   output        cfg_din3142,
   output        cfg_din3143,
   output        cfg_din3144,
   output        cfg_din3145,
   output        cfg_din3146,
   output        cfg_din3147,
   output        cfg_din3148,
   output        cfg_din3149,
   output        cfg_din3150,
   output        cfg_din3151,
   output        cfg_din3152,
   output        cfg_din3153,
   output        cfg_din3154,
   output        cfg_din3155,
   output        cfg_din3156,
   output        cfg_din3157,
   output        cfg_din3158,
   output        cfg_din3159,
   output        cfg_din3160,
   output        cfg_din3161,
   output        cfg_din3162,
   output        cfg_din3163,
   output        cfg_din3164,
   output        cfg_din3165,
   output        cfg_din3166,
   output        cfg_din3167,
   output        cfg_din3168,
   output        cfg_din3169,
   output        cfg_din3170,
   output        cfg_din3171,
   output        cfg_din3172,
   output        cfg_din3173,
   output        cfg_din3174,
   output        cfg_din3175,
   output        cfg_din3176,
   output        cfg_din3177,
   output        cfg_din3178,
   output        cfg_din3179,
   output        cfg_din3180,
   output        cfg_din3181,
   output        cfg_din3182,
   output        cfg_din3183,
   output        cfg_din3184,
   output        cfg_din3185,
   output        cfg_din3186,
   output        cfg_din3187,
   output        cfg_din3188,
   output        cfg_din3189,
   output        cfg_din3190,
   output        cfg_din3191,
   output        cfg_din3192,
   output        cfg_din3193,
   output        cfg_din3194,
   output        cfg_din3195,
   output        cfg_din3196,
   output        cfg_din3197,
   output        cfg_din3198,
   output        cfg_din3199,
   output        cfg_din3200,
   output        cfg_din3201,
   output        cfg_din3202,
   output        cfg_din3203,
   output        cfg_din3204,
   output        cfg_din3205,
   output        cfg_din3206,
   output        cfg_din3207,
   output        cfg_din3208,
   output        cfg_din3209,
   output        cfg_din3210,
   output        cfg_din3211,
   output        cfg_din3212,
   output        cfg_din3213,
   output        cfg_din3214,
   output        cfg_din3215,
   output        cfg_din3216,
   output        cfg_din3217,
   output        cfg_din3218,
   output        cfg_din3219,
   output        cfg_din3220,
   output        cfg_din3221,
   output        cfg_din3222,
   output        cfg_din3223,
   output        cfg_din3224,
   output        cfg_din3225,
   output        cfg_din3226,
   output        cfg_din3227,
   output        cfg_din3228,
   output        cfg_din3229,
   output        cfg_din3230,
   output        cfg_din3231,
   output        cfg_din3232,
   output        cfg_din3233,
   output        cfg_din3234,
   output        cfg_din3235,
   output        cfg_din3236,
   output        cfg_din3237,
   output        cfg_din3238,
   output        cfg_din3239,
   output        cfg_din3240,
   output        cfg_din3241,
   output        cfg_din3242,
   output        cfg_din3243,
   output        cfg_din3244,
   output        cfg_din3245,
   output        cfg_din3246,
   output        cfg_din3247,
   output        cfg_din3248,
   output        cfg_din3249,
   output        cfg_din3250,
   output        cfg_din3251,
   output        cfg_din3252,
   output        cfg_din3253,
   output        cfg_din3254,
   output        cfg_din3255,
   output        cfg_din3256,
   output        cfg_din3257,
   output        cfg_din3258,
   output        cfg_din3259,
   output        cfg_din3260,
   output        cfg_din3261,
   output        cfg_din3262,
   output        cfg_din3263,
   output        cfg_din3264,
   output        cfg_din3265,
   output        cfg_din3266,
   output        cfg_din3267,
   output        cfg_din3268,
   output        cfg_din3269,
   output        cfg_din3270,
   output        cfg_din3271,
   output        cfg_din3272,
   output        cfg_din3273,
   output        cfg_din3274,
   output        cfg_din3275,
   output        cfg_din3276,
   output        cfg_din3277,
   output        cfg_din3278,
   output        cfg_din3279,
   output        cfg_din3280,
   output        cfg_din3281,
   output        cfg_din3282,
   output        cfg_din3283,
   output        cfg_din3284,
   output        cfg_din3285,
   output        cfg_din3286,
   output        cfg_din3287,
   output        cfg_din3288,
   output        cfg_din3289,
   output        cfg_din3290,
   output        cfg_din3291,
   output        cfg_din3292,
   output        cfg_din3293,
   output        cfg_din3294,
   output        cfg_din3295,
   output        cfg_din3296,
   output        cfg_din3297,
   output        cfg_din3298,
   output        cfg_din3299,
   output        cfg_din3300,
   output        cfg_din3301,
   output        cfg_din3302,
   output        cfg_din3303,
   output        cfg_din3304,
   output        cfg_din3305,
   output        cfg_din3306,
   output        cfg_din3307,
   output        cfg_din3308,
   output        cfg_din3309,
   output        cfg_din3310,
   output        cfg_din3311,
   output        cfg_din3312,
   output        cfg_din3313,
   output        cfg_din3314,
   output        cfg_din3315,
   output        cfg_din3316,
   output        cfg_din3317,
   output        cfg_din3318,
   output        cfg_din3319,
   output        cfg_din3320,
   output        cfg_din3321,
   output        cfg_din3322,
   output        cfg_din3323,
   output        cfg_din3324,
   output        cfg_din3325,
   output        cfg_din3326,
   output        cfg_din3327,
   output        cfg_din3328,
   output        cfg_din3329,
   output        cfg_din3330,
   output        cfg_din3331,
   output        cfg_din3332,
   output        cfg_din3333,
   output        cfg_din3334,
   output        cfg_din3335,
   output        cfg_din3336,
   output        cfg_din3337,
   output        cfg_din3338,
   output        cfg_din3339,
   output        cfg_din3340,
   output        cfg_din3341,
   output        cfg_din3342,
   output        cfg_din3343,
   output        cfg_din3344,
   output        cfg_din3345,
   output        cfg_din3346,
   output        cfg_din3347,
   output        cfg_din3348,
   output        cfg_din3349,
   output        cfg_din3350,
   output        cfg_din3351,
   output        cfg_din3352,
   output        cfg_din3353,
   output        cfg_din3354,
   output        cfg_din3355,
   output        cfg_din3356,
   output        cfg_din3357,
   output        cfg_din3358,
   output        cfg_din3359,
   output        cfg_din3360,
   output        cfg_din3361,
   output        cfg_din3362,
   output        cfg_din3363,
   output        cfg_din3364,
   output        cfg_din3365,
   output        cfg_din3366,
   output        cfg_din3367,
   output        cfg_din3368,
   output        cfg_din3369,
   output        cfg_din3370,
   output        cfg_din3371,
   output        cfg_din3372,
   output        cfg_din3373,
   output        cfg_din3374,
   output        cfg_din3375,
   output        cfg_din3376,
   output        cfg_din3377,
   output        cfg_din3378,
   output        cfg_din3379,
   output        cfg_din3380,
   output        cfg_din3381,
   output        cfg_din3382,
   output        cfg_din3383,
   output        cfg_din3384,
   output        cfg_din3385,
   output        cfg_din3386,
   output        cfg_din3387,
   output        cfg_din3388,
   output        cfg_din3389,
   output        cfg_din3390,
   output        cfg_din3391,
   output        cfg_din3392,
   output        cfg_din3393,
   output        cfg_din3394,
   output        cfg_din3395,
   output        cfg_din3396,
   output        cfg_din3397,
   output        cfg_din3398,
   output        cfg_din3399,
   output        cfg_din3400,
   output        cfg_din3401,
   output        cfg_din3402,
   output        cfg_din3403,
   output        cfg_din3404,
   output        cfg_din3405,
   output        cfg_din3406,
   output        cfg_din3407,
   output        cfg_din3408,
   output        cfg_din3409,
   output        cfg_din3410,
   output        cfg_din3411,
   output        cfg_din3412,
   output        cfg_din3413,
   output        cfg_din3414,
   output        cfg_din3415,
   output        cfg_din3416,
   output        cfg_din3417,
   output        cfg_din3418,
   output        cfg_din3419,
   output        cfg_din3420,
   output        cfg_din3421,
   output        cfg_din3422,
   output        cfg_din3423,
   output        cfg_din3424,
   output        cfg_din3425,
   output        cfg_din3426,
   output        cfg_din3427,
   output        cfg_din3428,
   output        cfg_din3429,
   output        cfg_din3430,
   output        cfg_din3431,
   output        cfg_din3432,
   output        cfg_din3433,
   output        cfg_din3434,
   output        cfg_din3435,
   output        cfg_din3436,
   output        cfg_din3437,
   output        cfg_din3438,
   output        cfg_din3439,
   output        cfg_din3440,
   output        cfg_din3441,
   output        cfg_din3442,
   output        cfg_din3443,
   output        cfg_din3444,
   output        cfg_din3445,
   output        cfg_din3446,
   output        cfg_din3447,
   output        cfg_din3448,
   output        cfg_din3449,
   output        cfg_din3450,
   output        cfg_din3451,
   output        cfg_din3452,
   output        cfg_din3453,
   output        cfg_din3454,
   output        cfg_din3455,
   output        cfg_din3456,
   output        cfg_din3457,
   output        cfg_din3458,
   output        cfg_din3459,
   output        cfg_din3460,
   output        cfg_din3461,
   output        cfg_din3462,
   output        cfg_din3463,
   output        cfg_din3464,
   output        cfg_din3465,
   output        cfg_din3466,
   output        cfg_din3467,
   output        cfg_din3468,
   output        cfg_din3469,
   output        cfg_din3470,
   output        cfg_din3471,
   output        cfg_din3472,
   output        cfg_din3473,
   output        cfg_din3474,
   output        cfg_din3475,
   output        cfg_din3476,
   output        cfg_din3477,
   output        cfg_din3478,
   output        cfg_din3479,
   output        cfg_din3480,
   output        cfg_din3481,
   output        cfg_din3482,
   output        cfg_din3483,
   output        cfg_din3484,
   output        cfg_din3485,
   output        cfg_din3486,
   output        cfg_din3487,
   output        cfg_din3488,
   output        cfg_din3489,
   output        cfg_din3490,
   output        cfg_din3491,
   output        cfg_din3492,
   output        cfg_din3493,
   output        cfg_din3494,
   output        cfg_din3495,
   output        cfg_din3496,
   output        cfg_din3497,
   output        cfg_din3498,
   output        cfg_din3499,
   output        cfg_din3500,
   output        cfg_din3501,
   output        cfg_din3502,
   output        cfg_din3503,
   output        cfg_din3504,
   output        cfg_din3505,
   output        cfg_din3506,
   output        cfg_din3507,
   output        cfg_din3508,
   output        cfg_din3509,
   output        cfg_din3510,
   output        cfg_din3511,
   output        cfg_din3512,
   output        cfg_din3513,
   output        cfg_din3514,
   output        cfg_din3515,
   output        cfg_din3516,
   output        cfg_din3517,
   output        cfg_din3518,
   output        cfg_din3519,
   output        cfg_din3520,
   output        cfg_din3521,
   output        cfg_din3522,
   output        cfg_din3523,
   output        cfg_din3524,
   output        cfg_din3525,
   output        cfg_din3526,
   output        cfg_din3527,
   output        cfg_din3528,
   output        cfg_din3529,
   output        cfg_din3530,
   output        cfg_din3531,
   output        cfg_din3532,
   output        cfg_din3533,
   output        cfg_din3534,
   output        cfg_din3535,
   output        cfg_din3536,
   output        cfg_din3537,
   output        cfg_din3538,
   output        cfg_din3539,
   output        cfg_din3540,
   output        cfg_din3541,
   output        cfg_din3542,
   output        cfg_din3543,
   output        cfg_din3544,
   output        cfg_din3545,
   output        cfg_din3546,
   output        cfg_din3547,
   output        cfg_din3548,
   output        cfg_din3549,
   output        cfg_din3550,
   output        cfg_din3551,
   output        cfg_din3552,
   output        cfg_din3553,
   output        cfg_din3554,
   output        cfg_din3555,
   output        cfg_din3556,
   output        cfg_din3557,
   output        cfg_din3558,
   output        cfg_din3559,
   output        cfg_din3560,
   output        cfg_din3561,
   output        cfg_din3562,
   output        cfg_din3563,
   output        cfg_din3564,
   output        cfg_din3565,
   output        cfg_din3566,
   output        cfg_din3567,
   output        cfg_din3568,
   output        cfg_din3569,
   output        cfg_din3570,
   output        cfg_din3571,
   output        cfg_din3572,
   output        cfg_din3573,
   output        cfg_din3574,
   output        cfg_din3575,
   output        cfg_din3576,
   output        cfg_din3577,
   output        cfg_din3578,
   output        cfg_din3579,
   output        cfg_din3580,
   output        cfg_din3581,
   output        cfg_din3582,
   output        cfg_din3583,
   output        cfg_din3584,
   output        cfg_din3585,
   output        cfg_din3586,
   output        cfg_din3587,
   output        cfg_din3588,
   output        cfg_din3589,
   output        cfg_din3590,
   output        cfg_din3591,
   output        cfg_din3592,
   output        cfg_din3593,
   output        cfg_din3594,
   output        cfg_din3595,
   output        cfg_din3596,
   output        cfg_din3597,
   output        cfg_din3598,
   output        cfg_din3599,
   output        cfg_din3600,
   output        cfg_din3601,
   output        cfg_din3602,
   output        cfg_din3603,
   output        cfg_din3604,
   output        cfg_din3605,
   output        cfg_din3606,
   output        cfg_din3607,
   output        cfg_din3608,
   output        cfg_din3609,
   output        cfg_din3610,
   output        cfg_din3611,
   output        cfg_din3612,
   output        cfg_din3613,
   output        cfg_din3614,
   output        cfg_din3615,
   output        cfg_din3616,
   output        cfg_din3617,
   output        cfg_din3618,
   output        cfg_din3619,
   output        cfg_din3620,
   output        cfg_din3621,
   output        cfg_din3622,
   output        cfg_din3623,
   output        cfg_din3624,
   output        cfg_din3625,
   output        cfg_din3626,
   output        cfg_din3627,
   output        cfg_din3628,
   output        cfg_din3629,
   output        cfg_din3630,
   output        cfg_din3631,
   output        cfg_din3632,
   output        cfg_din3633,
   output        cfg_din3634,
   output        cfg_din3635,
   output        cfg_din3636,
   output        cfg_din3637,
   output        cfg_din3638,
   output        cfg_din3639,
   output        cfg_din3640,
   output        cfg_din3641,
   output        cfg_din3642,
   output        cfg_din3643,
   output        cfg_din3644,
   output        cfg_din3645,
   output        cfg_din3646,
   output        cfg_din3647,
   output        cfg_din3648,
   output        cfg_din3649,
   output        cfg_din3650,
   output        cfg_din3651,
   output        cfg_din3652,
   output        cfg_din3653,
   output        cfg_din3654,
   output        cfg_din3655,
   output        cfg_din3656,
   output        cfg_din3657,
   output        cfg_din3658,
   output        cfg_din3659,
   output        cfg_din3660,
   output        cfg_din3661,
   output        cfg_din3662,
   output        cfg_din3663,
   output        cfg_din3664,
   output        cfg_din3665,
   output        cfg_din3666,
   output        cfg_din3667,
   output        cfg_din3668,
   output        cfg_din3669,
   output        cfg_din3670,
   output        cfg_din3671,
   output        cfg_din3672,
   output        cfg_din3673,
   output        cfg_din3674,
   output        cfg_din3675,
   output        cfg_din3676,
   output        cfg_din3677,
   output        cfg_din3678,
   output        cfg_din3679,
   output        cfg_din3680,
   output        cfg_din3681,
   output        cfg_din3682,
   output        cfg_din3683,
   output        cfg_din3684,
   output        cfg_din3685,
   output        cfg_din3686,
   output        cfg_din3687,
   output        cfg_din3688,
   output        cfg_din3689,
   output        cfg_din3690,
   output        cfg_din3691,
   output        cfg_din3692,
   output        cfg_din3693,
   output        cfg_din3694,
   output        cfg_din3695,
   output        cfg_din3696,
   output        cfg_din3697,
   output        cfg_din3698,
   output        cfg_din3699,
   output        cfg_din3700,
   output        cfg_din3701,
   output        cfg_din3702,
   output        cfg_din3703,
   output        cfg_din3704,
   output        cfg_din3705,
   output        cfg_din3706,
   output        cfg_din3707,
   output        cfg_din3708,
   output        cfg_din3709,
   output        cfg_din3710,
   output        cfg_din3711,
   output        cfg_din3712,
   output        cfg_din3713,
   output        cfg_din3714,
   output        cfg_din3715,
   output        cfg_din3716,
   output        cfg_din3717,
   output        cfg_din3718,
   output        cfg_din3719,
   output        cfg_din3720,
   output        cfg_din3721,
   output        cfg_din3722,
   output        cfg_din3723,
   output        cfg_din3724,
   output        cfg_din3725,
   output        cfg_din3726,
   output        cfg_din3727,
   output        cfg_din3728,
   output        cfg_din3729,
   output        cfg_din3730,
   output        cfg_din3731,
   output        cfg_din3732,
   output        cfg_din3733,
   output        cfg_din3734,
   output        cfg_din3735,
   output        cfg_din3736,
   output        cfg_din3737,
   output        cfg_din3738,
   output        cfg_din3739,
   output        cfg_din3740,
   output        cfg_din3741,
   output        cfg_din3742,
   output        cfg_din3743,
   output        cfg_din3744,
   output        cfg_din3745,
   output        cfg_din3746,
   output        cfg_din3747,
   output        cfg_din3748,
   output        cfg_din3749,
   output        cfg_din3750,
   output        cfg_din3751,
   output        cfg_din3752,
   output        cfg_din3753,
   output        cfg_din3754,
   output        cfg_din3755,
   output        cfg_din3756,
   output        cfg_din3757,
   output        cfg_din3758,
   output        cfg_din3759,
   output        cfg_din3760,
   output        cfg_din3761,
   output        cfg_din3762,
   output        cfg_din3763,
   output        cfg_din3764,
   output        cfg_din3765,
   output        cfg_din3766,
   output        cfg_din3767,
   output        cfg_din3768,
   output        cfg_din3769,
   output        cfg_din3770,
   output        cfg_din3771,
   output        cfg_din3772,
   output        cfg_din3773,
   output        cfg_din3774,
   output        cfg_din3775,
   output        cfg_din3776,
   output        cfg_din3777,
   output        cfg_din3778,
   output        cfg_din3779,
   output        cfg_din3780,
   output        cfg_din3781,
   output        cfg_din3782,
   output        cfg_din3783,
   output        cfg_din3784,
   output        cfg_din3785,
   output        cfg_din3786,
   output        cfg_din3787,
   output        cfg_din3788,
   output        cfg_din3789,
   output        cfg_din3790,
   output        cfg_din3791,
   output        cfg_din3792,
   output        cfg_din3793,
   output        cfg_din3794,
   output        cfg_din3795,
   output        cfg_din3796,
   output        cfg_din3797,
   output        cfg_din3798,
   output        cfg_din3799,
   output        cfg_din3800,
   output        cfg_din3801,
   output        cfg_din3802,
   output        cfg_din3803,
   output        cfg_din3804,
   output        cfg_din3805,
   output        cfg_din3806,
   output        cfg_din3807,
   output        cfg_din3808,
   output        cfg_din3809,
   output        cfg_din3810,
   output        cfg_din3811,
   output        cfg_din3812,
   output        cfg_din3813,
   output        cfg_din3814,
   output        cfg_din3815,
   output        cfg_din3816,
   output        cfg_din3817,
   output        cfg_din3818,
   output        cfg_din3819,
   output        cfg_din3820,
   output        cfg_din3821,
   output        cfg_din3822,
   output        cfg_din3823,
   output        cfg_din3824,
   output        cfg_din3825,
   output        cfg_din3826,
   output        cfg_din3827,
   output        cfg_din3828,
   output        cfg_din3829,
   output        cfg_din3830,
   output        cfg_din3831,
   output        cfg_din3832,
   output        cfg_din3833,
   output        cfg_din3834,
   output        cfg_din3835,
   output        cfg_din3836,
   output        cfg_din3837,
   output        cfg_din3838,
   output        cfg_din3839,
   output        cfg_din3840,
   output        cfg_din3841,
   output        cfg_din3842,
   output        cfg_din3843,
   output        cfg_din3844,
   output        cfg_din3845,
   output        cfg_din3846,
   output        cfg_din3847,
   output        cfg_din3848,
   output        cfg_din3849,
   output        cfg_din3850,
   output        cfg_din3851,
   output        cfg_din3852,
   output        cfg_din3853,
   output        cfg_din3854,
   output        cfg_din3855,
   output        cfg_din3856,
   output        cfg_din3857,
   output        cfg_din3858,
   output        cfg_din3859,
   output        cfg_din3860,
   output        cfg_din3861,
   output        cfg_din3862,
   output        cfg_din3863,
   output        cfg_din3864,
   output        cfg_din3865,
   output        cfg_din3866,
   output        cfg_din3867,
   output        cfg_din3868,
   output        cfg_din3869,
   output        cfg_din3870,
   output        cfg_din3871,
   output        cfg_din3872,
   output        cfg_din3873,
   output        cfg_din3874,
   output        cfg_din3875,
   output        cfg_din3876,
   output        cfg_din3877,
   output        cfg_din3878,
   output        cfg_din3879,
   output        cfg_din3880,
   output        cfg_din3881,
   output        cfg_din3882,
   output        cfg_din3883,
   output        cfg_din3884,
   output        cfg_din3885,
   output        cfg_din3886,
   output        cfg_din3887,
   output        cfg_din3888,
   output        cfg_din3889,
   output        cfg_din3890,
   output        cfg_din3891,
   output        cfg_din3892,
   output        cfg_din3893,
   output        cfg_din3894,
   output        cfg_din3895,
   output        cfg_din3896,
   output        cfg_din3897,
   output        cfg_din3898,
   output        cfg_din3899,
   output        cfg_din3900,
   output        cfg_din3901,
   output        cfg_din3902,
   output        cfg_din3903,
   output        cfg_din3904,
   output        cfg_din3905,
   output        cfg_din3906,
   output        cfg_din3907,
   output        cfg_din3908,
   output        cfg_din3909,
   output        cfg_din3910,
   output        cfg_din3911,
   output        cfg_din3912,
   output        cfg_din3913,
   output        cfg_din3914,
   output        cfg_din3915,
   output        cfg_din3916,
   output        cfg_din3917,
   output        cfg_din3918,
   output        cfg_din3919,
   output        cfg_din3920,
   output        cfg_din3921,
   output        cfg_din3922,
   output        cfg_din3923,
   output        cfg_din3924,
   output        cfg_din3925,
   output        cfg_din3926,
   output        cfg_din3927,
   output        cfg_din3928,
   output        cfg_din3929,
   output        cfg_din3930,
   output        cfg_din3931,
   output        cfg_din3932,
   output        cfg_din3933,
   output        cfg_din3934,
   output        cfg_din3935,
   output        cfg_din3936,
   output        cfg_din3937,
   output        cfg_din3938,
   output        cfg_din3939,
   output        cfg_din3940,
   output        cfg_din3941,
   output        cfg_din3942,
   output        cfg_din3943,
   output        cfg_din3944,
   output        cfg_din3945,
   output        cfg_din3946,
   output        cfg_din3947,
   output        cfg_din3948,
   output        cfg_din3949,
   output        cfg_din3950,
   output        cfg_din3951,
   output        cfg_din3952,
   output        cfg_din3953,
   output        cfg_din3954,
   output        cfg_din3955,
   output        cfg_din3956,
   output        cfg_din3957,
   output        cfg_din3958,
   output        cfg_din3959,
   output        cfg_din3960,
   output        cfg_din3961,
   output        cfg_din3962,
   output        cfg_din3963,
   output        cfg_din3964,
   output        cfg_din3965,
   output        cfg_din3966,
   output        cfg_din3967,
   output        cfg_din3968,
   output        cfg_din3969,
   output        cfg_din3970,
   output        cfg_din3971,
   output        cfg_din3972,
   output        cfg_din3973,
   output        cfg_din3974,
   output        cfg_din3975,
   output        cfg_din3976,
   output        cfg_din3977,
   output        cfg_din3978,
   output        cfg_din3979,
   output        cfg_din3980,
   output        cfg_din3981,
   output        cfg_din3982,
   output        cfg_din3983,
   output        cfg_din3984,
   output        cfg_din3985,
   output        cfg_din3986,
   output        cfg_din3987,
   output        cfg_din3988,
   output        cfg_din3989,
   output        cfg_din3990,
   output        cfg_din3991,
   output        cfg_din3992,
   output        cfg_din3993,
   output        cfg_din3994,
   output        cfg_din3995,
   output        cfg_din3996,
   output        cfg_din3997,
   output        cfg_din3998,
   output        cfg_din3999,
   output        cfg_din4000,
   output        cfg_din4001,
   output        cfg_din4002,
   output        cfg_din4003,
   output        cfg_din4004,
   output        cfg_din4005,
   output        cfg_din4006,
   output        cfg_din4007,
   output        cfg_din4008,
   output        cfg_din4009,
   output        cfg_din4010,
   output        cfg_din4011,
   output        cfg_din4012,
   output        cfg_din4013,
   output        cfg_din4014,
   output        cfg_din4015,
   output        cfg_din4016,
   output        cfg_din4017,
   output        cfg_din4018,
   output        cfg_din4019,
   output        cfg_din4020,
   output        cfg_din4021,
   output        cfg_din4022,
   output        cfg_din4023,
   output        cfg_din4024,
   output        cfg_din4025,
   output        cfg_din4026,
   output        cfg_din4027,
   output        cfg_din4028,
   output        cfg_din4029,
   output        cfg_din4030,
   output        cfg_din4031,
   output        cfg_din4032,
   output        cfg_din4033,
   output        cfg_din4034,
   output        cfg_din4035,
   output        cfg_din4036,
   output        cfg_din4037,
   output        cfg_din4038,
   output        cfg_din4039,
   output        cfg_din4040,
   output        cfg_din4041,
   output        cfg_din4042,
   output        cfg_din4043,
   output        cfg_din4044,
   output        cfg_din4045,
   output        cfg_din4046,
   output        cfg_din4047,
   output        cfg_din4048,
   output        cfg_din4049,
   output        cfg_din4050,
   output        cfg_din4051,
   output        cfg_din4052,
   output        cfg_din4053,
   output        cfg_din4054,
   output        cfg_din4055,
   output        cfg_din4056,
   output        cfg_din4057,
   output        cfg_din4058,
   output        cfg_din4059,
   output        cfg_din4060,
   output        cfg_din4061,
   output        cfg_din4062,
   output        cfg_din4063,
   output        cfg_din4064,
   output        cfg_din4065,
   output        cfg_din4066,
   output        cfg_din4067,
   output        cfg_din4068,
   output        cfg_din4069,
   output        cfg_din4070,
   output        cfg_din4071,
   output        cfg_din4072,
   output        cfg_din4073,
   output        cfg_din4074,
   output        cfg_din4075,
   output        cfg_din4076,
   output        cfg_din4077,
   output        cfg_din4078,
   output        cfg_din4079,
   output        cfg_din4080,
   output        cfg_din4081,
   output        cfg_din4082,
   output        cfg_din4083,
   output        cfg_din4084,
   output        cfg_din4085,
   output        cfg_din4086,
   output        cfg_din4087,
   output        cfg_din4088,
   output        cfg_din4089,
   output        cfg_din4090,
   output        cfg_din4091,
   output        cfg_din4092,
   output        cfg_din4093,
   output        cfg_din4094,
   output        cfg_din4095,
   output        cfg_din4096,
   output        cfg_din4097,
   output        cfg_din4098,
   output        cfg_din4099,
   output        cfg_din4100,
   output        cfg_din4101,
   output        cfg_din4102,
   output        cfg_din4103,
   output        cfg_din4104,
   output        cfg_din4105,
   output        cfg_din4106,
   output        cfg_din4107,
   output        cfg_din4108,
   output        cfg_din4109,
   output        cfg_din4110,
   output        cfg_din4111,
   output        cfg_din4112,
   output        cfg_din4113,
   output        cfg_din4114,
   output        cfg_din4115,
   output        cfg_din4116,
   output        cfg_din4117,
   output        cfg_din4118,
   output        cfg_din4119,
   output        cfg_din4120,
   output        cfg_din4121,
   output        cfg_din4122,
   output        cfg_din4123,
   output        cfg_din4124,
   output        cfg_din4125,
   output        cfg_din4126,
   output        cfg_din4127,
   output        cfg_din4128,
   output        cfg_din4129,
   output        cfg_din4130,
   output        cfg_din4131,
   output        cfg_din4132,
   output        cfg_din4133,
   output        cfg_din4134,
   output        cfg_din4135,
   output        cfg_din4136,
   output        cfg_din4137,
   output        cfg_din4138,
   output        cfg_din4139,
   output        cfg_din4140,
   output        cfg_din4141,
   output        cfg_din4142,
   output        cfg_din4143,
   output        cfg_din4144,
   output        cfg_din4145,
   output        cfg_din4146,
   output        cfg_din4147,
   output        cfg_din4148,
   output        cfg_din4149,
   output        cfg_din4150,
   output        cfg_din4151,
   output        cfg_din4152,
   output        cfg_din4153,
   output        cfg_din4154,
   output        cfg_din4155,
   output        cfg_din4156,
   output        cfg_din4157,
   output        cfg_din4158,
   output        cfg_din4159,
   output        cfg_din4160,
   output        cfg_din4161,
   output        cfg_din4162,
   output        cfg_din4163,
   output        cfg_din4164,
   output        cfg_din4165,
   output        cfg_din4166,
   output        cfg_din4167,
   output        cfg_din4168,
   output        cfg_din4169,
   output        cfg_din4170,
   output        cfg_din4171,
   output        cfg_din4172,
   output        cfg_din4173,
   output        cfg_din4174,
   output        cfg_din4175,
   output        cfg_din4176,
   output        cfg_din4177,
   output        cfg_din4178,
   output        cfg_din4179,
   output        cfg_din4180,
   output        cfg_din4181,
   output        cfg_din4182,
   output        cfg_din4183,
   output        cfg_din4184,
   output        cfg_din4185,
   output        cfg_din4186,
   output        cfg_din4187,
   output        cfg_din4188,
   output        cfg_din4189,
   output        cfg_din4190,
   output        cfg_din4191,
   output        cfg_din4192,
   output        cfg_din4193,
   output        cfg_din4194,
   output        cfg_din4195,
   output        cfg_din4196,
   output        cfg_din4197,
   output        cfg_din4198,
   output        cfg_din4199,
   output        cfg_din4200,
   output        cfg_din4201,
   output        cfg_din4202,
   output        cfg_din4203,
   output        cfg_din4204,
   output        cfg_din4205,
   output        cfg_din4206,
   output        cfg_din4207,
   output        cfg_din4208,
   output        cfg_din4209,
   output        cfg_din4210,
   output        cfg_din4211,
   output        cfg_din4212,
   output        cfg_din4213,
   output        cfg_din4214,
   output        cfg_din4215,
   output        cfg_din4216,
   output        cfg_din4217,
   output        cfg_din4218,
   output        cfg_din4219,
   output        cfg_din4220,
   output        cfg_din4221,
   output        cfg_din4222,
   output        cfg_din4223,
   output        cfg_din4224,
   output        cfg_din4225,
   output        cfg_din4226,
   output        cfg_din4227,
   output        cfg_din4228,
   output        cfg_din4229,
   output        cfg_din4230,
   output        cfg_din4231,
   output        cfg_din4232,
   output        cfg_din4233,
   output        cfg_din4234,
   output        cfg_din4235,
   output        cfg_din4236,
   output        cfg_din4237,
   output        cfg_din4238,
   output        cfg_din4239,
   output        cfg_din4240,
   output        cfg_din4241,
   output        cfg_din4242,
   output        cfg_din4243,
   output        cfg_din4244,
   output        cfg_din4245,
   output        cfg_din4246,
   output        cfg_din4247,
   output        cfg_din4248,
   output        cfg_din4249,
   output        cfg_din4250,
   output        cfg_din4251,
   output        cfg_din4252,
   output        cfg_din4253,
   output        cfg_din4254,
   output        cfg_din4255,
   output        cfg_din4256,
   output        cfg_din4257,
   output        cfg_din4258,
   output        cfg_din4259,
   output        cfg_din4260,
   output        cfg_din4261,
   output        cfg_din4262,
   output        cfg_din4263,
   output        cfg_din4264,
   output        cfg_din4265,
   output        cfg_din4266,
   output        cfg_din4267,
   output        cfg_din4268,
   output        cfg_din4269,
   output        cfg_din4270,
   output        cfg_din4271,
   output        cfg_din4272,
   output        cfg_din4273,
   output        cfg_din4274,
   output        cfg_din4275,
   output        cfg_din4276,
   output        cfg_din4277,
   output        cfg_din4278,
   output        cfg_din4279,
   output        cfg_din4280,
   output        cfg_din4281,
   output        cfg_din4282,
   output        cfg_din4283,
   output        cfg_din4284,
   output        cfg_din4285,
   output        cfg_din4286,
   output        cfg_din4287,
   output        cfg_din4288,
   output        cfg_din4289,
   output        cfg_din4290,
   output        cfg_din4291,
   output        cfg_din4292,
   output        cfg_din4293,
   output        cfg_din4294,
   output        cfg_din4295,
   output        cfg_din4296,
   output        cfg_din4297,
   output        cfg_din4298,
   output        cfg_din4299,
   output        cfg_din4300,
   output        cfg_din4301,
   output        cfg_din4302,
   output        cfg_din4303,
   output        cfg_din4304,
   output        cfg_din4305,
   output        cfg_din4306,
   output        cfg_din4307,
   output        cfg_din4308,
   output        cfg_din4309,
   output        cfg_din4310,
   output        cfg_din4311,
   output        cfg_din4312,
   output        cfg_din4313,
   output        cfg_din4314,
   output        cfg_din4315,
   output        cfg_din4316,
   output        cfg_din4317,
   output        cfg_din4318,
   output        cfg_din4319,
   output        cfg_din4320,
   output        cfg_din4321,
   output        cfg_din4322,
   output        cfg_din4323,
   output        cfg_din4324,
   output        cfg_din4325,
   output        cfg_din4326,
   output        cfg_din4327,
   output        cfg_din4328,
   output        cfg_din4329,
   output        cfg_din4330,
   output        cfg_din4331,
   output        cfg_din4332,
   output        cfg_din4333,
   output        cfg_din4334,
   output        cfg_din4335,
   output        cfg_din4336,
   output        cfg_din4337,
   output        cfg_din4338,
   output        cfg_din4339,
   output        cfg_din4340,
   output        cfg_din4341,
   output        cfg_din4342,
   output        cfg_din4343,
   output        cfg_din4344,
   output        cfg_din4345,
   output        cfg_din4346,
   output        cfg_din4347,
   output        cfg_din4348,
   output        cfg_din4349,
   output        cfg_din4350,
   output        cfg_din4351,
   output        cfg_din4352,
   output        cfg_din4353,
   output        cfg_din4354,
   output        cfg_din4355,
   output        cfg_din4356,
   output        cfg_din4357,
   output        cfg_din4358,
   output        cfg_din4359,
   output        cfg_din4360,
   output        cfg_din4361,
   output        cfg_din4362,
   output        cfg_din4363,
   output        cfg_din4364,
   output        cfg_din4365,
   output        cfg_din4366,
   output        cfg_din4367,
   output        cfg_din4368,
   output        cfg_din4369,
   output        cfg_din4370,
   output        cfg_din4371,
   output        cfg_din4372,
   output        cfg_din4373,
   output        cfg_din4374,
   output        cfg_din4375,
   output        cfg_din4376,
   output        cfg_din4377,
   output        cfg_din4378,
   output        cfg_din4379,
   output        cfg_din4380,
   output        cfg_din4381,
   output        cfg_din4382,
   output        cfg_din4383,
   output        cfg_din4384,
   output        cfg_din4385,
   output        cfg_din4386,
   output        cfg_din4387,
   output        cfg_din4388,
   output        cfg_din4389,
   output        cfg_din4390,
   output        cfg_din4391,
   output        cfg_din4392,
   output        cfg_din4393,
   output        cfg_din4394,
   output        cfg_din4395,
   output        cfg_din4396,
   output        cfg_din4397,
   output        cfg_din4398,
   output        cfg_din4399,
   output        cfg_din4400,
   output        cfg_din4401,
   output        cfg_din4402,
   output        cfg_din4403,
   output        cfg_din4404,
   output        cfg_din4405,
   output        cfg_din4406,
   output        cfg_din4407,
   output        cfg_din4408,
   output        cfg_din4409,
   output        cfg_din4410,
   output        cfg_din4411,
   output        cfg_din4412,
   output        cfg_din4413,
   output        cfg_din4414,
   output        cfg_din4415,
   output        cfg_din4416,
   output        cfg_din4417,
   output        cfg_din4418,
   output        cfg_din4419,
   output        cfg_din4420,
   output        cfg_din4421,
   output        cfg_din4422,
   output        cfg_din4423,
   output        cfg_din4424,
   output        cfg_din4425,
   output        cfg_din4426,
   output        cfg_din4427,
   output        cfg_din4428,
   output        cfg_din4429,
   output        cfg_din4430,
   output        cfg_din4431,
   output        cfg_din4432,
   output        cfg_din4433,
   output        cfg_din4434,
   output        cfg_din4435,
   output        cfg_din4436,
   output        cfg_din4437,
   output        cfg_din4438,
   output        cfg_din4439,
   output        cfg_din4440,
   output        cfg_din4441,
   output        cfg_din4442,
   output        cfg_din4443,
   output        cfg_din4444,
   output        cfg_din4445,
   output        cfg_din4446,
   output        cfg_din4447,
   output        cfg_din4448,
   output        cfg_din4449,
   output        cfg_din4450,
   output        cfg_din4451,
   output        cfg_din4452,
   output        cfg_din4453,
   output        cfg_din4454,
   output        cfg_din4455,
   output        cfg_din4456,
   output        cfg_din4457,
   output        cfg_din4458,
   output        cfg_din4459,
   output        cfg_din4460,
   output        cfg_din4461,
   output        cfg_din4462,
   output        cfg_din4463,
   output        cfg_din4464,
   output        cfg_din4465,
   output        cfg_din4466,
   output        cfg_din4467,
   output        cfg_din4468,
   output        cfg_din4469,
   output        cfg_din4470,
   output        cfg_din4471,
   output        cfg_din4472,
   output        cfg_din4473,
   output        cfg_din4474,
   output        cfg_din4475,
   output        cfg_din4476,
   output        cfg_din4477,
   output        cfg_din4478,
   output        cfg_din4479,
   output        cfg_din4480,
   output        cfg_din4481,
   output        cfg_din4482,
   output        cfg_din4483,
   output        cfg_din4484,
   output        cfg_din4485,
   output        cfg_din4486,
   output        cfg_din4487,
   output        cfg_din4488,
   output        cfg_din4489,
   output        cfg_din4490,
   output        cfg_din4491,
   output        cfg_din4492,
   output        cfg_din4493,
   output        cfg_din4494,
   output        cfg_din4495,
   output        cfg_din4496,
   output        cfg_din4497,
   output        cfg_din4498,
   output        cfg_din4499,
   output        cfg_din4500,
   output        cfg_din4501,
   output        cfg_din4502,
   output        cfg_din4503,
   output        cfg_din4504,
   output        cfg_din4505,
   output        cfg_din4506,
   output        cfg_din4507,
   output        cfg_din4508,
   output        cfg_din4509,
   output        cfg_din4510,
   output        cfg_din4511,
   output        cfg_din4512,
   output        cfg_din4513,
   output        cfg_din4514,
   output        cfg_din4515,
   output        cfg_din4516,
   output        cfg_din4517,
   output        cfg_din4518,
   output        cfg_din4519,
   output        cfg_din4520,
   output        cfg_din4521,
   output        cfg_din4522,
   output        cfg_din4523,
   output        cfg_din4524,
   output        cfg_din4525,
   output        cfg_din4526,
   output        cfg_din4527,
   output        cfg_din4528,
   output        cfg_din4529,
   output        cfg_din4530,
   output        cfg_din4531,
   output        cfg_din4532,
   output        cfg_din4533,
   output        cfg_din4534,
   output        cfg_din4535,
   output        cfg_din4536,
   output        cfg_din4537,
   output        cfg_din4538,
   output        cfg_din4539,
   output        cfg_din4540,
   output        cfg_din4541,
   output        cfg_din4542,
   output        cfg_din4543,
   output        cfg_din4544,
   output        cfg_din4545,
   output        cfg_din4546,
   output        cfg_din4547,
   output        cfg_din4548,
   output        cfg_din4549,
   output        cfg_din4550,
   output        cfg_din4551,
   output        cfg_din4552,
   output        cfg_din4553,
   output        cfg_din4554,
   output        cfg_din4555,
   output        cfg_din4556,
   output        cfg_din4557,
   output        cfg_din4558,
   output        cfg_din4559,
   output        cfg_din4560,
   output        cfg_din4561,
   output        cfg_din4562,
   output        cfg_din4563,
   output        cfg_din4564,
   output        cfg_din4565,
   output        cfg_din4566,
   output        cfg_din4567,
   output        cfg_din4568,
   output        cfg_din4569,
   output        cfg_din4570,
   output        cfg_din4571,
   output        cfg_din4572,
   output        cfg_din4573,
   output        cfg_din4574,
   output        cfg_din4575,
   output        cfg_din4576,
   output        cfg_din4577,
   output        cfg_din4578,
   output        cfg_din4579,
   output        cfg_din4580,
   output        cfg_din4581,
   output        cfg_din4582,
   output        cfg_din4583,
   output        cfg_din4584,
   output        cfg_din4585,
   output        cfg_din4586,
   output        cfg_din4587,
   output        cfg_din4588,
   output        cfg_din4589,
   output        cfg_din4590,
   output        cfg_din4591,
   output        cfg_din4592,
   output        cfg_din4593,
   output        cfg_din4594,
   output        cfg_din4595,
   output        cfg_din4596,
   output        cfg_din4597,
   output        cfg_din4598,
   output        cfg_din4599,
   output        cfg_din4600,
   output        cfg_din4601,
   output        cfg_din4602,
   output        cfg_din4603,
   output        cfg_din4604,
   output        cfg_din4605,
   output        cfg_din4606,
   output        cfg_din4607,
   output        cfg_din4608,
   output        cfg_din4609,
   output        cfg_din4610,
   output        cfg_din4611,
   output        cfg_din4612,
   output        cfg_din4613,
   output        cfg_din4614,
   output        cfg_din4615,
   output        cfg_din4616,
   output        cfg_din4617,
   output        cfg_din4618,
   output        cfg_din4619,
   output        cfg_din4620,
   output        cfg_din4621,
   output        cfg_din4622,
   output        cfg_din4623,
   output        cfg_din4624,
   output        cfg_din4625,
   output        cfg_din4626,
   output        cfg_din4627,
   output        cfg_din4628,
   output        cfg_din4629,
   output        cfg_din4630,
   output        cfg_din4631,
   output        cfg_din4632,
   output        cfg_din4633,
   output        cfg_din4634,
   output        cfg_din4635,
   output        cfg_din4636,
   output        cfg_din4637,
   output        cfg_din4638,
   output        cfg_din4639,
   output        cfg_din4640,
   output        cfg_din4641,
   output        cfg_din4642,
   output        cfg_din4643,
   output        cfg_din4644,
   output        cfg_din4645,
   output        cfg_din4646,
   output        cfg_din4647,
   output        cfg_din4648,
   output        cfg_din4649,
   output        cfg_din4650,
   output        cfg_din4651,
   output        cfg_din4652,
   output        cfg_din4653,
   output        cfg_din4654,
   output        cfg_din4655,
   output        cfg_din4656,
   output        cfg_din4657,
   output        cfg_din4658,
   output        cfg_din4659,
   output        cfg_din4660,
   output        cfg_din4661,
   output        cfg_din4662,
   output        cfg_din4663,
   output        cfg_din4664,
   output        cfg_din4665,
   output        cfg_din4666,
   output        cfg_din4667,
   output        cfg_din4668,
   output        cfg_din4669,
   output        cfg_din4670,
   output        cfg_din4671,
   output        cfg_din4672,
   output        cfg_din4673,
   output        cfg_din4674,
   output        cfg_din4675,
   output        cfg_din4676,
   output        cfg_din4677,
   output        cfg_din4678,
   output        cfg_din4679,
   output        cfg_din4680,
   output        cfg_din4681,
   output        cfg_din4682,
   output        cfg_din4683,
   output        cfg_din4684,
   output        cfg_din4685,
   output        cfg_din4686,
   output        cfg_din4687,
   output        cfg_din4688,
   output        cfg_din4689,
   output        cfg_din4690,
   output        cfg_din4691,
   output        cfg_din4692,
   output        cfg_din4693,
   output        cfg_din4694,
   output        cfg_din4695,
   output        cfg_din4696,
   output        cfg_din4697,
   output        cfg_din4698,
   output        cfg_din4699,
   output        cfg_din4700,
   output        cfg_din4701,
   output        cfg_din4702,
   output        cfg_din4703,
   output        cfg_din4704,
   output        cfg_din4705,
   output        cfg_din4706,
   output        cfg_din4707,
   output        cfg_din4708,
   output        cfg_din4709,
   output        cfg_din4710,
   output        cfg_din4711,
   output        cfg_din4712,
   output        cfg_din4713,
   output        cfg_din4714,
   output        cfg_din4715,
   output        cfg_din4716,
   output        cfg_din4717,
   output        cfg_din4718,
   output        cfg_din4719,
   output        cfg_din4720,
   output        cfg_din4721,
   output        cfg_din4722,
   output        cfg_din4723,
   output        cfg_din4724,
   output        cfg_din4725,
   output        cfg_din4726,
   output        cfg_din4727,
   output        cfg_din4728,
   output        cfg_din4729,
   output        cfg_din4730,
   output        cfg_din4731,
   output        cfg_din4732,
   output        cfg_din4733,
   output        cfg_din4734,
   output        cfg_din4735,
   output        cfg_din4736,
   output        cfg_din4737,
   output        cfg_din4738,
   output        cfg_din4739,
   output        cfg_din4740,
   output        cfg_din4741,
   output        cfg_din4742,
   output        cfg_din4743,
   output        cfg_din4744,
   output        cfg_din4745,
   output        cfg_din4746,
   output        cfg_din4747,
   output        cfg_din4748,
   output        cfg_din4749,
   output        cfg_din4750,
   output        cfg_din4751,
   output        cfg_din4752,
   output        cfg_din4753,
   output        cfg_din4754,
   output        cfg_din4755,
   output        cfg_din4756,
   output        cfg_din4757,
   output        cfg_din4758,
   output        cfg_din4759,
   output        cfg_din4760,
   output        cfg_din4761,
   output        cfg_din4762,
   output        cfg_din4763,
   output        cfg_din4764,
   output        cfg_din4765,
   output        cfg_din4766,
   output        cfg_din4767,
   output        cfg_din4768,
   output        cfg_din4769,
   output        cfg_din4770,
   output        cfg_din4771,
   output        cfg_din4772,
   output        cfg_din4773,
   output        cfg_din4774,
   output        cfg_din4775,
   output        cfg_din4776,
   output        cfg_din4777,
   output        cfg_din4778,
   output        cfg_din4779,
   output        cfg_din4780,
   output        cfg_din4781,
   output        cfg_din4782,
   output        cfg_din4783,
   output        cfg_din4784,
   output        cfg_din4785,
   output        cfg_din4786,
   output        cfg_din4787,
   output        cfg_din4788,
   output        cfg_din4789,
   output        cfg_din4790,
   output        cfg_din4791,
   output        cfg_din4792,
   output        cfg_din4793,
   output        cfg_din4794,
   output        cfg_din4795,
   output        cfg_din4796,
   output        cfg_din4797,
   output        cfg_din4798,
   output        cfg_din4799,
   output        cfg_din4800,
   output        cfg_din4801,
   output        cfg_din4802,
   output        cfg_din4803,
   output        cfg_din4804,
   output        cfg_din4805,
   output        cfg_din4806,
   output        cfg_din4807,
   output        cfg_din4808,
   output        cfg_din4809,
   output        cfg_din4810,
   output        cfg_din4811,
   output        cfg_din4812,
   output        cfg_din4813,
   output        cfg_din4814,
   output        cfg_din4815,
   output        cfg_din4816,
   output        cfg_din4817,
   output        cfg_din4818,
   output        cfg_din4819,
   output        cfg_din4820,
   output        cfg_din4821,
   output        cfg_din4822,
   output        cfg_din4823,
   output        cfg_din4824,
   output        cfg_din4825,
   output        cfg_din4826,
   output        cfg_din4827,
   output        cfg_din4828,
   output        cfg_din4829,
   output        cfg_din4830,
   output        cfg_din4831,
   output        cfg_din4832,
   output        cfg_din4833,
   output        cfg_din4834,
   output        cfg_din4835,
   output        cfg_din4836,
   output        cfg_din4837,
   output        cfg_din4838,
   output        cfg_din4839,
   output        cfg_din4840,
   output        cfg_din4841,
   output        cfg_din4842,
   output        cfg_din4843,
   output        cfg_din4844,
   output        cfg_din4845,
   output        cfg_din4846,
   output        cfg_din4847,
   output        cfg_din4848,
   output        cfg_din4849,
   output        cfg_din4850,
   output        cfg_din4851,
   output        cfg_din4852,
   output        cfg_din4853,
   output        cfg_din4854,
   output        cfg_din4855,
   output        cfg_din4856,
   output        cfg_din4857,
   output        cfg_din4858,
   output        cfg_din4859,
   output        cfg_din4860,
   output        cfg_din4861,
   output        cfg_din4862,
   output        cfg_din4863,
   output        cfg_din4864,
   output        cfg_din4865,
   output        cfg_din4866,
   output        cfg_din4867,
   output        cfg_din4868,
   output        cfg_din4869,
   output        cfg_din4870,
   output        cfg_din4871,
   output        cfg_din4872,
   output        cfg_din4873,
   output        cfg_din4874,
   output        cfg_din4875,
   output        cfg_din4876,
   output        cfg_din4877,
   output        cfg_din4878,
   output        cfg_din4879,
   output        cfg_din4880,
   output        cfg_din4881,
   output        cfg_din4882,
   output        cfg_din4883,
   output        cfg_din4884,
   output        cfg_din4885,
   output        cfg_din4886,
   output        cfg_din4887,
   output        cfg_din4888,
   output        cfg_din4889,
   output        cfg_din4890,
   output        cfg_din4891,
   output        cfg_din4892,
   output        cfg_din4893,
   output        cfg_din4894,
   output        cfg_din4895,
   output        cfg_din4896,
   output        cfg_din4897,
   output        cfg_din4898,
   output        cfg_din4899,
   output        cfg_din4900,
   output        cfg_din4901,
   output        cfg_din4902,
   output        cfg_din4903,
   output        cfg_din4904,
   output        cfg_din4905,
   output        cfg_din4906,
   output        cfg_din4907,
   output        cfg_din4908,
   output        cfg_din4909,
   output        cfg_din4910,
   output        cfg_din4911,
   output        cfg_din4912,
   output        cfg_din4913,
   output        cfg_din4914,
   output        cfg_din4915,
   output        cfg_din4916,
   output        cfg_din4917,
   output        cfg_din4918,
   output        cfg_din4919,
   output        cfg_din4920,
   output        cfg_din4921,
   output        cfg_din4922,
   output        cfg_din4923,
   output        cfg_din4924,
   output        cfg_din4925,
   output        cfg_din4926,
   output        cfg_din4927,
   output        cfg_din4928,
   output        cfg_din4929,
   output        cfg_din4930,
   output        cfg_din4931,
   output        cfg_din4932,
   output        cfg_din4933,
   output        cfg_din4934,
   output        cfg_din4935,
   output        cfg_din4936,
   output        cfg_din4937,
   output        cfg_din4938,
   output        cfg_din4939,
   output        cfg_din4940,
   output        cfg_din4941,
   output        cfg_din4942,
   output        cfg_din4943,
   output        cfg_din4944,
   output        cfg_din4945,
   output        cfg_din4946,
   output        cfg_din4947,
   output        cfg_din4948,
   output        cfg_din4949,
   output        cfg_din4950,
   output        cfg_din4951,
   output        cfg_din4952,
   output        cfg_din4953,
   output        cfg_din4954,
   output        cfg_din4955,
   output        cfg_din4956,
   output        cfg_din4957,
   output        cfg_din4958,
   output        cfg_din4959,
   output        cfg_din4960,
   output        cfg_din4961,
   output        cfg_din4962,
   output        cfg_din4963,
   output        cfg_din4964,
   output        cfg_din4965,
   output        cfg_din4966,
   output        cfg_din4967,
   output        cfg_din4968,
   output        cfg_din4969,
   output        cfg_din4970,
   output        cfg_din4971,
   output        cfg_din4972,
   output        cfg_din4973,
   output        cfg_din4974,
   output        cfg_din4975,
   output        cfg_din4976,
   output        cfg_din4977,
   output        cfg_din4978,
   output        cfg_din4979,
   output        cfg_din4980,
   output        cfg_din4981,
   output        cfg_din4982,
   output        cfg_din4983,
   output        cfg_din4984,
   output        cfg_din4985,
   output        cfg_din4986,
   output        cfg_din4987,
   output        cfg_din4988,
   output        cfg_din4989,
   output        cfg_din4990,
   output        cfg_din4991,
   output        cfg_din4992,
   output        cfg_din4993,
   output        cfg_din4994,
   output        cfg_din4995,
   output        cfg_din4996,
   output        cfg_din4997,
   output        cfg_din4998,
   output        cfg_din4999,
   output        cfg_din5000,
   output        cfg_din5001,
   output        cfg_din5002,
   output        cfg_din5003,
   output        cfg_din5004,
   output        cfg_din5005,
   output        cfg_din5006,
   output        cfg_din5007,
   output        cfg_din5008,
   output        cfg_din5009,
   output        cfg_din5010,
   output        cfg_din5011,
   output        cfg_din5012,
   output        cfg_din5013,
   output        cfg_din5014,
   output        cfg_din5015,
   output        cfg_din5016,
   output        cfg_din5017,
   output        cfg_din5018,
   output        cfg_din5019,
   output        cfg_din5020,
   output        cfg_din5021,
   output        cfg_din5022,
   output        cfg_din5023,
   output        cfg_din5024,
   output        cfg_din5025,
   output        cfg_din5026,
   output        cfg_din5027,
   output        cfg_din5028,
   output        cfg_din5029,
   output        cfg_din5030,
   output        cfg_din5031,
   output        cfg_din5032,
   output        cfg_din5033,
   output        cfg_din5034,
   output        cfg_din5035,
   output        cfg_din5036,
   output        cfg_din5037,
   output        cfg_din5038,
   output        cfg_din5039,
   output        cfg_din5040,
   output        cfg_din5041,
   output        cfg_din5042,
   output        cfg_din5043,
   output        cfg_din5044,
   output        cfg_din5045,
   output        cfg_din5046,
   output        cfg_din5047,
   output        cfg_din5048,
   output        cfg_din5049,
   output        cfg_din5050,
   output        cfg_din5051,
   output        cfg_din5052,
   output        cfg_din5053,
   output        cfg_din5054,
   output        cfg_din5055,
   output        cfg_din5056,
   output        cfg_din5057,
   output        cfg_din5058,
   output        cfg_din5059,
   output        cfg_din5060,
   output        cfg_din5061,
   output        cfg_din5062,
   output        cfg_din5063,
   output        cfg_din5064,
   output        cfg_din5065,
   output        cfg_din5066,
   output        cfg_din5067,
   output        cfg_din5068,
   output        cfg_din5069,
   output        cfg_din5070,
   output        cfg_din5071,
   output        cfg_din5072,
   output        cfg_din5073,
   output        cfg_din5074,
   output        cfg_din5075,
   output        cfg_din5076,
   output        cfg_din5077,
   output        cfg_din5078,
   output        cfg_din5079,
   output        cfg_din5080,
   output        cfg_din5081,
   output        cfg_din5082,
   output        cfg_din5083,
   output        cfg_din5084,
   output        cfg_din5085,
   output        cfg_din5086,
   output        cfg_din5087,
   output        cfg_din5088,
   output        cfg_din5089,
   output        cfg_din5090,
   output        cfg_din5091,
   output        cfg_din5092,
   output        cfg_din5093,
   output        cfg_din5094,
   output        cfg_din5095,
   output        cfg_din5096,
   output        cfg_din5097,
   output        cfg_din5098,
   output        cfg_din5099,
   output        cfg_din5100,
   output        cfg_din5101,
   output        cfg_din5102,
   output        cfg_din5103,
   output        cfg_din5104,
   output        cfg_din5105,
   output        cfg_din5106,
   output        cfg_din5107,
   output        cfg_din5108,
   output        cfg_din5109,
   output        cfg_din5110,
   output        cfg_din5111,
   output        cfg_din5112,
   output        cfg_din5113,
   output        cfg_din5114,
   output        cfg_din5115,
   output        cfg_din5116,
   output        cfg_din5117,
   output        cfg_din5118,
   output        cfg_din5119,
   output        cfg_din5120,
   output        cfg_din5121,
   output        cfg_din5122,
   output        cfg_din5123,
   output        cfg_din5124,
   output        cfg_din5125,
   output        cfg_din5126,
   output        cfg_din5127,
   output        cfg_din5128,
   output        cfg_din5129,
   output        cfg_din5130,
   output        cfg_din5131,
   output        cfg_din5132,
   output        cfg_din5133,
   output        cfg_din5134,
   output        cfg_din5135,
   output        cfg_din5136,
   output        cfg_din5137,
   output        cfg_din5138,
   output        cfg_din5139,
   output        cfg_din5140,
   output        cfg_din5141,
   output        cfg_din5142,
   output        cfg_din5143,
   output        cfg_din5144,
   output        cfg_din5145,
   output        cfg_din5146,
   output        cfg_din5147,
   output        cfg_din5148,
   output        cfg_din5149,
   output        cfg_din5150,
   output        cfg_din5151,
   output        cfg_din5152,
   output        cfg_din5153,
   output        cfg_din5154,
   output        cfg_din5155,
   output        cfg_din5156,
   output        cfg_din5157,
   output        cfg_din5158,
   output        cfg_din5159,
   output        cfg_din5160,
   output        cfg_din5161,
   output        cfg_din5162,
   output        cfg_din5163,
   output        cfg_din5164,
   output        cfg_din5165,
   output        cfg_din5166,
   output        cfg_din5167,
   output        cfg_din5168,
   output        cfg_din5169,
   output        cfg_din5170,
   output        cfg_din5171,
   output        cfg_din5172,
   output        cfg_din5173,
   output        cfg_din5174,
   output        cfg_din5175,
   output        cfg_din5176,
   output        cfg_din5177,
   output        cfg_din5178,
   output        cfg_din5179,
   output        cfg_din5180,
   output        cfg_din5181,
   output        cfg_din5182,
   output        cfg_din5183,
   output        cfg_din5184,
   output        cfg_din5185,
   output        cfg_din5186,
   output        cfg_din5187,
   output        cfg_din5188,
   output        cfg_din5189,
   output        cfg_din5190,
   output        cfg_din5191,
   output        cfg_din5192,
   output        cfg_din5193,
   output        cfg_din5194,
   output        cfg_din5195,
   output        cfg_din5196,
   output        cfg_din5197,
   output        cfg_din5198,
   output        cfg_din5199,
   output        cfg_din5200,
   output        cfg_din5201,
   output        cfg_din5202,
   output        cfg_din5203,
   output        cfg_din5204,
   output        cfg_din5205,
   output        cfg_din5206,
   output        cfg_din5207,
   output        cfg_din5208,
   output        cfg_din5209,
   output        cfg_din5210,
   output        cfg_din5211,
   output        cfg_din5212,
   output        cfg_din5213,
   output        cfg_din5214,
   output        cfg_din5215,
   output        cfg_din5216,
   output        cfg_din5217,
   output        cfg_din5218,
   output        cfg_din5219,
   output        cfg_din5220,
   output        cfg_din5221,
   output        cfg_din5222,
   output        cfg_din5223,
   output        cfg_din5224,
   output        cfg_din5225,
   output        cfg_din5226,
   output        cfg_din5227,
   output        cfg_din5228,
   output        cfg_din5229,
   output        cfg_din5230,
   output        cfg_din5231,
   output        cfg_din5232,
   output        cfg_din5233,
   output        cfg_din5234,
   output        cfg_din5235,
   output        cfg_din5236,
   output        cfg_din5237,
   output        cfg_din5238,
   output        cfg_din5239,
   output        cfg_din5240,
   output        cfg_din5241,
   output        cfg_din5242,
   output        cfg_din5243,
   output        cfg_din5244,
   output        cfg_din5245,
   output        cfg_din5246,
   output        cfg_din5247,
   output        cfg_din5248,
   output        cfg_din5249,
   output        cfg_din5250,
   output        cfg_din5251,
   output        cfg_din5252,
   output        cfg_din5253,
   output        cfg_din5254,
   output        cfg_din5255,
   output        cfg_din5256,
   output        cfg_din5257,
   output        cfg_din5258,
   output        cfg_din5259,
   output        cfg_din5260,
   output        cfg_din5261,
   output        cfg_din5262,
   output        cfg_din5263,
   output        cfg_din5264,
   output        cfg_din5265,
   output        cfg_din5266,
   output        cfg_din5267,
   output        cfg_din5268,
   output        cfg_din5269,
   output        cfg_din5270,
   output        cfg_din5271,
   output        cfg_din5272,
   output        cfg_din5273,
   output        cfg_din5274,
   output        cfg_din5275,
   output        cfg_din5276,
   output        cfg_din5277,
   output        cfg_din5278,
   output        cfg_din5279,
   output        cfg_din5280,
   output        cfg_din5281,
   output        cfg_din5282,
   output        cfg_din5283,
   output        cfg_din5284,
   output        cfg_din5285,
   output        cfg_din5286,
   output        cfg_din5287,
   output        cfg_din5288,
   output        cfg_din5289,
   output        cfg_din5290,
   output        cfg_din5291,
   output        cfg_din5292,
   output        cfg_din5293,
   output        cfg_din5294,
   output        cfg_din5295,
   output        cfg_din5296,
   output        cfg_din5297,
   output        cfg_din5298,
   output        cfg_din5299,
   output        cfg_din5300,
   output        cfg_din5301,
   output        cfg_din5302,
   output        cfg_din5303,
   output        cfg_din5304,
   output        cfg_din5305,
   output        cfg_din5306,
   output        cfg_din5307,
   output        cfg_din5308,
   output        cfg_din5309,
   output        cfg_din5310,
   output        cfg_din5311,
   output        cfg_din5312,
   output        cfg_din5313,
   output        cfg_din5314,
   output        cfg_din5315,
   output        cfg_din5316,
   output        cfg_din5317,
   output        cfg_din5318,
   output        cfg_din5319,
   output        cfg_din5320,
   output        cfg_din5321,
   output        cfg_din5322,
   output        cfg_din5323,
   output        cfg_din5324,
   output        cfg_din5325,
   output        cfg_din5326,
   output        cfg_din5327,
   output        cfg_din5328,
   output        cfg_din5329,
   output        cfg_din5330,
   output        cfg_din5331,
   output        cfg_din5332,
   output        cfg_din5333,
   output        cfg_din5334,
   output        cfg_din5335,
   output        cfg_din5336,
   output        cfg_din5337,
   output        cfg_din5338,
   output        cfg_din5339,
   output        cfg_din5340,
   output        cfg_din5341,
   output        cfg_din5342,
   output        cfg_din5343,
   output        cfg_din5344,
   output        cfg_din5345,
   output        cfg_din5346,
   output        cfg_din5347,
   output        cfg_din5348,
   output        cfg_din5349,
   output        cfg_din5350,
   output        cfg_din5351,
   output        cfg_din5352,
   output        cfg_din5353,
   output        cfg_din5354,
   output        cfg_din5355,
   output        cfg_din5356,
   output        cfg_din5357,
   output        cfg_din5358,
   output        cfg_din5359,
   output        cfg_din5360,
   output        cfg_din5361,
   output        cfg_din5362,
   output        cfg_din5363,
   output        cfg_din5364,
   output        cfg_din5365,
   output        cfg_din5366,
   output        cfg_din5367,
   output        cfg_din5368,
   output        cfg_din5369,
   output        cfg_din5370,
   output        cfg_din5371,
   output        cfg_din5372,
   output        cfg_din5373,
   output        cfg_din5374,
   output        cfg_din5375,
   output        cfg_din5376,
   output        cfg_din5377,
   output        cfg_din5378,
   output        cfg_din5379,
   output        cfg_din5380,
   output        cfg_din5381,
   output        cfg_din5382,
   output        cfg_din5383,
   output        cfg_din5384,
   output        cfg_din5385,
   output        cfg_din5386,
   output        cfg_din5387,
   output        cfg_din5388,
   output        cfg_din5389,
   output        cfg_din5390,
   output        cfg_din5391,
   output        cfg_din5392,
   output        cfg_din5393,
   output        cfg_din5394,
   output        cfg_din5395,
   output        cfg_din5396,
   output        cfg_din5397,
   output        cfg_din5398,
   output        cfg_din5399,
   output        cfg_din5400,
   output        cfg_din5401,
   output        cfg_din5402,
   output        cfg_din5403,
   output        cfg_din5404,
   output        cfg_din5405,
   output        cfg_din5406,
   output        cfg_din5407,
   output        cfg_din5408,
   output        cfg_din5409,
   output        cfg_din5410,
   output        cfg_din5411,
   output        cfg_din5412,
   output        cfg_din5413,
   output        cfg_din5414,
   output        cfg_din5415,
   output        cfg_din5416,
   output        cfg_din5417,
   output        cfg_din5418,
   output        cfg_din5419,
   output        cfg_din5420,
   output        cfg_din5421,
   output        cfg_din5422,
   output        cfg_din5423,
   output        cfg_din5424,
   output        cfg_din5425,
   output        cfg_din5426,
   output        cfg_din5427,
   output        cfg_din5428,
   output        cfg_din5429,
   output        cfg_din5430,
   output        cfg_din5431,
   output        cfg_din5432,
   output        cfg_din5433,
   output        cfg_din5434,
   output        cfg_din5435,
   output        cfg_din5436,
   output        cfg_din5437,
   output        cfg_din5438,
   output        cfg_din5439,
   output        cfg_din5440,
   output        cfg_din5441,
   output        cfg_din5442,
   output        cfg_din5443,
   output        cfg_din5444,
   output        cfg_din5445,
   output        cfg_din5446,
   output        cfg_din5447,
   output        cfg_din5448,
   output        cfg_din5449,
   output        cfg_din5450,
   output        cfg_din5451,
   output        cfg_din5452,
   output        cfg_din5453,
   output        cfg_din5454,
   output        cfg_din5455,
   output        cfg_din5456,
   output        cfg_din5457,
   output        cfg_din5458,
   output        cfg_din5459,
   output        cfg_din5460,
   output        cfg_din5461,
   output        cfg_din5462,
   output        cfg_din5463,
   output        cfg_din5464,
   output        cfg_din5465,
   output        cfg_din5466,
   output        cfg_din5467,
   output        cfg_din5468,
   output        cfg_din5469,
   output        cfg_din5470,
   output        cfg_din5471,
   output        cfg_din5472,
   output        cfg_din5473,
   output        cfg_din5474,
   output        cfg_din5475,
   output        cfg_din5476,
   output        cfg_din5477,
   output        cfg_din5478,
   output        cfg_din5479,
   output        cfg_din5480,
   output        cfg_din5481,
   output        cfg_din5482,
   output        cfg_din5483,
   output        cfg_din5484,
   output        cfg_din5485,
   output        cfg_din5486,
   output        cfg_din5487,
   output        cfg_din5488,
   output        cfg_din5489,
   output        cfg_din5490,
   output        cfg_din5491,
   output        cfg_din5492,
   output        cfg_din5493,
   output        cfg_din5494,
   output        cfg_din5495,
   output        cfg_din5496,
   output        cfg_din5497,
   output        cfg_din5498,
   output        cfg_din5499,
   output        cfg_din5500,
   output        cfg_din5501,
   output        cfg_din5502,
   output        cfg_din5503,
   output        cfg_din5504,
   output        cfg_din5505,
   output        cfg_din5506,
   output        cfg_din5507,
   output        cfg_din5508,
   output        cfg_din5509,
   output        cfg_din5510,
   output        cfg_din5511,
   output        cfg_din5512,
   output        cfg_din5513,
   output        cfg_din5514,
   output        cfg_din5515,
   output        cfg_din5516,
   output        cfg_din5517,
   output        cfg_din5518,
   output        cfg_din5519,
   output        cfg_din5520,
   output        cfg_din5521,
   output        cfg_din5522,
   output        cfg_din5523,
   output        cfg_din5524,
   output        cfg_din5525,
   output        cfg_din5526,
   output        cfg_din5527,
   output        cfg_din5528,
   output        cfg_din5529,
   output        cfg_din5530,
   output        cfg_din5531,
   output        cfg_din5532,
   output        cfg_din5533,
   output        cfg_din5534,
   output        cfg_din5535,
   output        cfg_din5536,
   output        cfg_din5537,
   output        cfg_din5538,
   output        cfg_din5539,
   output        cfg_din5540,
   output        cfg_din5541,
   output        cfg_din5542,
   output        cfg_din5543,
   output        cfg_din5544,
   output        cfg_din5545,
   output        cfg_din5546,
   output        cfg_din5547,
   output        cfg_din5548,
   output        cfg_din5549,
   output        cfg_din5550,
   output        cfg_din5551,
   output        cfg_din5552,
   output        cfg_din5553,
   output        cfg_din5554,
   output        cfg_din5555,
   output        cfg_din5556,
   output        cfg_din5557,
   output        cfg_din5558,
   output        cfg_din5559,
   output        cfg_din5560,
   output        cfg_din5561,
   output        cfg_din5562,
   output        cfg_din5563,
   output        cfg_din5564,
   output        cfg_din5565,
   output        cfg_din5566,
   output        cfg_din5567,
   output        cfg_din5568,
   output        cfg_din5569,
   output        cfg_din5570,
   output        cfg_din5571,
   output        cfg_din5572,
   output        cfg_din5573,
   output        cfg_din5574,
   output        cfg_din5575,
   output        cfg_din5576,
   output        cfg_din5577,
   output        cfg_din5578,
   output        cfg_din5579,
   output        cfg_din5580,
   output        cfg_din5581,
   output        cfg_din5582,
   output        cfg_din5583,
   output        cfg_din5584,
   output        cfg_din5585,
   output        cfg_din5586,
   output        cfg_din5587,
   output        cfg_din5588,
   output        cfg_din5589,
   output        cfg_din5590,
   output        cfg_din5591,
   output        cfg_din5592,
   output        cfg_din5593,
   output        cfg_din5594,
   output        cfg_din5595,
   output        cfg_din5596,
   output        cfg_din5597,
   output        cfg_din5598,
   output        cfg_din5599,
   output        cfg_din5600,
   output        cfg_din5601,
   output        cfg_din5602,
   output        cfg_din5603,
   output        cfg_din5604,
   output        cfg_din5605,
   output        cfg_din5606,
   output        cfg_din5607,
   output        cfg_din5608,
   output        cfg_din5609,
   output        cfg_din5610,
   output        cfg_din5611,
   output        cfg_din5612,
   output        cfg_din5613,
   output        cfg_din5614,
   output        cfg_din5615,
   output        cfg_din5616,
   output        cfg_din5617,
   output        cfg_din5618,
   output        cfg_din5619,
   output        cfg_din5620,
   output        cfg_din5621,
   output        cfg_din5622,
   output        cfg_din5623,
   output        cfg_din5624,
   output        cfg_din5625,
   output        cfg_din5626,
   output        cfg_din5627,
   output        cfg_din5628,
   output        cfg_din5629,
   output        cfg_din5630,
   output        cfg_din5631,
   output        cfg_din5632,
   output        cfg_din5633,
   output        cfg_din5634,
   output        cfg_din5635,
   output        cfg_din5636,
   output        cfg_din5637,
   output        cfg_din5638,
   output        cfg_din5639,
   output        cfg_din5640,
   output        cfg_din5641,
   output        cfg_din5642,
   output        cfg_din5643,
   output        cfg_din5644,
   output        cfg_din5645,
   output        cfg_din5646,
   output        cfg_din5647,
   output        cfg_din5648,
   output        cfg_din5649,
   output        cfg_din5650,
   output        cfg_din5651,
   output        cfg_din5652,
   output        cfg_din5653,
   output        cfg_din5654,
   output        cfg_din5655,
   output        cfg_din5656,
   output        cfg_din5657,
   output        cfg_din5658,
   output        cfg_din5659,
   output        cfg_din5660,
   output        cfg_din5661,
   output        cfg_din5662,
   output        cfg_din5663,
   output        cfg_din5664,
   output        cfg_din5665,
   output        cfg_din5666,
   output        cfg_din5667,
   output        cfg_din5668,
   output        cfg_din5669,
   output        cfg_din5670,
   output        cfg_din5671,
   output        cfg_din5672,
   output        cfg_din5673,
   output        cfg_din5674,
   output        cfg_din5675,
   output        cfg_din5676,
   output        cfg_din5677,
   output        cfg_din5678,
   output        cfg_din5679,
   output        cfg_din5680,
   output        cfg_din5681,
   output        cfg_din5682,
   output        cfg_din5683,
   output        cfg_din5684,
   output        cfg_din5685,
   output        cfg_din5686,
   output        cfg_din5687,
   output        cfg_din5688,
   output        cfg_din5689,
   output        cfg_din5690,
   output        cfg_din5691,
   output        cfg_din5692,
   output        cfg_din5693,
   output        cfg_din5694,
   output        cfg_din5695,
   output        cfg_din5696,
   output        cfg_din5697,
   output        cfg_din5698,
   output        cfg_din5699,
   output        cfg_din5700,
   output        cfg_din5701,
   output        cfg_din5702,
   output        cfg_din5703,
   output        cfg_din5704,
   output        cfg_din5705,
   output        cfg_din5706,
   output        cfg_din5707,
   output        cfg_din5708,
   output        cfg_din5709,
   output        cfg_din5710,
   output        cfg_din5711,
   output        cfg_din5712,
   output        cfg_din5713,
   output        cfg_din5714,
   output        cfg_din5715,
   output        cfg_din5716,
   output        cfg_din5717,
   output        cfg_din5718,
   output        cfg_din5719,
   output        cfg_din5720,
   output        cfg_din5721,
   output        cfg_din5722,
   output        cfg_din5723,
   output        cfg_din5724,
   output        cfg_din5725,
   output        cfg_din5726,
   output        cfg_din5727,
   output        cfg_din5728,
   output        cfg_din5729,
   output        cfg_din5730,
   output        cfg_din5731,
   output        cfg_din5732,
   output        cfg_din5733,
   output        cfg_din5734,
   output        cfg_din5735,
   output        cfg_din5736,
   output        cfg_din5737,
   output        cfg_din5738,
   output        cfg_din5739,
   output        cfg_din5740,
   output        cfg_din5741,
   output        cfg_din5742,
   output        cfg_din5743,
   output        cfg_din5744,
   output        cfg_din5745,
   output        cfg_din5746,
   output        cfg_din5747,
   output        cfg_din5748,
   output        cfg_din5749,
   output        cfg_din5750,
   output        cfg_din5751,
   output        cfg_din5752,
   output        cfg_din5753,
   output        cfg_din5754,
   output        cfg_din5755,
   output        cfg_din5756,
   output        cfg_din5757,
   output        cfg_din5758,
   output        cfg_din5759,
   output        cfg_din5760,
   output        cfg_din5761,
   output        cfg_din5762,
   output        cfg_din5763,
   output        cfg_din5764,
   output        cfg_din5765,
   output        cfg_din5766,
   output        cfg_din5767,
   output        cfg_din5768,
   output        cfg_din5769,
   output        cfg_din5770,
   output        cfg_din5771,
   output        cfg_din5772,
   output        cfg_din5773,
   output        cfg_din5774,
   output        cfg_din5775,
   output        cfg_din5776,
   output        cfg_din5777,
   output        cfg_din5778,
   output        cfg_din5779,
   output        cfg_din5780,
   output        cfg_din5781,
   output        cfg_din5782,
   output        cfg_din5783,
   output        cfg_din5784,
   output        cfg_din5785,
   output        cfg_din5786,
   output        cfg_din5787,
   output        cfg_din5788,
   output        cfg_din5789,
   output        cfg_din5790,
   output        cfg_din5791,
   output        cfg_din5792,
   output        cfg_din5793,
   output        cfg_din5794,
   output        cfg_din5795,
   output        cfg_din5796,
   output        cfg_din5797,
   output        cfg_din5798,
   output        cfg_din5799,
   output        cfg_din5800,
   output        cfg_din5801,
   output        cfg_din5802,
   output        cfg_din5803,
   output        cfg_din5804,
   output        cfg_din5805,
   output        cfg_din5806,
   output        cfg_din5807,
   output        cfg_din5808,
   output        cfg_din5809,
   output        cfg_din5810,
   output        cfg_din5811,
   output        cfg_din5812,
   output        cfg_din5813,
   output        cfg_din5814,
   output        cfg_din5815,
   output        cfg_din5816,
   output        cfg_din5817,
   output        cfg_din5818,
   output        cfg_din5819,
   output        cfg_din5820,
   output        cfg_din5821,
   output        cfg_din5822,
   output        cfg_din5823,
   output        cfg_din5824,
   output        cfg_din5825,
   output        cfg_din5826,
   output        cfg_din5827,
   output        cfg_din5828,
   output        cfg_din5829,
   output        cfg_din5830,
   output        cfg_din5831,
   output        cfg_din5832,
   output        cfg_din5833,
   output        cfg_din5834,
   output        cfg_din5835,
   output        cfg_din5836,
   output        cfg_din5837,
   output        cfg_din5838,
   output        cfg_din5839,
   output        cfg_din5840,
   output        cfg_din5841,
   output        cfg_din5842,
   output        cfg_din5843,
   output        cfg_din5844,
   output        cfg_din5845,
   output        cfg_din5846,
   output        cfg_din5847,
   output        cfg_din5848,
   output        cfg_din5849,
   output        cfg_din5850,
   output        cfg_din5851,
   output        cfg_din5852,
   output        cfg_din5853,
   output        cfg_din5854,
   output        cfg_din5855,
   output        cfg_din5856,
   output        cfg_din5857,
   output        cfg_din5858,
   output        cfg_din5859,
   output        cfg_din5860,
   output        cfg_din5861,
   output        cfg_din5862,
   output        cfg_din5863,
   output        cfg_din5864,
   output        cfg_din5865,
   output        cfg_din5866,
   output        cfg_din5867,
   output        cfg_din5868,
   output        cfg_din5869,
   output        cfg_din5870,
   output        cfg_din5871,
   output        cfg_din5872,
   output        cfg_din5873,
   output        cfg_din5874,
   output        cfg_din5875,
   output        cfg_din5876,
   output        cfg_din5877,
   output        cfg_din5878,
   output        cfg_din5879,
   output        cfg_din5880,
   output        cfg_din5881,
   output        cfg_din5882,
   output        cfg_din5883,
   output        cfg_din5884,
   output        cfg_din5885,
   output        cfg_din5886,
   output        cfg_din5887,
   output        cfg_din5888,
   output        cfg_din5889,
   output        cfg_din5890,
   output        cfg_din5891,
   output        cfg_din5892,
   output        cfg_din5893,
   output        cfg_din5894,
   output        cfg_din5895,
   output        cfg_din5896,
   output        cfg_din5897,
   output        cfg_din5898,
   output        cfg_din5899,
   output        cfg_din5900,
   output        cfg_din5901,
   output        cfg_din5902,
   output        cfg_din5903,
   output        cfg_din5904,
   output        cfg_din5905,
   output        cfg_din5906,
   output        cfg_din5907,
   output        cfg_din5908,
   output        cfg_din5909,
   output        cfg_din5910,
   output        cfg_din5911,
   output        cfg_din5912,
   output        cfg_din5913,
   output        cfg_din5914,
   output        cfg_din5915,
   output        cfg_din5916,
   output        cfg_din5917,
   output        cfg_din5918,
   output        cfg_din5919,
   output        cfg_din5920,
   output        cfg_din5921,
   output        cfg_din5922,
   output        cfg_din5923,
   output        cfg_din5924,
   output        cfg_din5925,
   output        cfg_din5926,
   output        cfg_din5927,
   output        cfg_din5928,
   output        cfg_din5929,
   output        cfg_din5930,
   output        cfg_din5931,
   output        cfg_din5932,
   output        cfg_din5933,
   output        cfg_din5934,
   output        cfg_din5935,
   output        cfg_din5936,
   output        cfg_din5937,
   output        cfg_din5938,
   output        cfg_din5939,
   output        cfg_din5940,
   output        cfg_din5941,
   output        cfg_din5942,
   output        cfg_din5943,
   output        cfg_din5944,
   output        cfg_din5945,
   output        cfg_din5946,
   output        cfg_din5947,
   output        cfg_din5948,
   output        cfg_din5949,
   output        cfg_din5950,
   output        cfg_din5951,
   output        cfg_din5952,
   output        cfg_din5953,
   output        cfg_din5954,
   output        cfg_din5955,
   output        cfg_din5956,
   output        cfg_din5957,
   output        cfg_din5958,
   output        cfg_din5959,
   output        cfg_din5960,
   output        cfg_din5961,
   output        cfg_din5962,
   output        cfg_din5963,
   output        cfg_din5964,
   output        cfg_din5965,
   output        cfg_din5966,
   output        cfg_din5967,
   output        cfg_din5968,
   output        cfg_din5969,
   output        cfg_din5970,
   output        cfg_din5971,
   output        cfg_din5972,
   output        cfg_din5973,
   output        cfg_din5974,
   output        cfg_din5975,
   output        cfg_din5976,
   output        cfg_din5977,
   output        cfg_din5978,
   output        cfg_din5979,
   output        cfg_din5980,
   output        cfg_din5981,
   output        cfg_din5982,
   output        cfg_din5983,
   output        cfg_din5984,
   output        cfg_din5985,
   output        cfg_din5986,
   output        cfg_din5987,
   output        cfg_din5988,
   output        cfg_din5989,
   output        cfg_din5990,
   output        cfg_din5991,
   output        cfg_din5992,
   output        cfg_din5993,
   output        cfg_din5994,
   output        cfg_din5995,
   output        cfg_din5996,
   output        cfg_din5997,
   output        cfg_din5998,
   output        cfg_din5999,
   output        cfg_din6000,
   output        cfg_din6001,
   output        cfg_din6002,
   output        cfg_din6003,
   output        cfg_din6004,
   output        cfg_din6005,
   output        cfg_din6006,
   output        cfg_din6007,
   output        cfg_din6008,
   output        cfg_din6009,
   output        cfg_din6010,
   output        cfg_din6011,
   output        cfg_din6012,
   output        cfg_din6013,
   output        cfg_din6014,
   output        cfg_din6015,
   output        cfg_din6016,
   output        cfg_din6017,
   output        cfg_din6018,
   output        cfg_din6019,
   output        cfg_din6020,
   output        cfg_din6021,
   output        cfg_din6022,
   output        cfg_din6023,
   output        cfg_din6024,
   output        cfg_din6025,
   output        cfg_din6026,
   output        cfg_din6027,
   output        cfg_din6028,
   output        cfg_din6029,
   output        cfg_din6030,
   output        cfg_din6031,
   output        cfg_din6032,
   output        cfg_din6033,
   output        cfg_din6034,
   output        cfg_din6035,
   output        cfg_din6036,
   output        cfg_din6037,
   output        cfg_din6038,
   output        cfg_din6039,
   output        cfg_din6040,
   output        cfg_din6041,
   output        cfg_din6042,
   output        cfg_din6043,
   output        cfg_din6044,
   output        cfg_din6045,
   output        cfg_din6046,
   output        cfg_din6047,
   output        cfg_din6048,
   output        cfg_din6049,
   output        cfg_din6050,
   output        cfg_din6051,
   output        cfg_din6052,
   output        cfg_din6053,
   output        cfg_din6054,
   output        cfg_din6055,
   output        cfg_din6056,
   output        cfg_din6057,
   output        cfg_din6058,
   output        cfg_din6059,
   output        cfg_din6060,
   output        cfg_din6061,
   output        cfg_din6062,
   output        cfg_din6063,
   output        cfg_din6064,
   output        cfg_din6065,
   output        cfg_din6066,
   output        cfg_din6067,
   output        cfg_din6068,
   output        cfg_din6069,
   output        cfg_din6070,
   output        cfg_din6071,
   output        cfg_din6072,
   output        cfg_din6073,
   output        cfg_din6074,
   output        cfg_din6075,
   output        cfg_din6076,
   output        cfg_din6077,
   output        cfg_din6078,
   output        cfg_din6079,
   output        cfg_din6080,
   output        cfg_din6081,
   output        cfg_din6082,
   output        cfg_din6083,
   output        cfg_din6084,
   output        cfg_din6085,
   output        cfg_din6086,
   output        cfg_din6087,
   output        cfg_din6088,
   output        cfg_din6089,
   output        cfg_din6090,
   output        cfg_din6091,
   output        cfg_din6092,
   output        cfg_din6093,
   output        cfg_din6094,
   output        cfg_din6095,
   output        cfg_din6096,
   output        cfg_din6097,
   output        cfg_din6098,
   output        cfg_din6099,
   output        cfg_din6100,
   output        cfg_din6101,
   output        cfg_din6102,
   output        cfg_din6103,
   output        cfg_din6104,
   output        cfg_din6105,
   output        cfg_din6106,
   output        cfg_din6107,
   output        cfg_din6108,
   output        cfg_din6109,
   output        cfg_din6110,
   output        cfg_din6111,
   output        cfg_din6112,
   output        cfg_din6113,
   output        cfg_din6114,
   output        cfg_din6115,
   output        cfg_din6116,
   output        cfg_din6117,
   output        cfg_din6118,
   output        cfg_din6119,
   output        cfg_din6120,
   output        cfg_din6121,
   output        cfg_din6122,
   output        cfg_din6123,
   output        cfg_din6124,
   output        cfg_din6125,
   output        cfg_din6126,
   output        cfg_din6127,
   output        cfg_din6128,
   output        cfg_din6129,
   output        cfg_din6130,
   output        cfg_din6131,
   output        cfg_din6132,
   output        cfg_din6133,
   output        cfg_din6134,
   output        cfg_din6135,
   output        cfg_din6136,
   output        cfg_din6137,
   output        cfg_din6138,
   output        cfg_din6139,
   output        cfg_din6140,
   output        cfg_din6141,
   output        cfg_din6142,
   output        cfg_din6143,
   output        cfg_din6144,
   output        cfg_din6145,
   output        cfg_din6146,
   output        cfg_din6147,
   output        cfg_din6148,
   output        cfg_din6149,
   output        cfg_din6150,
   output        cfg_din6151,
   output        cfg_din6152,
   output        cfg_din6153,
   output        cfg_din6154,
   output        cfg_din6155,
   output        cfg_din6156,
   output        cfg_din6157,
   output        cfg_din6158,
   output        cfg_din6159,
   output        cfg_din6160,
   output        cfg_din6161,
   output        cfg_din6162,
   output        cfg_din6163,
   output        cfg_din6164,
   output        cfg_din6165,
   output        cfg_din6166,
   output        cfg_din6167,
   output        cfg_din6168,
   output        cfg_din6169,
   output        cfg_din6170,
   output        cfg_din6171,
   output        cfg_din6172,
   output        cfg_din6173,
   output        cfg_din6174,
   output        cfg_din6175,
   output        cfg_din6176,
   output        cfg_din6177,
   output        cfg_din6178,
   output        cfg_din6179,
   output        cfg_din6180,
   output        cfg_din6181,
   output        cfg_din6182,
   output        cfg_din6183,
   output        cfg_din6184,
   output        cfg_din6185,
   output        cfg_din6186,
   output        cfg_din6187,
   output        cfg_din6188,
   output        cfg_din6189,
   output        cfg_din6190,
   output        cfg_din6191,
   output        cfg_din6192,
   output        cfg_din6193,
   output        cfg_din6194,
   output        cfg_din6195,
   output        cfg_din6196,
   output        cfg_din6197,
   output        cfg_din6198,
   output        cfg_din6199,
   output        cfg_din6200,
   output        cfg_din6201,
   output        cfg_din6202,
   output        cfg_din6203,
   output        cfg_din6204,
   output        cfg_din6205,
   output        cfg_din6206,
   output        cfg_din6207,
   output        cfg_din6208,
   output        cfg_din6209,
   output        cfg_din6210,
   output        cfg_din6211,
   output        cfg_din6212,
   output        cfg_din6213,
   output        cfg_din6214,
   output        cfg_din6215,
   output        cfg_din6216,
   output        cfg_din6217,
   output        cfg_din6218,
   output        cfg_din6219,
   output        cfg_din6220,
   output        cfg_din6221,
   output        cfg_din6222,
   output        cfg_din6223,
   output        cfg_din6224,
   output        cfg_din6225,
   output        cfg_din6226,
   output        cfg_din6227,
   output        cfg_din6228,
   output        cfg_din6229,
   output        cfg_din6230,
   output        cfg_din6231,
   output        cfg_din6232,
   output        cfg_din6233,
   output        cfg_din6234,
   output        cfg_din6235,
   output        cfg_din6236,
   output        cfg_din6237,
   output        cfg_din6238,
   output        cfg_din6239,
   output        cfg_din6240,
   output        cfg_din6241,
   output        cfg_din6242,
   output        cfg_din6243,
   output        cfg_din6244,
   output        cfg_din6245,
   output        cfg_din6246,
   output        cfg_din6247,
   output        cfg_din6248,
   output        cfg_din6249,
   output        cfg_din6250,
   output        cfg_din6251,
   output        cfg_din6252,
   output        cfg_din6253,
   output        cfg_din6254,
   output        cfg_din6255,
   output        cfg_din6256,
   output        cfg_din6257,
   output        cfg_din6258,
   output        cfg_din6259,
   output        cfg_din6260,
   output        cfg_din6261,
   output        cfg_din6262,
   output        cfg_din6263,
   output        cfg_din6264,
   output        cfg_din6265,
   output        cfg_din6266,
   output        cfg_din6267,
   output        cfg_din6268,
   output        cfg_din6269,
   output        cfg_din6270,
   output        cfg_din6271,
   output        cfg_din6272,
   output        cfg_din6273,
   output        cfg_din6274,
   output        cfg_din6275,
   output        cfg_din6276,
   output        cfg_din6277,
   output        cfg_din6278,
   output        cfg_din6279,
   output        cfg_din6280,
   output        cfg_din6281,
   output        cfg_din6282,
   output        cfg_din6283,
   output        cfg_din6284,
   output        cfg_din6285,
   output        cfg_din6286,
   output        cfg_din6287,
   output        cfg_din6288,
   output        cfg_din6289,
   output        cfg_din6290,
   output        cfg_din6291,
   output        cfg_din6292,
   output        cfg_din6293,
   output        cfg_din6294,
   output        cfg_din6295,
   output        cfg_din6296,
   output        cfg_din6297,
   output        cfg_din6298,
   output        cfg_din6299,
   output        cfg_din6300,
   output        cfg_din6301,
   output        cfg_din6302,
   output        cfg_din6303,
   output        cfg_din6304,
   output        cfg_din6305,
   output        cfg_din6306,
   output        cfg_din6307,
   output        cfg_din6308,
   output        cfg_din6309,
   output        cfg_din6310,
   output        cfg_din6311,
   output        cfg_din6312,
   output        cfg_din6313,
   output        cfg_din6314,
   output        cfg_din6315,
   output        cfg_din6316,
   output        cfg_din6317,
   output        cfg_din6318,
   output        cfg_din6319,
   output        cfg_din6320,
   output        cfg_din6321,
   output        cfg_din6322,
   output        cfg_din6323,
   output        cfg_din6324,
   output        cfg_din6325,
   output        cfg_din6326,
   output        cfg_din6327,
   output        cfg_din6328,
   output        cfg_din6329,
   output        cfg_din6330,
   output        cfg_din6331,
   output        cfg_din6332,
   output        cfg_din6333,
   output        cfg_din6334,
   output        cfg_din6335,
   output        cfg_din6336,
   output        cfg_din6337,
   output        cfg_din6338,
   output        cfg_din6339,
   output        cfg_din6340,
   output        cfg_din6341,
   output        cfg_din6342,
   output        cfg_din6343,
   output        cfg_din6344,
   output        cfg_din6345,
   output        cfg_din6346,
   output        cfg_din6347,
   output        cfg_din6348,
   output        cfg_din6349,
   output        cfg_din6350,
   output        cfg_din6351,
   output        cfg_din6352,
   output        cfg_din6353,
   output        cfg_din6354,
   output        cfg_din6355,
   output        cfg_din6356,
   output        cfg_din6357,
   output        cfg_din6358,
   output        cfg_din6359,
   output        cfg_din6360,
   output        cfg_din6361,
   output        cfg_din6362,
   output        cfg_din6363,
   output        cfg_din6364,
   output        cfg_din6365,
   output        cfg_din6366,
   output        cfg_din6367,
   output        cfg_din6368,
   output        cfg_din6369,
   output        cfg_din6370,
   output        cfg_din6371,
   output        cfg_din6372,
   output        cfg_din6373,
   output        cfg_din6374,
   output        cfg_din6375,
   output        cfg_din6376,
   output        cfg_din6377,
   output        cfg_din6378,
   output        cfg_din6379,
   output        cfg_din6380,
   output        cfg_din6381,
   output        cfg_din6382,
   output        cfg_din6383,
   output        cfg_din6384,
   output        cfg_din6385,
   output        cfg_din6386,
   output        cfg_din6387,
   output        cfg_din6388,
   output        cfg_din6389,
   output        cfg_din6390,
   output        cfg_din6391,
   output        cfg_din6392,
   output        cfg_din6393,
   output        cfg_din6394,
   output        cfg_din6395,
   output        cfg_din6396,
   output        cfg_din6397,
   output        cfg_din6398,
   output        cfg_din6399,
   output        cfg_din6400,
   output        cfg_din6401,
   output        cfg_din6402,
   output        cfg_din6403,
   output        cfg_din6404,
   output        cfg_din6405,
   output        cfg_din6406,
   output        cfg_din6407,
   output        cfg_din6408,
   output        cfg_din6409,
   output        cfg_din6410,
   output        cfg_din6411,
   output        cfg_din6412,
   output        cfg_din6413,
   output        cfg_din6414,
   output        cfg_din6415,
   output        cfg_din6416,
   output        cfg_din6417,
   output        cfg_din6418,
   output        cfg_din6419,
   output        cfg_din6420,
   output        cfg_din6421,
   output        cfg_din6422,
   output        cfg_din6423,
   output        cfg_din6424,
   output        cfg_din6425,
   output        cfg_din6426,
   output        cfg_din6427,
   output        cfg_din6428,
   output        cfg_din6429,
   output        cfg_din6430,
   output        cfg_din6431,
   output        cfg_din6432,
   output        cfg_din6433,
   output        cfg_din6434,
   output        cfg_din6435,
   output        cfg_din6436,
   output        cfg_din6437,
   output        cfg_din6438,
   output        cfg_din6439,
   output        cfg_din6440,
   output        cfg_din6441,
   output        cfg_din6442,
   output        cfg_din6443,
   output        cfg_din6444,
   output        cfg_din6445,
   output        cfg_din6446,
   output        cfg_din6447,
   output        cfg_din6448,
   output        cfg_din6449,
   output        cfg_din6450,
   output        cfg_din6451,
   output        cfg_din6452,
   output        cfg_din6453,
   output        cfg_din6454,
   output        cfg_din6455,
   output        cfg_din6456,
   output        cfg_din6457,
   output        cfg_din6458,
   output        cfg_din6459,
   output        cfg_din6460,
   output        cfg_din6461,
   output        cfg_din6462,
   output        cfg_din6463,
   output        cfg_din6464,
   output        cfg_din6465,
   output        cfg_din6466,
   output        cfg_din6467,
   output        cfg_din6468,
   output        cfg_din6469,
   output        cfg_din6470,
   output        cfg_din6471,
   output        cfg_din6472,
   output        cfg_din6473,
   output        cfg_din6474,
   output        cfg_din6475,
   output        cfg_din6476,
   output        cfg_din6477,
   output        cfg_din6478,
   output        cfg_din6479,
   output        cfg_din6480,
   output        cfg_din6481,
   output        cfg_din6482,
   output        cfg_din6483,
   output        cfg_din6484,
   output        cfg_din6485,
   output        cfg_din6486,
   output        cfg_din6487,
   output        cfg_din6488,
   output        cfg_din6489,
   output        cfg_din6490,
   output        cfg_din6491,
   output        cfg_din6492,
   output        cfg_din6493,
   output        cfg_din6494,
   output        cfg_din6495,
   output        cfg_din6496,
   output        cfg_din6497,
   output        cfg_din6498,
   output        cfg_din6499,
   output        cfg_din6500,
   output        cfg_din6501,
   output        cfg_din6502,
   output        cfg_din6503,
   output        cfg_din6504,
   output        cfg_din6505,
   output        cfg_din6506,
   output        cfg_din6507,
   output        cfg_din6508,
   output        cfg_din6509,
   output        cfg_din6510,
   output        cfg_din6511,
   output        cfg_din6512,
   output        cfg_din6513,
   output        cfg_din6514,
   output        cfg_din6515,
   output        cfg_din6516,
   output        cfg_din6517,
   output        cfg_din6518,
   output        cfg_din6519,
   output        cfg_din6520,
   output        cfg_din6521,
   output        cfg_din6522,
   output        cfg_din6523,
   output        cfg_din6524,
   output        cfg_din6525,
   output        cfg_din6526,
   output        cfg_din6527,
   output        cfg_din6528,
   output        cfg_din6529,
   output        cfg_din6530,
   output        cfg_din6531,
   output        cfg_din6532,
   output        cfg_din6533,
   output        cfg_din6534,
   output        cfg_din6535,
   output        cfg_din6536,
   output        cfg_din6537,
   output        cfg_din6538,
   output        cfg_din6539,
   output        cfg_din6540,
   output        cfg_din6541,
   output        cfg_din6542,
   output        cfg_din6543,
   output        cfg_din6544,
   output        cfg_din6545,
   output        cfg_din6546,
   output        cfg_din6547,
   output        cfg_din6548,
   output        cfg_din6549,
   output        cfg_din6550,
   output        cfg_din6551,
   output        cfg_din6552,
   output        cfg_din6553,
   output        cfg_din6554,
   output        cfg_din6555,
   output        cfg_din6556,
   output        cfg_din6557,
   output        cfg_din6558,
   output        cfg_din6559,
   output        cfg_din6560,
   output        cfg_din6561,
   output        cfg_din6562,
   output        cfg_din6563,
   output        cfg_din6564,
   output        cfg_din6565,
   output        cfg_din6566,
   output        cfg_din6567,
   output        cfg_din6568,
   output        cfg_din6569,
   output        cfg_din6570,
   output        cfg_din6571,
   output        cfg_din6572,
   output        cfg_din6573,
   output        cfg_din6574,
   output        cfg_din6575,
   output        cfg_din6576,
   output        cfg_din6577,
   output        cfg_din6578,
   output        cfg_din6579,
   output        cfg_din6580,
   output        cfg_din6581,
   output        cfg_din6582,
   output        cfg_din6583,
   output        cfg_din6584,
   output        cfg_din6585,
   output        cfg_din6586,
   output        cfg_din6587,
   output        cfg_din6588,
   output        cfg_din6589,
   output        cfg_din6590,
   output        cfg_din6591,
   output        cfg_din6592,
   output        cfg_din6593,
   output        cfg_din6594,
   output        cfg_din6595,
   output        cfg_din6596,
   output        cfg_din6597,
   output        cfg_din6598,
   output        cfg_din6599,
   output        cfg_din6600,
   output        cfg_din6601,
   output        cfg_din6602,
   output        cfg_din6603,
   output        cfg_din6604,
   output        cfg_din6605,
   output        cfg_din6606,
   output        cfg_din6607,
   output        cfg_din6608,
   output        cfg_din6609,
   output        cfg_din6610,
   output        cfg_din6611,
   output        cfg_din6612,
   output        cfg_din6613,
   output        cfg_din6614,
   output        cfg_din6615,
   output        cfg_din6616,
   output        cfg_din6617,
   output        cfg_din6618,
   output        cfg_din6619,
   output        cfg_din6620,
   output        cfg_din6621,
   output        cfg_din6622,
   output        cfg_din6623,
   output        cfg_din6624,
   output        cfg_din6625,
   output        cfg_din6626,
   output        cfg_din6627,
   output        cfg_din6628,
   output        cfg_din6629,
   output        cfg_din6630,
   output        cfg_din6631,
   output        cfg_din6632,
   output        cfg_din6633,
   output        cfg_din6634,
   output        cfg_din6635,
   output        cfg_din6636,
   output        cfg_din6637,
   output        cfg_din6638,
   output        cfg_din6639,
   output        cfg_din6640,
   output        cfg_din6641,
   output        cfg_din6642,
   output        cfg_din6643,
   output        cfg_din6644,
   output        cfg_din6645,
   output        cfg_din6646,
   output        cfg_din6647,
   output        cfg_din6648,
   output        cfg_din6649,
   output        cfg_din6650,
   output        cfg_din6651,
   output        cfg_din6652,
   output        cfg_din6653,
   output        cfg_din6654,
   output        cfg_din6655,
   output        cfg_din6656,
   output        cfg_din6657,
   output        cfg_din6658,
   output        cfg_din6659,
   output        cfg_din6660,
   output        cfg_din6661,
   output        cfg_din6662,
   output        cfg_din6663,
   output        cfg_din6664,
   output        cfg_din6665,
   output        cfg_din6666,
   output        cfg_din6667,
   output        cfg_din6668,
   output        cfg_din6669,
   output        cfg_din6670,
   output        cfg_din6671,
   output        cfg_din6672,
   output        cfg_din6673,
   output        cfg_din6674,
   output        cfg_din6675,
   output        cfg_din6676,
   output        cfg_din6677,
   output        cfg_din6678,
   output        cfg_din6679,
   output        cfg_din6680,
   output        cfg_din6681,
   output        cfg_din6682,
   output        cfg_din6683,
   output        cfg_din6684,
   output        cfg_din6685,
   output        cfg_din6686,
   output        cfg_din6687,
   output        cfg_din6688,
   output        cfg_din6689,
   output        cfg_din6690,
   output        cfg_din6691,
   output        cfg_din6692,
   output        cfg_din6693,
   output        cfg_din6694,
   output        cfg_din6695,
   output        cfg_din6696,
   output        cfg_din6697,
   output        cfg_din6698,
   output        cfg_din6699,
   output        cfg_din6700,
   output        cfg_din6701,
   output        cfg_din6702,
   output        cfg_din6703,
   output        cfg_din6704,
   output        cfg_din6705,
   output        cfg_din6706,
   output        cfg_din6707,
   output        cfg_din6708,
   output        cfg_din6709,
   output        cfg_din6710,
   output        cfg_din6711,
   output        cfg_din6712,
   output        cfg_din6713,
   output        cfg_din6714,
   output        cfg_din6715,
   output        cfg_din6716,
   output        cfg_din6717,
   output        cfg_din6718,
   output        cfg_din6719,
   output        cfg_din6720,
   output        cfg_din6721,
   output        cfg_din6722,
   output        cfg_din6723,
   output        cfg_din6724,
   output        cfg_din6725,
   output        cfg_din6726,
   output        cfg_din6727,
   output        cfg_din6728,
   output        cfg_din6729,
   output        cfg_din6730,
   output        cfg_din6731,
   output        cfg_din6732,
   output        cfg_din6733,
   output        cfg_din6734,
   output        cfg_din6735,
   output        cfg_din6736,
   output        cfg_din6737,
   output        cfg_din6738,
   output        cfg_din6739,
   output        cfg_din6740,
   output        cfg_din6741,
   output        cfg_din6742,
   output        cfg_din6743,
   output        cfg_din6744,
   output        cfg_din6745,
   output        cfg_din6746,
   output        cfg_din6747,
   output        cfg_din6748,
   output        cfg_din6749,
   output        cfg_din6750,
   output        cfg_din6751,
   output        cfg_din6752,
   output        cfg_din6753,
   output        cfg_din6754,
   output        cfg_din6755,
   output        cfg_din6756,
   output        cfg_din6757,
   output        cfg_din6758,
   output        cfg_din6759,
   output        cfg_din6760,
   output        cfg_din6761,
   output        cfg_din6762,
   output        cfg_din6763,
   output        cfg_din6764,
   output        cfg_din6765,
   output        cfg_din6766,
   output        cfg_din6767,
   output        cfg_din6768,
   output        cfg_din6769,
   output        cfg_din6770,
   output        cfg_din6771,
   output        cfg_din6772,
   output        cfg_din6773,
   output        cfg_din6774,
   output        cfg_din6775,
   output        cfg_din6776,
   output        cfg_din6777,
   output        cfg_din6778,
   output        cfg_din6779,
   output        cfg_din6780,
   output        cfg_din6781,
   output        cfg_din6782,
   output        cfg_din6783,
   output        cfg_din6784,
   output        cfg_din6785,
   output        cfg_din6786,
   output        cfg_din6787,
   output        cfg_din6788,
   output        cfg_din6789,
   output        cfg_din6790,
   output        cfg_din6791,
   output        cfg_din6792,
   output        cfg_din6793,
   output        cfg_din6794,
   output        cfg_din6795,
   output        cfg_din6796,
   output        cfg_din6797,
   output        cfg_din6798,
   output        cfg_din6799,
   output        cfg_din6800,
   output        cfg_din6801,
   output        cfg_din6802,
   output        cfg_din6803,
   output        cfg_din6804,
   output        cfg_din6805,
   output        cfg_din6806,
   output        cfg_din6807,
   output        cfg_din6808,
   output        cfg_din6809,
   output        cfg_din6810,
   output        cfg_din6811,
   output        cfg_din6812,
   output        cfg_din6813,
   output        cfg_din6814,
   output        cfg_din6815,
   output        cfg_din6816,
   output        cfg_din6817,
   output        cfg_din6818,
   output        cfg_din6819,
   output        cfg_din6820,
   output        cfg_din6821,
   output        cfg_din6822,
   output        cfg_din6823,
   output        cfg_din6824,
   output        cfg_din6825,
   output        cfg_din6826,
   output        cfg_din6827,
   output        cfg_din6828,
   output        cfg_din6829,
   output        cfg_din6830,
   output        cfg_din6831,
   output        cfg_din6832,
   output        cfg_din6833,
   output        cfg_din6834,
   output        cfg_din6835,
   output        cfg_din6836,
   output        cfg_din6837,
   output        cfg_din6838,
   output        cfg_din6839,
   output        cfg_din6840,
   output        cfg_din6841,
   output        cfg_din6842,
   output        cfg_din6843,
   output        cfg_din6844,
   output        cfg_din6845,
   output        cfg_din6846,
   output        cfg_din6847,
   output        cfg_din6848,
   output        cfg_din6849,
   output        cfg_din6850,
   output        cfg_din6851,
   output        cfg_din6852,
   output        cfg_din6853,
   output        cfg_din6854,
   output        cfg_din6855,
   output        cfg_din6856,
   output        cfg_din6857,
   output        cfg_din6858,
   output        cfg_din6859,
   output        cfg_din6860,
   output        cfg_din6861,
   output        cfg_din6862,
   output        cfg_din6863,
   output        cfg_din6864,
   output        cfg_din6865,
   output        cfg_din6866,
   output        cfg_din6867,
   output        cfg_din6868,
   output        cfg_din6869,
   output        cfg_din6870,
   output        cfg_din6871,
   output        cfg_din6872,
   output        cfg_din6873,
   output        cfg_din6874,
   output        cfg_din6875,
   output        cfg_din6876,
   output        cfg_din6877,
   output        cfg_din6878,
   output        cfg_din6879,
   output        cfg_din6880,
   output        cfg_din6881,
   output        cfg_din6882,
   output        cfg_din6883,
   output        cfg_din6884,
   output        cfg_din6885,
   output        cfg_din6886,
   output        cfg_din6887,
   output        cfg_din6888,
   output        cfg_din6889,
   output        cfg_din6890,
   output        cfg_din6891,
   output        cfg_din6892,
   output        cfg_din6893,
   output        cfg_din6894,
   output        cfg_din6895,
   output        cfg_din6896,
   output        cfg_din6897,
   output        cfg_din6898,
   output        cfg_din6899,
   output        cfg_din6900,
   output        cfg_din6901,
   output        cfg_din6902,
   output        cfg_din6903,
   output        cfg_din6904,
   output        cfg_din6905,
   output        cfg_din6906,
   output        cfg_din6907,
   output        cfg_din6908,
   output        cfg_din6909,
   output        cfg_din6910,
   output        cfg_din6911,
   output        cfg_din6912,
   output        cfg_din6913,
   output        cfg_din6914,
   output        cfg_din6915,
   output        cfg_din6916,
   output        cfg_din6917,
   output        cfg_din6918,
   output        cfg_din6919,
   output        cfg_din6920,
   output        cfg_din6921,
   output        cfg_din6922,
   output        cfg_din6923,
   output        cfg_din6924,
   output        cfg_din6925,
   output        cfg_din6926,
   output        cfg_din6927,
   output        cfg_din6928,
   output        cfg_din6929,
   output        cfg_din6930,
   output        cfg_din6931,
   output        cfg_din6932,
   output        cfg_din6933,
   output        cfg_din6934,
   output        cfg_din6935,
   output        cfg_din6936,
   output        cfg_din6937,
   output        cfg_din6938,
   output        cfg_din6939,
   output        cfg_din6940,
   output        cfg_din6941,
   output        cfg_din6942,
   output        cfg_din6943,
   output        cfg_din6944,
   output        cfg_din6945,
   output        cfg_din6946,
   output        cfg_din6947,
   output        cfg_din6948,
   output        cfg_din6949,
   output        cfg_din6950,
   output        cfg_din6951,
   output        cfg_din6952,
   output        cfg_din6953,
   output        cfg_din6954,
   output        cfg_din6955,
   output        cfg_din6956,
   output        cfg_din6957,
   output        cfg_din6958,
   output        cfg_din6959,
   output        cfg_din6960,
   output        cfg_din6961,
   output        cfg_din6962,
   output        cfg_din6963,
   output        cfg_din6964,
   output        cfg_din6965,
   output        cfg_din6966,
   output        cfg_din6967,
   output        cfg_din6968,
   output        cfg_din6969,
   output        cfg_din6970,
   output        cfg_din6971,
   output        cfg_din6972,
   output        cfg_din6973,
   output        cfg_din6974,
   output        cfg_din6975,
   output        cfg_din6976,
   output        cfg_din6977,
   output        cfg_din6978,
   output        cfg_din6979,
   output        cfg_din6980,
   output        cfg_din6981,
   output        cfg_din6982,
   output        cfg_din6983,
   output        cfg_din6984,
   output        cfg_din6985,
   output        cfg_din6986,
   output        cfg_din6987,
   output        cfg_din6988,
   output        cfg_din6989,
   output        cfg_din6990,
   output        cfg_din6991,
   output        cfg_din6992,
   output        cfg_din6993,
   output        cfg_din6994,
   output        cfg_din6995,
   output        cfg_din6996,
   output        cfg_din6997,
   output        cfg_din6998,
   output        cfg_din6999,
   output        cfg_din7000,
   output        cfg_din7001,
   output        cfg_din7002,
   output        cfg_din7003,
   output        cfg_din7004,
   output        cfg_din7005,
   output        cfg_din7006,
   output        cfg_din7007,
   output        cfg_din7008,
   output        cfg_din7009,
   output        cfg_din7010,
   output        cfg_din7011,
   output        cfg_din7012,
   output        cfg_din7013,
   output        cfg_din7014,
   output        cfg_din7015,
   output        cfg_din7016,
   output        cfg_din7017,
   output        cfg_din7018,
   output        cfg_din7019,
   output        cfg_din7020,
   output        cfg_din7021,
   output        cfg_din7022,
   output        cfg_din7023,
   output        cfg_din7024,
   output        cfg_din7025,
   output        cfg_din7026,
   output        cfg_din7027,
   output        cfg_din7028,
   output        cfg_din7029,
   output        cfg_din7030,
   output        cfg_din7031,
   output        cfg_din7032,
   output        cfg_din7033,
   output        cfg_din7034,
   output        cfg_din7035,
   output        cfg_din7036,
   output        cfg_din7037,
   output        cfg_din7038,
   output        cfg_din7039,
   output        cfg_din7040,
   output        cfg_din7041,
   output        cfg_din7042,
   output        cfg_din7043,
   output        cfg_din7044,
   output        cfg_din7045,
   output        cfg_din7046,
   output        cfg_din7047,
   output        cfg_din7048,
   output        cfg_din7049,
   output        cfg_din7050,
   output        cfg_din7051,
   output        cfg_din7052,
   output        cfg_din7053,
   output        cfg_din7054,
   output        cfg_din7055,
   output        cfg_din7056,
   output        cfg_din7057,
   output        cfg_din7058,
   output        cfg_din7059,
   output        cfg_din7060,
   output        cfg_din7061,
   output        cfg_din7062,
   output        cfg_din7063,
   output        cfg_din7064,
   output        cfg_din7065,
   output        cfg_din7066,
   output        cfg_din7067,
   output        cfg_din7068,
   output        cfg_din7069,
   output        cfg_din7070,
   output        cfg_din7071,
   output        cfg_din7072,
   output        cfg_din7073,
   output        cfg_din7074,
   output        cfg_din7075,
   output        cfg_din7076,
   output        cfg_din7077,
   output        cfg_din7078,
   output        cfg_din7079,
   output        cfg_din7080,
   output        cfg_din7081,
   output        cfg_din7082,
   output        cfg_din7083,
   output        cfg_din7084,
   output        cfg_din7085,
   output        cfg_din7086,
   output        cfg_din7087,
   output        cfg_din7088,
   output        cfg_din7089,
   output        cfg_din7090,
   output        cfg_din7091,
   output        cfg_din7092,
   output        cfg_din7093,
   output        cfg_din7094,
   output        cfg_din7095,
   output        cfg_din7096,
   output        cfg_din7097,
   output        cfg_din7098,
   output        cfg_din7099,
   output        cfg_din7100,
   output        cfg_din7101,
   output        cfg_din7102,
   output        cfg_din7103,
   output        cfg_din7104,
   output        cfg_din7105,
   output        cfg_din7106,
   output        cfg_din7107,
   output        cfg_din7108,
   output        cfg_din7109,
   output        cfg_din7110,
   output        cfg_din7111,
   output        cfg_din7112,
   output        cfg_din7113,
   output        cfg_din7114,
   output        cfg_din7115,
   output        cfg_din7116,
   output        cfg_din7117,
   output        cfg_din7118,
   output        cfg_din7119,
   output        cfg_din7120,
   output        cfg_din7121,
   output        cfg_din7122,
   output        cfg_din7123,
   output        cfg_din7124,
   output        cfg_din7125,
   output        cfg_din7126,
   output        cfg_din7127,
   output        cfg_din7128,
   output        cfg_din7129,
   output        cfg_din7130,
   output        cfg_din7131,
   output        cfg_din7132,
   output        cfg_din7133,
   output        cfg_din7134,
   output        cfg_din7135,
   output        cfg_din7136,
   output        cfg_din7137,
   output        cfg_din7138,
   output        cfg_din7139,
   output        cfg_din7140,
   output        cfg_din7141,
   output        cfg_din7142,
   output        cfg_din7143,
   output        cfg_din7144,
   output        cfg_din7145,
   output        cfg_din7146,
   output        cfg_din7147,
   output        cfg_din7148,
   output        cfg_din7149,
   output        cfg_din7150,
   output        cfg_din7151,
   output        cfg_din7152,
   output        cfg_din7153,
   output        cfg_din7154,
   output        cfg_din7155,
   output        cfg_din7156,
   output        cfg_din7157,
   output        cfg_din7158,
   output        cfg_din7159,
   output        cfg_din7160,
   output        cfg_din7161,
   output        cfg_din7162,
   output        cfg_din7163,
   output        cfg_din7164,
   output        cfg_din7165,
   output        cfg_din7166,
   output        cfg_din7167,
   output        cfg_din7168,
   output        cfg_din7169,
   output        cfg_din7170,
   output        cfg_din7171,
   output        cfg_din7172,
   output        cfg_din7173,
   output        cfg_din7174,
   output        cfg_din7175,
   output        cfg_din7176,
   output        cfg_din7177,
   output        cfg_din7178,
   output        cfg_din7179,
   output        cfg_din7180,
   output        cfg_din7181,
   output        cfg_din7182,
   output        cfg_din7183,
   output        cfg_din7184,
   output        cfg_din7185,
   output        cfg_din7186,
   output        cfg_din7187,
   output        cfg_din7188,
   output        cfg_din7189,
   output        cfg_din7190,
   output        cfg_din7191,
   output        cfg_din7192,
   output        cfg_din7193,
   output        cfg_din7194,
   output        cfg_din7195,
   output        cfg_din7196,
   output        cfg_din7197,
   output        cfg_din7198,
   output        cfg_din7199,
   output        cfg_din7200,
   output        cfg_din7201,
   output        cfg_din7202,
   output        cfg_din7203,
   output        cfg_din7204,
   output        cfg_din7205,
   output        cfg_din7206,
   output        cfg_din7207,
   output        cfg_din7208,
   output        cfg_din7209,
   output        cfg_din7210,
   output        cfg_din7211,
   output        cfg_din7212,
   output        cfg_din7213,
   output        cfg_din7214,
   output        cfg_din7215,
   output        cfg_din7216,
   output        cfg_din7217,
   output        cfg_din7218,
   output        cfg_din7219,
   output        cfg_din7220,
   output        cfg_din7221,
   output        cfg_din7222,
   output        cfg_din7223,
   output        cfg_din7224,
   output        cfg_din7225,
   output        cfg_din7226,
   output        cfg_din7227,
   output        cfg_din7228,
   output        cfg_din7229,
   output        cfg_din7230,
   output        cfg_din7231,
   output        cfg_din7232,
   output        cfg_din7233,
   output        cfg_din7234,
   output        cfg_din7235,
   output        cfg_din7236,
   output        cfg_din7237,
   output        cfg_din7238,
   output        cfg_din7239,
   output        cfg_din7240,
   output        cfg_din7241,
   output        cfg_din7242,
   output        cfg_din7243,
   output        cfg_din7244,
   output        cfg_din7245,
   output        cfg_din7246,
   output        cfg_din7247,
   output        cfg_din7248,
   output        cfg_din7249,
   output        cfg_din7250,
   output        cfg_din7251,
   output        cfg_din7252,
   output        cfg_din7253,
   output        cfg_din7254,
   output        cfg_din7255,
   output        cfg_din7256,
   output        cfg_din7257,
   output        cfg_din7258,
   output        cfg_din7259,
   output        cfg_din7260,
   output        cfg_din7261,
   output        cfg_din7262,
   output        cfg_din7263,
   output        cfg_din7264,
   output        cfg_din7265,
   output        cfg_din7266,
   output        cfg_din7267,
   output        cfg_din7268,
   output        cfg_din7269,
   output        cfg_din7270,
   output        cfg_din7271,
   output        cfg_din7272,
   output        cfg_din7273,
   output        cfg_din7274,
   output        cfg_din7275,
   output        cfg_din7276,
   output        cfg_din7277,
   output        cfg_din7278,
   output        cfg_din7279,
   output        cfg_din7280,
   output        cfg_din7281,
   output        cfg_din7282,
   output        cfg_din7283,
   output        cfg_din7284,
   output        cfg_din7285,
   output        cfg_din7286,
   output        cfg_din7287,
   output        cfg_din7288,
   output        cfg_din7289,
   output        cfg_din7290,
   output        cfg_din7291,
   output        cfg_din7292,
   output        cfg_din7293,
   output        cfg_din7294,
   output        cfg_din7295,
   output        cfg_din7296,
   output        cfg_din7297,
   output        cfg_din7298,
   output        cfg_din7299,
   output        cfg_din7300,
   output        cfg_din7301,
   output        cfg_din7302,
   output        cfg_din7303,
   output        cfg_din7304,
   output        cfg_din7305,
   output        cfg_din7306,
   output        cfg_din7307,
   output        cfg_din7308,
   output        cfg_din7309,
   output        cfg_din7310,
   output        cfg_din7311,
   output        cfg_din7312,
   output        cfg_din7313,
   output        cfg_din7314,
   output        cfg_din7315,
   output        cfg_din7316,
   output        cfg_din7317,
   output        cfg_din7318,
   output        cfg_din7319,
   output        cfg_din7320,
   output        cfg_din7321,
   output        cfg_din7322,
   output        cfg_din7323,
   output        cfg_din7324,
   output        cfg_din7325,
   output        cfg_din7326,
   output        cfg_din7327,
   output        cfg_din7328,
   output        cfg_din7329,
   output        cfg_din7330,
   output        cfg_din7331,
   output        cfg_din7332,
   output        cfg_din7333,
   output        cfg_din7334,
   output        cfg_din7335,
   output        cfg_din7336,
   output        cfg_din7337,
   output        cfg_din7338,
   output        cfg_din7339,
   output        cfg_din7340,
   output        cfg_din7341,
   output        cfg_din7342,
   output        cfg_din7343,
   output        cfg_din7344,
   output        cfg_din7345,
   output        cfg_din7346,
   output        cfg_din7347,
   output        cfg_din7348,
   output        cfg_din7349,
   output        cfg_din7350,
   output        cfg_din7351,
   output        cfg_din7352,
   output        cfg_din7353,
   output        cfg_din7354,
   output        cfg_din7355,
   output        cfg_din7356,
   output        cfg_din7357,
   output        cfg_din7358,
   output        cfg_din7359,
   output        cfg_din7360,
   output        cfg_din7361,
   output        cfg_din7362,
   output        cfg_din7363,
   output        cfg_din7364,
   output        cfg_din7365,
   output        cfg_din7366,
   output        cfg_din7367,
   output        cfg_din7368,
   output        cfg_din7369,
   output        cfg_din7370,
   output        cfg_din7371,
   output        cfg_din7372,
   output        cfg_din7373,
   output        cfg_din7374,
   output        cfg_din7375,
   output        cfg_din7376,
   output        cfg_din7377,
   output        cfg_din7378,
   output        cfg_din7379,
   output        cfg_din7380,
   output        cfg_din7381,
   output        cfg_din7382,
   output        cfg_din7383,
   output        cfg_din7384,
   output        cfg_din7385,
   output        cfg_din7386,
   output        cfg_din7387,
   output        cfg_din7388,
   output        cfg_din7389,
   output        cfg_din7390,
   output        cfg_din7391,
   output        cfg_din7392,
   output        cfg_din7393,
   output        cfg_din7394,
   output        cfg_din7395,
   output        cfg_din7396,
   output        cfg_din7397,
   output        cfg_din7398,
   output        cfg_din7399,
   output        cfg_din7400,
   output        cfg_din7401,
   output        cfg_din7402,
   output        cfg_din7403,
   output        cfg_din7404,
   output        cfg_din7405,
   output        cfg_din7406,
   output        cfg_din7407,
   output        cfg_din7408,
   output        cfg_din7409,
   output        cfg_din7410,
   output        cfg_din7411,
   output        cfg_din7412,
   output        cfg_din7413,
   output        cfg_din7414,
   output        cfg_din7415,
   output        cfg_din7416,
   output        cfg_din7417,
   output        cfg_din7418,
   output        cfg_din7419,
   output        cfg_din7420,
   output        cfg_din7421,
   output        cfg_din7422,
   output        cfg_din7423,
   output        cfg_din7424,
   output        cfg_din7425,
   output        cfg_din7426,
   output        cfg_din7427,
   output        cfg_din7428,
   output        cfg_din7429,
   output        cfg_din7430,
   output        cfg_din7431,
   output        cfg_din7432,
   output        cfg_din7433,
   output        cfg_din7434,
   output        cfg_din7435,
   output        cfg_din7436,
   output        cfg_din7437,
   output        cfg_din7438,
   output        cfg_din7439,
   output        cfg_din7440,
   output        cfg_din7441,
   output        cfg_din7442,
   output        cfg_din7443,
   output        cfg_din7444,
   output        cfg_din7445,
   output        cfg_din7446,
   output        cfg_din7447,
   output        cfg_din7448,
   output        cfg_din7449,
   output        cfg_din7450,
   output        cfg_din7451,
   output        cfg_din7452,
   output        cfg_din7453,
   output        cfg_din7454,
   output        cfg_din7455,
   output        cfg_din7456,
   output        cfg_din7457,
   output        cfg_din7458,
   output        cfg_din7459,
   output        cfg_din7460,
   output        cfg_din7461,
   output        cfg_din7462,
   output        cfg_din7463,
   output        cfg_din7464,
   output        cfg_din7465,
   output        cfg_din7466,
   output        cfg_din7467,
   output        cfg_din7468,
   output        cfg_din7469,
   output        cfg_din7470,
   output        cfg_din7471,
   output        cfg_din7472,
   output        cfg_din7473,
   output        cfg_din7474,
   output        cfg_din7475,
   output        cfg_din7476,
   output        cfg_din7477,
   output        cfg_din7478,
   output        cfg_din7479,
   output        cfg_din7480,
   output        cfg_din7481,
   output        cfg_din7482,
   output        cfg_din7483,
   output        cfg_din7484,
   output        cfg_din7485,
   output        cfg_din7486,
   output        cfg_din7487,
   output        cfg_din7488,
   output        cfg_din7489,
   output        cfg_din7490,
   output        cfg_din7491,
   output        cfg_din7492,
   output        cfg_din7493,
   output        cfg_din7494,
   output        cfg_din7495,
   output        cfg_din7496,
   output        cfg_din7497,
   output        cfg_din7498,
   output        cfg_din7499,
   output        cfg_din7500,
   output        cfg_din7501,
   output        cfg_din7502,
   output        cfg_din7503,
   output        cfg_din7504,
   output        cfg_din7505,
   output        cfg_din7506,
   output        cfg_din7507,
   output        cfg_din7508,
   output        cfg_din7509,
   output        cfg_din7510,
   output        cfg_din7511,
   output        cfg_din7512,
   output        cfg_din7513,
   output        cfg_din7514,
   output        cfg_din7515,
   output        cfg_din7516,
   output        cfg_din7517,
   output        cfg_din7518,
   output        cfg_din7519,
   output        cfg_din7520,
   output        cfg_din7521,
   output        cfg_din7522,
   output        cfg_din7523,
   output        cfg_din7524,
   output        cfg_din7525,
   output        cfg_din7526,
   output        cfg_din7527,
   output        cfg_din7528,
   output        cfg_din7529,
   output        cfg_din7530,
   output        cfg_din7531,
   output        cfg_din7532,
   output        cfg_din7533,
   output        cfg_din7534,
   output        cfg_din7535,
   output        cfg_din7536,
   output        cfg_din7537,
   output        cfg_din7538,
   output        cfg_din7539,
   output        cfg_din7540,
   output        cfg_din7541,
   output        cfg_din7542,
   output        cfg_din7543,
   output        cfg_din7544,
   output        cfg_din7545,
   output        cfg_din7546,
   output        cfg_din7547,
   output        cfg_din7548,
   output        cfg_din7549,
   output        cfg_din7550,
   output        cfg_din7551,
   output        cfg_din7552,
   output        cfg_din7553,
   output        cfg_din7554,
   output        cfg_din7555,
   output        cfg_din7556,
   output        cfg_din7557,
   output        cfg_din7558,
   output        cfg_din7559,
   output        cfg_din7560,
   output        cfg_din7561,
   output        cfg_din7562,
   output        cfg_din7563,
   output        cfg_din7564,
   output        cfg_din7565,
   output        cfg_din7566,
   output        cfg_din7567,
   output        cfg_din7568,
   output        cfg_din7569,
   output        cfg_din7570,
   output        cfg_din7571,
   output        cfg_din7572,
   output        cfg_din7573,
   output        cfg_din7574,
   output        cfg_din7575,
   output        cfg_din7576,
   output        cfg_din7577,
   output        cfg_din7578,
   output        cfg_din7579,
   output        cfg_din7580,
   output        cfg_din7581,
   output        cfg_din7582,
   output        cfg_din7583,
   output        cfg_din7584,
   output        cfg_din7585,
   output        cfg_din7586,
   output        cfg_din7587,
   output        cfg_din7588,
   output        cfg_din7589,
   output        cfg_din7590,
   output        cfg_din7591,
   output        cfg_din7592,
   output        cfg_din7593,
   output        cfg_din7594,
   output        cfg_din7595,
   output        cfg_din7596,
   output        cfg_din7597,
   output        cfg_din7598,
   output        cfg_din7599,
   output        cfg_din7600,
   output        cfg_din7601,
   output        cfg_din7602,
   output        cfg_din7603,
   output        cfg_din7604,
   output        cfg_din7605,
   output        cfg_din7606,
   output        cfg_din7607,
   output        cfg_din7608,
   output        cfg_din7609,
   output        cfg_din7610,
   output        cfg_din7611,
   output        cfg_din7612,
   output        cfg_din7613,
   output        cfg_din7614,
   output        cfg_din7615,
   output        cfg_din7616,
   output        cfg_din7617,
   output        cfg_din7618,
   output        cfg_din7619,
   output        cfg_din7620,
   output        cfg_din7621,
   output        cfg_din7622,
   output        cfg_din7623,
   output        cfg_din7624,
   output        cfg_din7625,
   output        cfg_din7626,
   output        cfg_din7627,
   output        cfg_din7628,
   output        cfg_din7629,
   output        cfg_din7630,
   output        cfg_din7631,
   output        cfg_din7632,
   output        cfg_din7633,
   output        cfg_din7634,
   output        cfg_din7635,
   output        cfg_din7636,
   output        cfg_din7637,
   output        cfg_din7638,
   output        cfg_din7639,
   output        cfg_din7640,
   output        cfg_din7641,
   output        cfg_din7642,
   output        cfg_din7643,
   output        cfg_din7644,
   output        cfg_din7645,
   output        cfg_din7646,
   output        cfg_din7647,
   output        cfg_din7648,
   output        cfg_din7649,
   output        cfg_din7650,
   output        cfg_din7651,
   output        cfg_din7652,
   output        cfg_din7653,
   output        cfg_din7654,
   output        cfg_din7655,
   output        cfg_din7656,
   output        cfg_din7657,
   output        cfg_din7658,
   output        cfg_din7659,
   output        cfg_din7660,
   output        cfg_din7661,
   output        cfg_din7662,
   output        cfg_din7663,
   output        cfg_din7664,
   output        cfg_din7665,
   output        cfg_din7666,
   output        cfg_din7667,
   output        cfg_din7668,
   output        cfg_din7669,
   output        cfg_din7670,
   output        cfg_din7671,
   output        cfg_din7672,
   output        cfg_din7673,
   output        cfg_din7674,
   output        cfg_din7675,
   output        cfg_din7676,
   output        cfg_din7677,
   output        cfg_din7678,
   output        cfg_din7679,
   output        cfg_din7680,
   output        cfg_din7681,
   output        cfg_din7682,
   output        cfg_din7683,
   output        cfg_din7684,
   output        cfg_din7685,
   output        cfg_din7686,
   output        cfg_din7687,
   output        cfg_din7688,
   output        cfg_din7689,
   output        cfg_din7690,
   output        cfg_din7691,
   output        cfg_din7692,
   output        cfg_din7693,
   output        cfg_din7694,
   output        cfg_din7695,
   output        cfg_din7696,
   output        cfg_din7697,
   output        cfg_din7698,
   output        cfg_din7699,
   output        cfg_din7700,
   output        cfg_din7701,
   output        cfg_din7702,
   output        cfg_din7703,
   output        cfg_din7704,
   output        cfg_din7705,
   output        cfg_din7706,
   output        cfg_din7707,
   output        cfg_din7708,
   output        cfg_din7709,
   output        cfg_din7710,
   output        cfg_din7711,
   output        cfg_din7712,
   output        cfg_din7713,
   output        cfg_din7714,
   output        cfg_din7715,
   output        cfg_din7716,
   output        cfg_din7717,
   output        cfg_din7718,
   output        cfg_din7719,
   output        cfg_din7720,
   output        cfg_din7721,
   output        cfg_din7722,
   output        cfg_din7723,
   output        cfg_din7724,
   output        cfg_din7725,
   output        cfg_din7726,
   output        cfg_din7727,
   output        cfg_din7728,
   output        cfg_din7729,
   output        cfg_din7730,
   output        cfg_din7731,
   output        cfg_din7732,
   output        cfg_din7733,
   output        cfg_din7734,
   output        cfg_din7735,
   output        cfg_din7736,
   output        cfg_din7737,
   output        cfg_din7738,
   output        cfg_din7739,
   output        cfg_din7740,
   output        cfg_din7741,
   output        cfg_din7742,
   output        cfg_din7743,
   output        cfg_din7744,
   output        cfg_din7745,
   output        cfg_din7746,
   output        cfg_din7747,
   output        cfg_din7748,
   output        cfg_din7749,
   output        cfg_din7750,
   output        cfg_din7751,
   output        cfg_din7752,
   output        cfg_din7753,
   output        cfg_din7754,
   output        cfg_din7755,
   output        cfg_din7756,
   output        cfg_din7757,
   output        cfg_din7758,
   output        cfg_din7759,
   output        cfg_din7760,
   output        cfg_din7761,
   output        cfg_din7762,
   output        cfg_din7763,
   output        cfg_din7764,
   output        cfg_din7765,
   output        cfg_din7766,
   output        cfg_din7767,
   output        cfg_din7768,
   output        cfg_din7769,
   output        cfg_din7770,
   output        cfg_din7771,
   output        cfg_din7772,
   output        cfg_din7773,
   output        cfg_din7774,
   output        cfg_din7775,
   output        cfg_din7776,
   output        cfg_din7777,
   output        cfg_din7778,
   output        cfg_din7779,
   output        cfg_din7780,
   output        cfg_din7781,
   output        cfg_din7782,
   output        cfg_din7783,
   output        cfg_din7784,
   output        cfg_din7785,
   output        cfg_din7786,
   output        cfg_din7787,
   output        cfg_din7788,
   output        cfg_din7789,
   output        cfg_din7790,
   output        cfg_din7791,
   output        cfg_din7792,
   output        cfg_din7793,
   output        cfg_din7794,
   output        cfg_din7795,
   output        cfg_din7796,
   output        cfg_din7797,
   output        cfg_din7798,
   output        cfg_din7799,
   output        cfg_din7800,
   output        cfg_din7801,
   output        cfg_din7802,
   output        cfg_din7803,
   output        cfg_din7804,
   output        cfg_din7805,
   output        cfg_din7806,
   output        cfg_din7807,
   output        cfg_din7808,
   output        cfg_din7809,
   output        cfg_din7810,
   output        cfg_din7811,
   output        cfg_din7812,
   output        cfg_din7813,
   output        cfg_din7814,
   output        cfg_din7815,
   output        cfg_din7816,
   output        cfg_din7817,
   output        cfg_din7818,
   output        cfg_din7819,
   output        cfg_din7820,
   output        cfg_din7821,
   output        cfg_din7822,
   output        cfg_din7823,
   output        cfg_din7824,
   output        cfg_din7825,
   output        cfg_din7826,
   output        cfg_din7827,
   output        cfg_din7828,
   output        cfg_din7829,
   output        cfg_din7830,
   output        cfg_din7831,
   output        cfg_din7832,
   output        cfg_din7833,
   output        cfg_din7834,
   output        cfg_din7835,
   output        cfg_din7836,
   output        cfg_din7837,
   output        cfg_din7838,
   output        cfg_din7839,
   output        cfg_din7840,
   output        cfg_din7841,
   output        cfg_din7842,
   output        cfg_din7843,
   output        cfg_din7844,
   output        cfg_din7845,
   output        cfg_din7846,
   output        cfg_din7847,
   output        cfg_din7848,
   output        cfg_din7849,
   output        cfg_din7850,
   output        cfg_din7851,
   output        cfg_din7852,
   output        cfg_din7853,
   output        cfg_din7854,
   output        cfg_din7855,
   output        cfg_din7856,
   output        cfg_din7857,
   output        cfg_din7858,
   output        cfg_din7859,
   output        cfg_din7860,
   output        cfg_din7861,
   output        cfg_din7862,
   output        cfg_din7863,
   output        cfg_din7864,
   output        cfg_din7865,
   output        cfg_din7866,
   output        cfg_din7867,
   output        cfg_din7868,
   output        cfg_din7869,
   output        cfg_din7870,
   output        cfg_din7871,
   output        cfg_din7872,
   output        cfg_din7873,
   output        cfg_din7874,
   output        cfg_din7875,
   output        cfg_din7876,
   output        cfg_din7877,
   output        cfg_din7878,
   output        cfg_din7879,
   output        cfg_din7880,
   output        cfg_din7881,
   output        cfg_din7882,
   output        cfg_din7883,
   output        cfg_din7884,
   output        cfg_din7885,
   output        cfg_din7886,
   output        cfg_din7887,
   output        cfg_din7888,
   output        cfg_din7889,
   output        cfg_din7890,
   output        cfg_din7891,
   output        cfg_din7892,
   output        cfg_din7893,
   output        cfg_din7894,
   output        cfg_din7895,
   output        cfg_din7896,
   output        cfg_din7897,
   output        cfg_din7898,
   output        cfg_din7899,
   output        cfg_din7900,
   output        cfg_din7901,
   output        cfg_din7902,
   output        cfg_din7903,
   output        cfg_din7904,
   output        cfg_din7905,
   output        cfg_din7906,
   output        cfg_din7907,
   output        cfg_din7908,
   output        cfg_din7909,
   output        cfg_din7910,
   output        cfg_din7911,
   output        cfg_din7912,
   output        cfg_din7913,
   output        cfg_din7914,
   output        cfg_din7915,
   output        cfg_din7916,
   output        cfg_din7917,
   output        cfg_din7918,
   output        cfg_din7919,
   output        cfg_din7920,
   output        cfg_din7921,
   output        cfg_din7922,
   output        cfg_din7923,
   output        cfg_din7924,
   output        cfg_din7925,
   output        cfg_din7926,
   output        cfg_din7927,
   output        cfg_din7928,
   output        cfg_din7929,
   output        cfg_din7930,
   output        cfg_din7931,
   output        cfg_din7932,
   output        cfg_din7933,
   output        cfg_din7934,
   output        cfg_din7935,
   output        cfg_din7936,
   output        cfg_din7937,
   output        cfg_din7938,
   output        cfg_din7939,
   output        cfg_din7940,
   output        cfg_din7941,
   output        cfg_din7942,
   output        cfg_din7943,
   output        cfg_din7944,
   output        cfg_din7945,
   output        cfg_din7946,
   output        cfg_din7947,
   output        cfg_din7948,
   output        cfg_din7949,
   output        cfg_din7950,
   output        cfg_din7951,
   output        cfg_din7952,
   output        cfg_din7953,
   output        cfg_din7954,
   output        cfg_din7955,
   output        cfg_din7956,
   output        cfg_din7957,
   output        cfg_din7958,
   output        cfg_din7959,
   output        cfg_din7960,
   output        cfg_din7961,
   output        cfg_din7962,
   output        cfg_din7963,
   output        cfg_din7964,
   output        cfg_din7965,
   output        cfg_din7966,
   output        cfg_din7967,
   output        cfg_din7968,
   output        cfg_din7969,
   output        cfg_din7970,
   output        cfg_din7971,
   output        cfg_din7972,
   output        cfg_din7973,
   output        cfg_din7974,
   output        cfg_din7975,
   output        cfg_din7976,
   output        cfg_din7977,
   output        cfg_din7978,
   output        cfg_din7979,
   output        cfg_din7980,
   output        cfg_din7981,
   output        cfg_din7982,
   output        cfg_din7983,
   output        cfg_din7984,
   output        cfg_din7985,
   output        cfg_din7986,
   output        cfg_din7987,
   output        cfg_din7988,
   output        cfg_din7989,
   output        cfg_din7990,
   output        cfg_din7991,
   output        cfg_din7992,
   output        cfg_din7993,
   output        cfg_din7994,
   output        cfg_din7995,
   output        cfg_din7996,
   output        cfg_din7997,
   output        cfg_din7998,
   output        cfg_din7999,
   output        cfg_din8000,
   output        cfg_din8001,
   output        cfg_din8002,
   output        cfg_din8003,
   output        cfg_din8004,
   output        cfg_din8005,
   output        cfg_din8006,
   output        cfg_din8007,
   output        cfg_din8008,
   output        cfg_din8009,
   output        cfg_din8010,
   output        cfg_din8011,
   output        cfg_din8012,
   output        cfg_din8013,
   output        cfg_din8014,
   output        cfg_din8015,
   output        cfg_din8016,
   output        cfg_din8017,
   output        cfg_din8018,
   output        cfg_din8019,
   output        cfg_din8020,
   output        cfg_din8021,
   output        cfg_din8022,
   output        cfg_din8023,
   output        cfg_din8024,
   output        cfg_din8025,
   output        cfg_din8026,
   output        cfg_din8027,
   output        cfg_din8028,
   output        cfg_din8029,
   output        cfg_din8030,
   output        cfg_din8031,
   output        cfg_din8032,
   output        cfg_din8033,
   output        cfg_din8034,
   output        cfg_din8035,
   output        cfg_din8036,
   output        cfg_din8037,
   output        cfg_din8038,
   output        cfg_din8039,
   output        cfg_din8040,
   output        cfg_din8041,
   output        cfg_din8042,
   output        cfg_din8043,
   output        cfg_din8044,
   output        cfg_din8045,
   output        cfg_din8046,
   output        cfg_din8047,
   output        cfg_din8048,
   output        cfg_din8049,
   output        cfg_din8050,
   output        cfg_din8051,
   output        cfg_din8052,
   output        cfg_din8053,
   output        cfg_din8054,
   output        cfg_din8055,
   output        cfg_din8056,
   output        cfg_din8057,
   output        cfg_din8058,
   output        cfg_din8059,
   output        cfg_din8060,
   output        cfg_din8061,
   output        cfg_din8062,
   output        cfg_din8063,
   output        cfg_din8064,
   output        cfg_din8065,
   output        cfg_din8066,
   output        cfg_din8067,
   output        cfg_din8068,
   output        cfg_din8069,
   output        cfg_din8070,
   output        cfg_din8071,
   output        cfg_din8072,
   output        cfg_din8073,
   output        cfg_din8074,
   output        cfg_din8075,
   output        cfg_din8076,
   output        cfg_din8077,
   output        cfg_din8078,
   output        cfg_din8079,
   output        cfg_din8080,
   output        cfg_din8081,
   output        cfg_din8082,
   output        cfg_din8083,
   output        cfg_din8084,
   output        cfg_din8085,
   output        cfg_din8086,
   output        cfg_din8087,
   output        cfg_din8088,
   output        cfg_din8089,
   output        cfg_din8090,
   output        cfg_din8091,
   output        cfg_din8092,
   output        cfg_din8093,
   output        cfg_din8094,
   output        cfg_din8095,
   output        cfg_din8096,
   output        cfg_din8097,
   output        cfg_din8098,
   output        cfg_din8099,
   output        cfg_din8100,
   output        cfg_din8101,
   output        cfg_din8102,
   output        cfg_din8103,
   output        cfg_din8104,
   output        cfg_din8105,
   output        cfg_din8106,
   output        cfg_din8107,
   output        cfg_din8108,
   output        cfg_din8109,
   output        cfg_din8110,
   output        cfg_din8111,
   output        cfg_din8112,
   output        cfg_din8113,
   output        cfg_din8114,
   output        cfg_din8115,
   output        cfg_din8116,
   output        cfg_din8117,
   output        cfg_din8118,
   output        cfg_din8119,
   output        cfg_din8120,
   output        cfg_din8121,
   output        cfg_din8122,
   output        cfg_din8123,
   output        cfg_din8124,
   output        cfg_din8125,
   output        cfg_din8126,
   output        cfg_din8127,
   output        cfg_din8128,
   output        cfg_din8129,
   output        cfg_din8130,
   output        cfg_din8131,
   output        cfg_din8132,
   output        cfg_din8133,
   output        cfg_din8134,
   output        cfg_din8135,
   output        cfg_din8136,
   output        cfg_din8137,
   output        cfg_din8138,
   output        cfg_din8139,
   output        cfg_din8140,
   output        cfg_din8141,
   output        cfg_din8142,
   output        cfg_din8143,
   output        cfg_din8144,
   output        cfg_din8145,
   output        cfg_din8146,
   output        cfg_din8147,
   output        cfg_din8148,
   output        cfg_din8149,
   output        cfg_din8150,
   output        cfg_din8151,
   output        cfg_din8152,
   output        cfg_din8153,
   output        cfg_din8154,
   output        cfg_din8155,
   output        cfg_din8156,
   output        cfg_din8157,
   output        cfg_din8158,
   output        cfg_din8159,
   output        cfg_din8160,
   output        cfg_din8161,
   output        cfg_din8162,
   output        cfg_din8163,
   output        cfg_din8164,
   output        cfg_din8165,
   output        cfg_din8166,
   output        cfg_din8167,
   output        cfg_din8168,
   output        cfg_din8169,
   output        cfg_din8170,
   output        cfg_din8171,
   output        cfg_din8172,
   output        cfg_din8173,
   output        cfg_din8174,
   output        cfg_din8175,
   output        cfg_din8176,
   output        cfg_din8177,
   output        cfg_din8178,
   output        cfg_din8179,
   output        cfg_din8180,
   output        cfg_din8181,
   output        cfg_din8182,
   output        cfg_din8183,
   output        cfg_din8184,
   output        cfg_din8185,
   output        cfg_din8186,
   output        cfg_din8187,
   output        cfg_din8188,
   output        cfg_din8189,
   output        cfg_din8190,
   output        cfg_din8191,
   output        tc_cfg_din,
   output        cc_cfg_din0,
   output        cc_cfg_din1,
   output        cc_cfg_din2,
   output        cc_cfg_din3,

