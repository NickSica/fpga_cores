    .INIT_00(256'h0207c40b00201f01001100202af2ff00001020202a601f000250003640e28000),
    .INIT_01(256'h00bc0c0b0020100100bd0d202b82003300be0e3240b2800000bf0f1d0022df02),
    .INIT_02(256'h0010802076c2df020207f5202c101f000250003240b320770207f21d00320566),
    .INIT_03(256'h001100010822202a0010002f01f2202a0207c42243c2202a0011010100228000),
    .INIT_04(256'h0250003242d2202a0207091d0022202a0207f22200a2202a0207e22057c2202a),
    .INIT_05(256'h0011013242d2202a0010801d0102202a0207a63242d2202a0207f81d0082202a),
    .INIT_06(256'h0207e2050402202a001100205512202a0010043641f2202a0207c41d0202202a),
    .INIT_07(256'h0207fb1d040280000250002243c2df020207150100201f010207f22055a2202a),
    .INIT_08(256'h0207c42055a1d004001101030bf32077001080205511d0010207ac3642620554),
    .INIT_09(256'h0207f23602a205570207e21d080323a10011002243c1d00800100801002322ca),
    .INIT_0A(256'h0207b6010022055a0207fe2055a01060025000030bf322ca020726205511d004),
    .INIT_0B(256'h00100c0b002205280207c4202802052000110120277205660010802243c0109f),
    .INIT_0C(256'h02073b0b002200370207f22028922bfc0207e232437204f20011001d00220538),
    .INIT_0D(256'h0368352076c0900200d008202922500000900e32437200630250001d0032004a),
    .INIT_0E(256'h032839010000d00100d0022055a0b00000900e0504032046025000205510d080),
    .INIT_0F(256'h03283d0900d0121f00d0022200a011ff00900f20594010ff0250002056636046),
    .INIT_10(256'h0328410900d3e04000d002250001b2000090103643f1b1000250000d08019001),
    .INIT_11(256'h032845014400d04000d0022500009001009011364432f0000250000d04001001),
    .INIT_12(256'h00100c0b0142b00c0008400b2152b00000095001300250000250000150a32046),
    .INIT_13(256'h0131000d0082d01001480814300010ff01490e142002bfff0011000d0102bf7e),
    .INIT_14(256'h036857011012d00101d100030070300f03684d1430009001019001142002d011),
    .INIT_15(256'h00d508224540900602500014106360590018ff3a4580d0200019ff190010900d),
    .INIT_16(256'h0018ff2d2090900d0019ff2d30a09006001102123500900603685d1024022054),
    .INIT_17(256'h00015001a002205b03e86a250000900701d1030201036060025000090080d080),
    .INIT_18(256'h01410e09c1c2053601180114b06250000018ff14b06090070000400bb1309007),
    .INIT_19(256'h00190b10ba02053a01180809f1f204f603e86209e1e2052a01400809d1d2051a),
    .INIT_1A(256'h00084013f002051200095013e002053402500013d002053800110410cb020528),
    .INIT_1B(256'h0011022043f204f603e87320489204fc01b90501b002053c01981801a04204f6),
    .INIT_1C(256'h0001802043f0101902500009d07250000018ff2043f204f20019ff09c07204fa),
    .INIT_1D(256'h01410601a732021f01490009f07250000141062043f3e07400381f09e0719001),
    .INIT_1E(256'h0011020b6120d0010149000b5110900d0141060b4102020d01490001b0120227),
    .INIT_1F(256'h01400612e600108001400612d50206b7000a9010c40206b0000080036013207a),
    .INIT_20(256'h0140063e47d1dc93014a001bb00207ef01400619a01207c401400613f0001101),
    .INIT_21(256'h01d90b20489207db03d00001b010100001da5d01a7401100014a00250003607d),
    .INIT_22(256'h001104204431d11203a88d2df070311e01d81420443001e003688b2500020890),
    .INIT_23(256'h025000204431d11603a88b2dd07320a201d808204431d1140250002de0732092),
    .INIT_24(256'h009508204432f23902f5032db0701220009508204432202a0208a42dc07320b0),
    .INIT_25(256'h009508015001400802f6050146c1410a02f50425000001e00096082da07000d0),
    .INIT_26(256'h0095080d0101d04802f6310b014320be02f5300b2151d05800960801300030f8),
    .INIT_27(256'h009508142001d0b802f6380d008320c102f537143001d08800960814200320be),
    .INIT_28(256'h025000190012f23902f606011010122002f53c030072202a00960814300320c1),
    .INIT_29(256'h02d5091024014008001100224a31410a00160714106001e00015ef3a4a7000d0),
    .INIT_2A(256'h001300090081d0880250002d209320c102d10b2d30a1d04802d60a12350030f8),
    .INIT_2B(256'h02f0162d0082202a0208c82d209320c400b1172d30a1d0b800b01606010320c4),
    .INIT_2C(256'h00b01814c00001e000130114b00000d002f22014a062f23902f1172500001230),
    .INIT_2D(256'h02f119250001d08802f01814f00030f80208c814e001400800b11914d001410a),
    .INIT_2E(256'h00b11b14c081d0e800b01a14d08320c100130214e081d0c802f22114f0e320be),
    .INIT_2F(256'h02f222110b92f00202f11b250000100202f01a14a082202a0208c814b08320c1),
    .INIT_30(256'h0208c819011220c600b11d390002f00200b01c190e90100300130339000220c6),
    .INIT_31(256'h025000190f60120302f223390002020902f11d110072f00202f01c3e4c901004),
    .INIT_32(256'h03100000c000100101f1ff250002f03a01d0ff1100a01000001200250002f201),
    .INIT_33(256'h014006204d32024d0140062054620244014006204dd20219014006204d32f024),
    .INIT_34(256'h01400e01100207ef014100250002026c014006205462023b014100204dd20232),
    .INIT_35(256'h00b224141002026c01003014c06207db01400e141000101001400e14c0601100),
    .INIT_36(256'h022bfc1410001100022bfc14c0620256022bfc141000110002500014c0601010),
    .INIT_37(256'h022bfc11107206b0022bfc3a4e020798022bfc1d10a207db022bfc2500001010),
    .INIT_38(256'h022bfc2054901101022bfc01a0001080022bfc25000206b0022bfc1113020766),
    .INIT_39(256'h022bfc0110401004022bfc3900001100022bfc204bf207ef022bfc09006207c4),
    .INIT_3A(256'h022bfc04a00207a6022bfc364e820232022bfc19101207a6022bfc204b1207db),
    .INIT_3B(256'h022bfc19201207a6022bfc2054620244022bfc204dd207a6022bfc001002023b),
    .INIT_3C(256'h022bfc22546206b0022bfc0110d20766022bfc25000206b0022bfc364e32024d),
    .INIT_3D(256'h022bfc2254601014022bfc0115f01100022bfc22546207ef022bfc011202026c),
    .INIT_3E(256'h022bfc22546207c4022bfc0113101101022bfc22546010c0022bfc0113e207db),
    .INIT_3F(256'h022bfc2254620256022bfc0113001100022bfc2254601014022bfc01133207a6),
    .INIT_40(256'h022bfc225460b002022bfc01132207db022bfc2254601014022bfc0113101100),
    .INIT_41(256'h022bfc22546206b0022bfc0113420798022bfc225463215f022bfc011331d002),
    .INIT_42(256'h022bfc22546206b0022bfc0113620766022bfc22546206b0022bfc0113520766),
    .INIT_43(256'h022bfc22546207ef022bfc01138207c4022bfc2254601101022bfc0113701080),
    .INIT_44(256'h022bfc22546207ac022bfc01141207db022bfc2254601008022bfc0113901100),
    .INIT_45(256'h022bfc22546207ac022bfc011432023b022bfc22546207ac022bfc0114220232),
    .INIT_46(256'h022bfc22546206b0022bfc011452024d022bfc22546207ac022bfc0114420244),
    .INIT_47(256'h022bfc22546206b0022bfc0114720766022bfc22546206b0022bfc0114620766),
    .INIT_48(256'h022bfc2254601018022bfc0114901100022bfc22546207ef022bfc011482026c),
    .INIT_49(256'h022bfc22546207c4022bfc0114b01101022bfc22546010c0022bfc0114a207db),
    .INIT_4A(256'h022bfc2254620256022bfc0114d01100022bfc2254601018022bfc0114c207ac),
    .INIT_4B(256'h022bfc225460b002022bfc0114f207db022bfc2254601018022bfc0114e01100),
    .INIT_4C(256'h022bfc22546206b0022bfc0115120798022bfc225463215f022bfc011501d003),
    .INIT_4D(256'h022bfc22546206b0022bfc0115320766022bfc22546206b0022bfc0115220766),
    .INIT_4E(256'h022bfc2254601101022bfc0115501080022bfc22546206b0022bfc0115420766),
    .INIT_4F(256'h022bfc225460100c022bfc0115701100022bfc22546207ef022bfc01156207c4),
    .INIT_50(256'h022bfc22546207b6022bfc0115920232022bfc22546207b6022bfc01158207db),
    .INIT_51(256'h022bfc2d106207b6022bfc2054d20244022bfc22546207b6022bfc0115a2023b),
    .INIT_52(256'h022bfc36549206b0022bfc0d02020766022bfc0900d206b0022bfc250002024d),
    .INIT_53(256'h022bfc3654d206b0022bfc0d01020766022bfc0900d206b0022bfc2500020766),
    .INIT_54(256'h022bfc250000101c022bfc0306001100022bfc09000207ef022bfc250002026c),
    .INIT_55(256'h022bfc09013207c4022bfc2500001101022bfc0309f010c0022bfc09000207db),
    .INIT_56(256'h022bfc0316020256022bfc0010001100022bfc250000101c022bfc03007207b6),
    .INIT_57(256'h022bfc2051c206bd022bfc2d100207db022bfc041000101c022bfc2055401100),
    .INIT_58(256'h022bfc204cb207a6022bfc20551206bd022bfc204f4207a6022bfc20516206ba),
    .INIT_59(256'h022bfc0319f32173022bfc001001d002022bfc250000b002022bfc204f2206ba),
    .INIT_5A(256'h022bfc20536206ba022bfc2d100207ac022bfc04100206bd022bfc20551207ac),
    .INIT_5B(256'h022bfc1d001207b6022bfc0b03232173022bfc204f41d003022bfc205160b002),
    .INIT_5C(256'h022bfc204f2202a6022bfc204cb206ba022bfc20554207b6022bfc32590206bd),
    .INIT_5D(256'h022bfc204f43217d022bfc205161d002022bfc205360b002022bfc25000202af),
    .INIT_5E(256'h022bfc250003217d022bfc204f21d003022bfc204cb0b002022bfc01002202b8),
    .INIT_5F(256'h022bfc0410001002022bfc205512b02e022bfc0319f2076c022bfc00100202c1),
    .INIT_60(256'h022bfc2057c01002022bfc010002d010022bfc2500001002022bfc2d1002d00f),
    .INIT_61(256'h022bfc205162083d022bfc205362b02e022bfc2d10320839022bfc0b1322d011),
    .INIT_62(256'h022bfc325901d002022bfc1d0010b002022bfc0b0322d00f022bfc204f401002),
    .INIT_63(256'h022bfc250002d010022bfc204f201002022bfc204cb20841022bfc0104032196),
    .INIT_64(256'h022bfc2500020845022bfc204f232196022bfc204cb1d003022bfc010200b002),
    .INIT_65(256'h022bfc2052e2b02e022bfc3259b20839022bfc1d0002d011022bfc2055401002),
    .INIT_66(256'h022bfc205220b002022bfc250002d00f022bfc204f401002022bfc204f82083d),
    .INIT_67(256'h022bfc204f401002022bfc2052c20841022bfc20536321a7022bfc225981d002),
    .INIT_68(256'h022bfc2056b321a7022bfc204f21d003022bfc204cc0b002022bfc00c302d010),
    .INIT_69(256'h022bfc204f420798022bfc205222d011022bfc2053401002022bfc2055f20845),
    .INIT_6A(256'h022bfc250002026c022bfc204f2206b0022bfc204cc20213022bfc0bc3a20209),
    .INIT_6B(256'h022bfc204fe01100022bfc204f420261022bfc2051c01100022bfc2052a01010),
    .INIT_6C(256'h022bfc0bc052026c022bfc204cc207a6022bfc0bc06207db022bfc204fe01010),
    .INIT_6D(256'h022bfc204f201100022bfc204cc20261022bfc0bc0401100022bfc204cc01014),
    .INIT_6E(256'h022bfc204f41d002022bfc205140b002022bfc20538207db022bfc2060201014),
    .INIT_6F(256'h022bfc2061401018022bfc3a5c12026c022bfc0d504207ac022bfc09502321d0),
    .INIT_70(256'h022bfc09e1e01018022bfc09d1d01100022bfc09c1c20261022bfc225d801100),
    .INIT_71(256'h022bfc14b06321d0022bfc14b061d003022bfc0bb130b002022bfc09f1f207db),
    .INIT_72(256'h022bfc13f0001100022bfc13e000101c022bfc13d002026c022bfc10cb0207b6),
    .INIT_73(256'h022bfc2fc34207db022bfc2fd350101c022bfc2fe3601100022bfc2ff3b20261),
    .INIT_74(256'h022bfc204cc0300f022bfc0bc3609001022bfc204cc2b04e022bfc0bc3b20209),
    .INIT_75(256'h022bfc204cc0d002022bfc0bc3409002022bfc204cc321f7022bfc0bc351d001),
    .INIT_76(256'h022bfc204f42b40f022bfc205142b20f022bfc205162076c022bfc204f2321e8),
    .INIT_77(256'h022bfc225f62b10f022bfc206142b08f022bfc3a5e02b04f022bfc0d5042b80f),
    .INIT_78(256'h022bfc0bf3b2d010022bfc0be360101c022bfc0bd352d010022bfc0bc34010e0),
    .INIT_79(256'h022bfc2043f2200a022bfc2048920594022bfc01b0020566022bfc01a0401002),
    .INIT_7A(256'h022bfc2043f1d002022bfc09e070b002022bfc2043f20280022bfc09f0720277),
    .INIT_7B(256'h022bfc204cc1d003022bfc09c070b002022bfc2043f20289022bfc09d07321f2),
    .INIT_7C(256'h022bfc204cc01000022bfc00ce02076c022bfc204cc20292022bfc00cd0321f2),
    .INIT_7D(256'h022bfc205162076c022bfc204f22200a022bfc204cc20594022bfc00cf020566),
    .INIT_7E(256'h022bfc01c002b04f022bfc204fe2b80f022bfc204f42b40f022bfc205282b20f),
    .INIT_7F(256'h022bfc204cc2d010022bfc11c01010e0022bfc14c002b10f022bfc0d5042b08f),
    .INITP_00(256'h727aeadc538f3bd9219076dfc5724df71e09689d20f3cb5a1605a5a1f7b3327c),
    .INITP_01(256'h579602dad50f03576fb4b057f7fdff891ef0813cee40724e4b49afacd515045c),
    .INITP_02(256'h13dd9e48b723834182e182177424dd3d3b9e87241d153afae82e0dd3eca69bd3),
    .INITP_03(256'h0706173a8d2d3180270a21b7966608a3abe704273618522e3804f90682243a29),
    .INITP_04(256'h12de69898ad2d5949d6a582f8ef61cc36c792167104c96ff9fc8a9aea9bea73f),
    .INITP_05(256'h43d965628321b963f0c0ea8fb936d052ee721707aafa6343419c3210e5cd5125),
    .INITP_06(256'h646a71f6715171dabc2a8ba8248e94a5861b988d57a007bb7ec16e6ce80920a1),
    .INITP_07(256'hf3d576d5f14cfe44766b7a4d72c97461c9575ef7faf24e6bc3daf45f5f747478),
    .INITP_08(256'h726e727472fc7762777077ee77647e527acdf7c9725472d5724f714bfac576cf),
    .INITP_09(256'hf8f67a69f7ec727172ec72f672f771f7fa7ef7eff36ef777f16afe78f7727a6e),
    .INITP_0A(256'he1f0dfd9c5f3774ac7f169d677615374ececc074f06dc07df44b7c697c6c7c7d),
    .INITP_0B(256'h52cd44f1785c48624dfc72f5c342d1c1cde1db6d7878dedcceecfc4447dbc667),
    .INITP_0C(256'hcf757aecf0eecf5eedc7ce51e5c65ae6e048d7d0da4b73cf7beee4ddd3e5fae7),
    .INITP_0D(256'h7ccc6dce58f66de4c05fea59f6dafac54143e56774c6d2f3c16fef52de5cd5c0),
    .INITP_0E(256'h4168dfe4d36d67ca52f65f68c26bc8e9e55251edf0d652537ae8c5ccfd784552),
    .INITP_0F(256'hc9c547f964cbd36d67595259564bdd4fc74d56e147e9d2cac1f5de617e51c06b),
