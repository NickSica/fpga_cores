      parameter integer C_PROBE0_WIDTH         = 1,
      parameter integer C_PROBE1_WIDTH         = 1,
      parameter integer C_PROBE2_WIDTH         = 1,
      parameter integer C_PROBE3_WIDTH         = 1,
      parameter integer C_PROBE4_WIDTH         = 1,
      parameter integer C_PROBE5_WIDTH         = 1,
      parameter integer C_PROBE6_WIDTH         = 1,
      parameter integer C_PROBE7_WIDTH         = 1,
      parameter integer C_PROBE8_WIDTH         = 1,
      parameter integer C_PROBE9_WIDTH         = 1,
      parameter integer C_PROBE10_WIDTH        = 1,
      parameter integer C_PROBE11_WIDTH        = 1,
      parameter integer C_PROBE12_WIDTH        = 1,
      parameter integer C_PROBE13_WIDTH        = 1,
      parameter integer C_PROBE14_WIDTH        = 1,
      parameter integer C_PROBE15_WIDTH        = 1,
      parameter integer C_PROBE16_WIDTH        = 1,
      parameter integer C_PROBE17_WIDTH        = 1,
      parameter integer C_PROBE18_WIDTH        = 1,
      parameter integer C_PROBE19_WIDTH        = 1,
      parameter integer C_PROBE20_WIDTH        = 1,
      parameter integer C_PROBE21_WIDTH        = 1,
      parameter integer C_PROBE22_WIDTH        = 1,
      parameter integer C_PROBE23_WIDTH        = 1,
      parameter integer C_PROBE24_WIDTH        = 1,
      parameter integer C_PROBE25_WIDTH        = 1,
      parameter integer C_PROBE26_WIDTH        = 1,
      parameter integer C_PROBE27_WIDTH        = 1,
      parameter integer C_PROBE28_WIDTH        = 1,
      parameter integer C_PROBE29_WIDTH        = 1,
      parameter integer C_PROBE30_WIDTH        = 1,
      parameter integer C_PROBE31_WIDTH        = 1,
      parameter integer C_PROBE32_WIDTH        = 1,
      parameter integer C_PROBE33_WIDTH        = 1,
      parameter integer C_PROBE34_WIDTH        = 1,
      parameter integer C_PROBE35_WIDTH        = 1,
      parameter integer C_PROBE36_WIDTH        = 1,
      parameter integer C_PROBE37_WIDTH        = 1,
      parameter integer C_PROBE38_WIDTH        = 1,
      parameter integer C_PROBE39_WIDTH        = 1,
      parameter integer C_PROBE40_WIDTH        = 1,
      parameter integer C_PROBE41_WIDTH        = 1,
      parameter integer C_PROBE42_WIDTH        = 1,
      parameter integer C_PROBE43_WIDTH        = 1,
      parameter integer C_PROBE44_WIDTH        = 1,
      parameter integer C_PROBE45_WIDTH        = 1,
      parameter integer C_PROBE46_WIDTH        = 1,
      parameter integer C_PROBE47_WIDTH        = 1,
      parameter integer C_PROBE48_WIDTH        = 1,
      parameter integer C_PROBE49_WIDTH        = 1,
      parameter integer C_PROBE50_WIDTH        = 1,
      parameter integer C_PROBE51_WIDTH        = 1,
      parameter integer C_PROBE52_WIDTH        = 1,
      parameter integer C_PROBE53_WIDTH        = 1,
      parameter integer C_PROBE54_WIDTH        = 1,
      parameter integer C_PROBE55_WIDTH        = 1,
      parameter integer C_PROBE56_WIDTH        = 1,
      parameter integer C_PROBE57_WIDTH        = 1,
      parameter integer C_PROBE58_WIDTH        = 1,
      parameter integer C_PROBE59_WIDTH        = 1,
      parameter integer C_PROBE60_WIDTH        = 1,
      parameter integer C_PROBE61_WIDTH        = 1,
      parameter integer C_PROBE62_WIDTH        = 1,
      parameter integer C_PROBE63_WIDTH        = 1,
      parameter integer C_PROBE64_WIDTH        = 1,
      parameter integer C_PROBE65_WIDTH        = 1,
      parameter integer C_PROBE66_WIDTH        = 1,
      parameter integer C_PROBE67_WIDTH        = 1,
      parameter integer C_PROBE68_WIDTH        = 1,
      parameter integer C_PROBE69_WIDTH        = 1,
      parameter integer C_PROBE70_WIDTH        = 1,
      parameter integer C_PROBE71_WIDTH        = 1,
      parameter integer C_PROBE72_WIDTH        = 1,
      parameter integer C_PROBE73_WIDTH        = 1,
      parameter integer C_PROBE74_WIDTH        = 1,
      parameter integer C_PROBE75_WIDTH        = 1,
      parameter integer C_PROBE76_WIDTH        = 1,
      parameter integer C_PROBE77_WIDTH        = 1,
      parameter integer C_PROBE78_WIDTH        = 1,
      parameter integer C_PROBE79_WIDTH        = 1,
      parameter integer C_PROBE80_WIDTH        = 1,
      parameter integer C_PROBE81_WIDTH        = 1,
      parameter integer C_PROBE82_WIDTH        = 1,
      parameter integer C_PROBE83_WIDTH        = 1,
      parameter integer C_PROBE84_WIDTH        = 1,
      parameter integer C_PROBE85_WIDTH        = 1,
      parameter integer C_PROBE86_WIDTH        = 1,
      parameter integer C_PROBE87_WIDTH        = 1,
      parameter integer C_PROBE88_WIDTH        = 1,
      parameter integer C_PROBE89_WIDTH        = 1,
      parameter integer C_PROBE90_WIDTH        = 1,
      parameter integer C_PROBE91_WIDTH        = 1,
      parameter integer C_PROBE92_WIDTH        = 1,
      parameter integer C_PROBE93_WIDTH        = 1,
      parameter integer C_PROBE94_WIDTH        = 1,
      parameter integer C_PROBE95_WIDTH        = 1,
      parameter integer C_PROBE96_WIDTH        = 1,
      parameter integer C_PROBE97_WIDTH        = 1,
      parameter integer C_PROBE98_WIDTH        = 1,
      parameter integer C_PROBE99_WIDTH        = 1,
      parameter integer C_PROBE100_WIDTH       = 1,
      parameter integer C_PROBE101_WIDTH       = 1,
      parameter integer C_PROBE102_WIDTH       = 1,
      parameter integer C_PROBE103_WIDTH       = 1,
      parameter integer C_PROBE104_WIDTH       = 1,
      parameter integer C_PROBE105_WIDTH       = 1,
      parameter integer C_PROBE106_WIDTH       = 1,
      parameter integer C_PROBE107_WIDTH       = 1,
      parameter integer C_PROBE108_WIDTH       = 1,
      parameter integer C_PROBE109_WIDTH       = 1,
      parameter integer C_PROBE110_WIDTH       = 1,
      parameter integer C_PROBE111_WIDTH       = 1,
      parameter integer C_PROBE112_WIDTH       = 1,
      parameter integer C_PROBE113_WIDTH       = 1,
      parameter integer C_PROBE114_WIDTH       = 1,
      parameter integer C_PROBE115_WIDTH       = 1,
      parameter integer C_PROBE116_WIDTH       = 1,
      parameter integer C_PROBE117_WIDTH       = 1,
      parameter integer C_PROBE118_WIDTH       = 1,
      parameter integer C_PROBE119_WIDTH       = 1,
      parameter integer C_PROBE120_WIDTH       = 1,
      parameter integer C_PROBE121_WIDTH       = 1,
      parameter integer C_PROBE122_WIDTH       = 1,
      parameter integer C_PROBE123_WIDTH       = 1,
      parameter integer C_PROBE124_WIDTH       = 1,
      parameter integer C_PROBE125_WIDTH       = 1,
      parameter integer C_PROBE126_WIDTH       = 1,
      parameter integer C_PROBE127_WIDTH       = 1,
      parameter integer C_PROBE128_WIDTH       = 1,
      parameter integer C_PROBE129_WIDTH       = 1,
      parameter integer C_PROBE130_WIDTH       = 1,
      parameter integer C_PROBE131_WIDTH       = 1,
      parameter integer C_PROBE132_WIDTH       = 1,
      parameter integer C_PROBE133_WIDTH       = 1,
      parameter integer C_PROBE134_WIDTH       = 1,
      parameter integer C_PROBE135_WIDTH       = 1,
      parameter integer C_PROBE136_WIDTH       = 1,
      parameter integer C_PROBE137_WIDTH       = 1,
      parameter integer C_PROBE138_WIDTH       = 1,
      parameter integer C_PROBE139_WIDTH       = 1,
      parameter integer C_PROBE140_WIDTH       = 1,
      parameter integer C_PROBE141_WIDTH       = 1,
      parameter integer C_PROBE142_WIDTH       = 1,
      parameter integer C_PROBE143_WIDTH       = 1,
      parameter integer C_PROBE144_WIDTH       = 1,
      parameter integer C_PROBE145_WIDTH       = 1,
      parameter integer C_PROBE146_WIDTH       = 1,
      parameter integer C_PROBE147_WIDTH       = 1,
      parameter integer C_PROBE148_WIDTH       = 1,
      parameter integer C_PROBE149_WIDTH       = 1,
      parameter integer C_PROBE150_WIDTH       = 1,
      parameter integer C_PROBE151_WIDTH       = 1,
      parameter integer C_PROBE152_WIDTH       = 1,
      parameter integer C_PROBE153_WIDTH       = 1,
      parameter integer C_PROBE154_WIDTH       = 1,
      parameter integer C_PROBE155_WIDTH       = 1,
      parameter integer C_PROBE156_WIDTH       = 1,
      parameter integer C_PROBE157_WIDTH       = 1,
      parameter integer C_PROBE158_WIDTH       = 1,
      parameter integer C_PROBE159_WIDTH       = 1,
      parameter integer C_PROBE160_WIDTH       = 1,
      parameter integer C_PROBE161_WIDTH       = 1,
      parameter integer C_PROBE162_WIDTH       = 1,
      parameter integer C_PROBE163_WIDTH       = 1,
      parameter integer C_PROBE164_WIDTH       = 1,
      parameter integer C_PROBE165_WIDTH       = 1,
      parameter integer C_PROBE166_WIDTH       = 1,
      parameter integer C_PROBE167_WIDTH       = 1,
      parameter integer C_PROBE168_WIDTH       = 1,
      parameter integer C_PROBE169_WIDTH       = 1,
      parameter integer C_PROBE170_WIDTH       = 1,
      parameter integer C_PROBE171_WIDTH       = 1,
      parameter integer C_PROBE172_WIDTH       = 1,
      parameter integer C_PROBE173_WIDTH       = 1,
      parameter integer C_PROBE174_WIDTH       = 1,
      parameter integer C_PROBE175_WIDTH       = 1,
      parameter integer C_PROBE176_WIDTH       = 1,
      parameter integer C_PROBE177_WIDTH       = 1,
      parameter integer C_PROBE178_WIDTH       = 1,
      parameter integer C_PROBE179_WIDTH       = 1,
      parameter integer C_PROBE180_WIDTH       = 1,
      parameter integer C_PROBE181_WIDTH       = 1,
      parameter integer C_PROBE182_WIDTH       = 1,
      parameter integer C_PROBE183_WIDTH       = 1,
      parameter integer C_PROBE184_WIDTH       = 1,
      parameter integer C_PROBE185_WIDTH       = 1,
      parameter integer C_PROBE186_WIDTH       = 1,
      parameter integer C_PROBE187_WIDTH       = 1,
      parameter integer C_PROBE188_WIDTH       = 1,
      parameter integer C_PROBE189_WIDTH       = 1,
      parameter integer C_PROBE190_WIDTH       = 1,
      parameter integer C_PROBE191_WIDTH       = 1,
      parameter integer C_PROBE192_WIDTH       = 1,
      parameter integer C_PROBE193_WIDTH       = 1,
      parameter integer C_PROBE194_WIDTH       = 1,
      parameter integer C_PROBE195_WIDTH       = 1,
      parameter integer C_PROBE196_WIDTH       = 1,
      parameter integer C_PROBE197_WIDTH       = 1,
      parameter integer C_PROBE198_WIDTH       = 1,
      parameter integer C_PROBE199_WIDTH       = 1,
      parameter integer C_PROBE200_WIDTH       = 1,
      parameter integer C_PROBE201_WIDTH       = 1,
      parameter integer C_PROBE202_WIDTH       = 1,
      parameter integer C_PROBE203_WIDTH       = 1,
      parameter integer C_PROBE204_WIDTH       = 1,
      parameter integer C_PROBE205_WIDTH       = 1,
      parameter integer C_PROBE206_WIDTH       = 1,
      parameter integer C_PROBE207_WIDTH       = 1,
      parameter integer C_PROBE208_WIDTH       = 1,
      parameter integer C_PROBE209_WIDTH       = 1,
      parameter integer C_PROBE210_WIDTH       = 1,
      parameter integer C_PROBE211_WIDTH       = 1,
      parameter integer C_PROBE212_WIDTH       = 1,
      parameter integer C_PROBE213_WIDTH       = 1,
      parameter integer C_PROBE214_WIDTH       = 1,
      parameter integer C_PROBE215_WIDTH       = 1,
      parameter integer C_PROBE216_WIDTH       = 1,
      parameter integer C_PROBE217_WIDTH       = 1,
      parameter integer C_PROBE218_WIDTH       = 1,
      parameter integer C_PROBE219_WIDTH       = 1,
      parameter integer C_PROBE220_WIDTH       = 1,
      parameter integer C_PROBE221_WIDTH       = 1,
      parameter integer C_PROBE222_WIDTH       = 1,
      parameter integer C_PROBE223_WIDTH       = 1,
      parameter integer C_PROBE224_WIDTH       = 1,
      parameter integer C_PROBE225_WIDTH       = 1,
      parameter integer C_PROBE226_WIDTH       = 1,
      parameter integer C_PROBE227_WIDTH       = 1,
      parameter integer C_PROBE228_WIDTH       = 1,
      parameter integer C_PROBE229_WIDTH       = 1,
      parameter integer C_PROBE230_WIDTH       = 1,
      parameter integer C_PROBE231_WIDTH       = 1,
      parameter integer C_PROBE232_WIDTH       = 1,
      parameter integer C_PROBE233_WIDTH       = 1,
      parameter integer C_PROBE234_WIDTH       = 1,
      parameter integer C_PROBE235_WIDTH       = 1,
      parameter integer C_PROBE236_WIDTH       = 1,
      parameter integer C_PROBE237_WIDTH       = 1,
      parameter integer C_PROBE238_WIDTH       = 1,
      parameter integer C_PROBE239_WIDTH       = 1,
      parameter integer C_PROBE240_WIDTH       = 1,
      parameter integer C_PROBE241_WIDTH       = 1,
      parameter integer C_PROBE242_WIDTH       = 1,
      parameter integer C_PROBE243_WIDTH       = 1,
      parameter integer C_PROBE244_WIDTH       = 1,
      parameter integer C_PROBE245_WIDTH       = 1,
      parameter integer C_PROBE246_WIDTH       = 1,
      parameter integer C_PROBE247_WIDTH       = 1,
      parameter integer C_PROBE248_WIDTH       = 1,
      parameter integer C_PROBE249_WIDTH       = 1,
      parameter integer C_PROBE250_WIDTH       = 1,
      parameter integer C_PROBE251_WIDTH       = 1,
      parameter integer C_PROBE252_WIDTH       = 1,
      parameter integer C_PROBE253_WIDTH       = 1,
      parameter integer C_PROBE254_WIDTH       = 1,
      parameter integer C_PROBE255_WIDTH       = 1,
      parameter integer C_PROBE256_WIDTH        = 1,
      parameter integer C_PROBE257_WIDTH        = 1,
      parameter integer C_PROBE258_WIDTH        = 1,
      parameter integer C_PROBE259_WIDTH        = 1,
      parameter integer C_PROBE260_WIDTH        = 1,
      parameter integer C_PROBE261_WIDTH        = 1,
      parameter integer C_PROBE262_WIDTH        = 1,
      parameter integer C_PROBE263_WIDTH        = 1,
      parameter integer C_PROBE264_WIDTH        = 1,
      parameter integer C_PROBE265_WIDTH        = 1,
      parameter integer C_PROBE266_WIDTH        = 1,
      parameter integer C_PROBE267_WIDTH        = 1,
      parameter integer C_PROBE268_WIDTH        = 1,
      parameter integer C_PROBE269_WIDTH        = 1,
      parameter integer C_PROBE270_WIDTH        = 1,
      parameter integer C_PROBE271_WIDTH        = 1,
      parameter integer C_PROBE272_WIDTH        = 1,
      parameter integer C_PROBE273_WIDTH        = 1,
      parameter integer C_PROBE274_WIDTH        = 1,
      parameter integer C_PROBE275_WIDTH        = 1,
      parameter integer C_PROBE276_WIDTH        = 1,
      parameter integer C_PROBE277_WIDTH        = 1,
      parameter integer C_PROBE278_WIDTH        = 1,
      parameter integer C_PROBE279_WIDTH        = 1,
      parameter integer C_PROBE280_WIDTH        = 1,
      parameter integer C_PROBE281_WIDTH        = 1,
      parameter integer C_PROBE282_WIDTH        = 1,
      parameter integer C_PROBE283_WIDTH        = 1,
      parameter integer C_PROBE284_WIDTH        = 1,
      parameter integer C_PROBE285_WIDTH        = 1,
      parameter integer C_PROBE286_WIDTH        = 1,
      parameter integer C_PROBE287_WIDTH        = 1,
      parameter integer C_PROBE288_WIDTH        = 1,
      parameter integer C_PROBE289_WIDTH        = 1,
      parameter integer C_PROBE290_WIDTH        = 1,
      parameter integer C_PROBE291_WIDTH        = 1,
      parameter integer C_PROBE292_WIDTH        = 1,
      parameter integer C_PROBE293_WIDTH        = 1,
      parameter integer C_PROBE294_WIDTH        = 1,
      parameter integer C_PROBE295_WIDTH        = 1,
      parameter integer C_PROBE296_WIDTH        = 1,
      parameter integer C_PROBE297_WIDTH        = 1,
      parameter integer C_PROBE298_WIDTH        = 1,
      parameter integer C_PROBE299_WIDTH        = 1,
      parameter integer C_PROBE300_WIDTH        = 1,
      parameter integer C_PROBE301_WIDTH        = 1,
      parameter integer C_PROBE302_WIDTH        = 1,
      parameter integer C_PROBE303_WIDTH        = 1,
      parameter integer C_PROBE304_WIDTH        = 1,
      parameter integer C_PROBE305_WIDTH        = 1,
      parameter integer C_PROBE306_WIDTH        = 1,
      parameter integer C_PROBE307_WIDTH        = 1,
      parameter integer C_PROBE308_WIDTH        = 1,
      parameter integer C_PROBE309_WIDTH        = 1,
      parameter integer C_PROBE310_WIDTH        = 1,
      parameter integer C_PROBE311_WIDTH        = 1,
      parameter integer C_PROBE312_WIDTH        = 1,
      parameter integer C_PROBE313_WIDTH        = 1,
      parameter integer C_PROBE314_WIDTH        = 1,
      parameter integer C_PROBE315_WIDTH        = 1,
      parameter integer C_PROBE316_WIDTH        = 1,
      parameter integer C_PROBE317_WIDTH        = 1,
      parameter integer C_PROBE318_WIDTH        = 1,
      parameter integer C_PROBE319_WIDTH        = 1,
      parameter integer C_PROBE320_WIDTH        = 1,
      parameter integer C_PROBE321_WIDTH        = 1,
      parameter integer C_PROBE322_WIDTH        = 1,
      parameter integer C_PROBE323_WIDTH        = 1,
      parameter integer C_PROBE324_WIDTH        = 1,
      parameter integer C_PROBE325_WIDTH        = 1,
      parameter integer C_PROBE326_WIDTH        = 1,
      parameter integer C_PROBE327_WIDTH        = 1,
      parameter integer C_PROBE328_WIDTH        = 1,
      parameter integer C_PROBE329_WIDTH        = 1,
      parameter integer C_PROBE330_WIDTH        = 1,
      parameter integer C_PROBE331_WIDTH        = 1,
      parameter integer C_PROBE332_WIDTH        = 1,
      parameter integer C_PROBE333_WIDTH        = 1,
      parameter integer C_PROBE334_WIDTH        = 1,
      parameter integer C_PROBE335_WIDTH        = 1,
      parameter integer C_PROBE336_WIDTH        = 1,
      parameter integer C_PROBE337_WIDTH        = 1,
      parameter integer C_PROBE338_WIDTH        = 1,
      parameter integer C_PROBE339_WIDTH        = 1,
      parameter integer C_PROBE340_WIDTH        = 1,
      parameter integer C_PROBE341_WIDTH        = 1,
      parameter integer C_PROBE342_WIDTH        = 1,
      parameter integer C_PROBE343_WIDTH        = 1,
      parameter integer C_PROBE344_WIDTH        = 1,
      parameter integer C_PROBE345_WIDTH        = 1,
      parameter integer C_PROBE346_WIDTH        = 1,
      parameter integer C_PROBE347_WIDTH        = 1,
      parameter integer C_PROBE348_WIDTH        = 1,
      parameter integer C_PROBE349_WIDTH        = 1,
      parameter integer C_PROBE350_WIDTH        = 1,
      parameter integer C_PROBE351_WIDTH        = 1,
      parameter integer C_PROBE352_WIDTH        = 1,
      parameter integer C_PROBE353_WIDTH        = 1,
      parameter integer C_PROBE354_WIDTH        = 1,
      parameter integer C_PROBE355_WIDTH        = 1,
      parameter integer C_PROBE356_WIDTH        = 1,
      parameter integer C_PROBE357_WIDTH        = 1,
      parameter integer C_PROBE358_WIDTH        = 1,
      parameter integer C_PROBE359_WIDTH        = 1,
      parameter integer C_PROBE360_WIDTH        = 1,
      parameter integer C_PROBE361_WIDTH        = 1,
      parameter integer C_PROBE362_WIDTH        = 1,
      parameter integer C_PROBE363_WIDTH        = 1,
      parameter integer C_PROBE364_WIDTH        = 1,
      parameter integer C_PROBE365_WIDTH        = 1,
      parameter integer C_PROBE366_WIDTH        = 1,
      parameter integer C_PROBE367_WIDTH        = 1,
      parameter integer C_PROBE368_WIDTH        = 1,
      parameter integer C_PROBE369_WIDTH        = 1,
      parameter integer C_PROBE370_WIDTH        = 1,
      parameter integer C_PROBE371_WIDTH        = 1,
      parameter integer C_PROBE372_WIDTH        = 1,
      parameter integer C_PROBE373_WIDTH        = 1,
      parameter integer C_PROBE374_WIDTH        = 1,
      parameter integer C_PROBE375_WIDTH        = 1,
      parameter integer C_PROBE376_WIDTH        = 1,
      parameter integer C_PROBE377_WIDTH        = 1,
      parameter integer C_PROBE378_WIDTH        = 1,
      parameter integer C_PROBE379_WIDTH        = 1,
      parameter integer C_PROBE380_WIDTH        = 1,
      parameter integer C_PROBE381_WIDTH        = 1,
      parameter integer C_PROBE382_WIDTH        = 1,
      parameter integer C_PROBE383_WIDTH        = 1,
      parameter integer C_PROBE384_WIDTH        = 1,
      parameter integer C_PROBE385_WIDTH        = 1,
      parameter integer C_PROBE386_WIDTH        = 1,
      parameter integer C_PROBE387_WIDTH        = 1,
      parameter integer C_PROBE388_WIDTH        = 1,
      parameter integer C_PROBE389_WIDTH        = 1,
      parameter integer C_PROBE390_WIDTH        = 1,
      parameter integer C_PROBE391_WIDTH        = 1,
      parameter integer C_PROBE392_WIDTH        = 1,
      parameter integer C_PROBE393_WIDTH        = 1,
      parameter integer C_PROBE394_WIDTH        = 1,
      parameter integer C_PROBE395_WIDTH        = 1,
      parameter integer C_PROBE396_WIDTH        = 1,
      parameter integer C_PROBE397_WIDTH        = 1,
      parameter integer C_PROBE398_WIDTH        = 1,
      parameter integer C_PROBE399_WIDTH        = 1,
      parameter integer C_PROBE400_WIDTH        = 1,
      parameter integer C_PROBE401_WIDTH        = 1,
      parameter integer C_PROBE402_WIDTH        = 1,
      parameter integer C_PROBE403_WIDTH        = 1,
      parameter integer C_PROBE404_WIDTH        = 1,
      parameter integer C_PROBE405_WIDTH        = 1,
      parameter integer C_PROBE406_WIDTH        = 1,
      parameter integer C_PROBE407_WIDTH        = 1,
      parameter integer C_PROBE408_WIDTH        = 1,
      parameter integer C_PROBE409_WIDTH        = 1,
      parameter integer C_PROBE410_WIDTH        = 1,
      parameter integer C_PROBE411_WIDTH        = 1,
      parameter integer C_PROBE412_WIDTH        = 1,
      parameter integer C_PROBE413_WIDTH        = 1,
      parameter integer C_PROBE414_WIDTH        = 1,
      parameter integer C_PROBE415_WIDTH        = 1,
      parameter integer C_PROBE416_WIDTH        = 1,
      parameter integer C_PROBE417_WIDTH        = 1,
      parameter integer C_PROBE418_WIDTH        = 1,
      parameter integer C_PROBE419_WIDTH        = 1,
      parameter integer C_PROBE420_WIDTH        = 1,
      parameter integer C_PROBE421_WIDTH        = 1,
      parameter integer C_PROBE422_WIDTH        = 1,
      parameter integer C_PROBE423_WIDTH        = 1,
      parameter integer C_PROBE424_WIDTH        = 1,
      parameter integer C_PROBE425_WIDTH        = 1,
      parameter integer C_PROBE426_WIDTH        = 1,
      parameter integer C_PROBE427_WIDTH        = 1,
      parameter integer C_PROBE428_WIDTH        = 1,
      parameter integer C_PROBE429_WIDTH        = 1,
      parameter integer C_PROBE430_WIDTH        = 1,
      parameter integer C_PROBE431_WIDTH        = 1,
      parameter integer C_PROBE432_WIDTH        = 1,
      parameter integer C_PROBE433_WIDTH        = 1,
      parameter integer C_PROBE434_WIDTH        = 1,
      parameter integer C_PROBE435_WIDTH        = 1,
      parameter integer C_PROBE436_WIDTH        = 1,
      parameter integer C_PROBE437_WIDTH        = 1,
      parameter integer C_PROBE438_WIDTH        = 1,
      parameter integer C_PROBE439_WIDTH        = 1,
      parameter integer C_PROBE440_WIDTH        = 1,
      parameter integer C_PROBE441_WIDTH        = 1,
      parameter integer C_PROBE442_WIDTH        = 1,
      parameter integer C_PROBE443_WIDTH        = 1,
      parameter integer C_PROBE444_WIDTH        = 1,
      parameter integer C_PROBE445_WIDTH        = 1,
      parameter integer C_PROBE446_WIDTH        = 1,
      parameter integer C_PROBE447_WIDTH        = 1,
      parameter integer C_PROBE448_WIDTH        = 1,
      parameter integer C_PROBE449_WIDTH        = 1,
      parameter integer C_PROBE450_WIDTH        = 1,
      parameter integer C_PROBE451_WIDTH        = 1,
      parameter integer C_PROBE452_WIDTH        = 1,
      parameter integer C_PROBE453_WIDTH        = 1,
      parameter integer C_PROBE454_WIDTH        = 1,
      parameter integer C_PROBE455_WIDTH        = 1,
      parameter integer C_PROBE456_WIDTH        = 1,
      parameter integer C_PROBE457_WIDTH        = 1,
      parameter integer C_PROBE458_WIDTH        = 1,
      parameter integer C_PROBE459_WIDTH        = 1,
      parameter integer C_PROBE460_WIDTH        = 1,
      parameter integer C_PROBE461_WIDTH        = 1,
      parameter integer C_PROBE462_WIDTH        = 1,
      parameter integer C_PROBE463_WIDTH        = 1,
      parameter integer C_PROBE464_WIDTH        = 1,
      parameter integer C_PROBE465_WIDTH        = 1,
      parameter integer C_PROBE466_WIDTH        = 1,
      parameter integer C_PROBE467_WIDTH        = 1,
      parameter integer C_PROBE468_WIDTH        = 1,
      parameter integer C_PROBE469_WIDTH        = 1,
      parameter integer C_PROBE470_WIDTH        = 1,
      parameter integer C_PROBE471_WIDTH        = 1,
      parameter integer C_PROBE472_WIDTH        = 1,
      parameter integer C_PROBE473_WIDTH        = 1,
      parameter integer C_PROBE474_WIDTH        = 1,
      parameter integer C_PROBE475_WIDTH        = 1,
      parameter integer C_PROBE476_WIDTH        = 1,
      parameter integer C_PROBE477_WIDTH        = 1,
      parameter integer C_PROBE478_WIDTH        = 1,
      parameter integer C_PROBE479_WIDTH        = 1,
      parameter integer C_PROBE480_WIDTH        = 1,
      parameter integer C_PROBE481_WIDTH        = 1,
      parameter integer C_PROBE482_WIDTH        = 1,
      parameter integer C_PROBE483_WIDTH        = 1,
      parameter integer C_PROBE484_WIDTH        = 1,
      parameter integer C_PROBE485_WIDTH        = 1,
      parameter integer C_PROBE486_WIDTH        = 1,
      parameter integer C_PROBE487_WIDTH        = 1,
      parameter integer C_PROBE488_WIDTH        = 1,
      parameter integer C_PROBE489_WIDTH        = 1,
      parameter integer C_PROBE490_WIDTH        = 1,
      parameter integer C_PROBE491_WIDTH        = 1,
      parameter integer C_PROBE492_WIDTH        = 1,
      parameter integer C_PROBE493_WIDTH        = 1,
      parameter integer C_PROBE494_WIDTH        = 1,
      parameter integer C_PROBE495_WIDTH        = 1,
      parameter integer C_PROBE496_WIDTH        = 1,
      parameter integer C_PROBE497_WIDTH        = 1,
      parameter integer C_PROBE498_WIDTH        = 1,
      parameter integer C_PROBE499_WIDTH        = 1,
      parameter integer C_PROBE500_WIDTH        = 1,
      parameter integer C_PROBE501_WIDTH        = 1,
      parameter integer C_PROBE502_WIDTH        = 1,
      parameter integer C_PROBE503_WIDTH        = 1,
      parameter integer C_PROBE504_WIDTH        = 1,
      parameter integer C_PROBE505_WIDTH        = 1,
      parameter integer C_PROBE506_WIDTH        = 1,
      parameter integer C_PROBE507_WIDTH        = 1,
      parameter integer C_PROBE508_WIDTH        = 1,
      parameter integer C_PROBE509_WIDTH        = 1,
      parameter integer C_PROBE510_WIDTH        = 1,
      parameter integer C_PROBE511_WIDTH        = 1,
