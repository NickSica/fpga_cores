
    axis_itct_v1_0_0_mu_itct
    #(
      .C_NUM_PROBES           (C_NUM_PROBES              )
     ) u_mu_itct
     (
      .cfg_clk                (cfg_clk                   ),
      .cfg_in                 (cfg_data_i                ),
      .cfg_en                 (cfg_en_i                  ),
      .aresetn                (resetn                    ),
      .curr_mu                (app_spec_i                ),
      .mu_sel                 (wr_mu_config_i            ),
      .tc_sel                 (wr_tc_config_i            ),
      .cc_sel                 (wr_cc_config_i            ),
      .cfg_out                (cfg_out_o                 ),
      .tc_cfg_out             (tc_cfg_dout               ),
      .cc_cfg_out0            (cc_cfg_dout0              ),
      .cc_cfg_out1            (cc_cfg_dout1              ),
      .cc_cfg_out2            (cc_cfg_dout2              ),
      .cc_cfg_out3            (cc_cfg_dout3              ),
      .tc_cfg_in              (tc_cfg_din                ),
      .cc_cfg_in0             (cc_cfg_din0               ),
      .cc_cfg_in1             (cc_cfg_din1               ),
      .cc_cfg_in2             (cc_cfg_din2               ),
      .cc_cfg_in3             (cc_cfg_din3               ),
      .tc_cfg_en              (tc_cfg_en                 ),
      .cc_cfg_en0             (cc_cfg_en0                ),
      .cc_cfg_en1             (cc_cfg_en1                ),
      .cc_cfg_en2             (cc_cfg_en2                ),
      .cc_cfg_en3             (cc_cfg_en3                ),
      .cfg_out0          (cfg_dout0            ),
      .cfg_out1          (cfg_dout1            ),
      .cfg_out2          (cfg_dout2            ),
      .cfg_out3          (cfg_dout3            ),
      .cfg_out4          (cfg_dout4            ),
      .cfg_out5          (cfg_dout5            ),
      .cfg_out6          (cfg_dout6            ),
      .cfg_out7          (cfg_dout7            ),
      .cfg_out8          (cfg_dout8            ),
      .cfg_out9          (cfg_dout9            ),
      .cfg_out10          (cfg_dout10            ),
      .cfg_out11          (cfg_dout11            ),
      .cfg_out12          (cfg_dout12            ),
      .cfg_out13          (cfg_dout13            ),
      .cfg_out14          (cfg_dout14            ),
      .cfg_out15          (cfg_dout15            ),
      .cfg_out16          (cfg_dout16            ),
      .cfg_out17          (cfg_dout17            ),
      .cfg_out18          (cfg_dout18            ),
      .cfg_out19          (cfg_dout19            ),
      .cfg_out20          (cfg_dout20            ),
      .cfg_out21          (cfg_dout21            ),
      .cfg_out22          (cfg_dout22            ),
      .cfg_out23          (cfg_dout23            ),
      .cfg_out24          (cfg_dout24            ),
      .cfg_out25          (cfg_dout25            ),
      .cfg_out26          (cfg_dout26            ),
      .cfg_out27          (cfg_dout27            ),
      .cfg_out28          (cfg_dout28            ),
      .cfg_out29          (cfg_dout29            ),
      .cfg_out30          (cfg_dout30            ),
      .cfg_out31          (cfg_dout31            ),
      .cfg_out32          (cfg_dout32            ),
      .cfg_out33          (cfg_dout33            ),
      .cfg_out34          (cfg_dout34            ),
      .cfg_out35          (cfg_dout35            ),
      .cfg_out36          (cfg_dout36            ),
      .cfg_out37          (cfg_dout37            ),
      .cfg_out38          (cfg_dout38            ),
      .cfg_out39          (cfg_dout39            ),
      .cfg_out40          (cfg_dout40            ),
      .cfg_out41          (cfg_dout41            ),
      .cfg_out42          (cfg_dout42            ),
      .cfg_out43          (cfg_dout43            ),
      .cfg_out44          (cfg_dout44            ),
      .cfg_out45          (cfg_dout45            ),
      .cfg_out46          (cfg_dout46            ),
      .cfg_out47          (cfg_dout47            ),
      .cfg_out48          (cfg_dout48            ),
      .cfg_out49          (cfg_dout49            ),
      .cfg_out50          (cfg_dout50            ),
      .cfg_out51          (cfg_dout51            ),
      .cfg_out52          (cfg_dout52            ),
      .cfg_out53          (cfg_dout53            ),
      .cfg_out54          (cfg_dout54            ),
      .cfg_out55          (cfg_dout55            ),
      .cfg_out56          (cfg_dout56            ),
      .cfg_out57          (cfg_dout57            ),
      .cfg_out58          (cfg_dout58            ),
      .cfg_out59          (cfg_dout59            ),
      .cfg_out60          (cfg_dout60            ),
      .cfg_out61          (cfg_dout61            ),
      .cfg_out62          (cfg_dout62            ),
      .cfg_out63          (cfg_dout63            ),
      .cfg_out64          (cfg_dout64            ),
      .cfg_out65          (cfg_dout65            ),
      .cfg_out66          (cfg_dout66            ),
      .cfg_out67          (cfg_dout67            ),
      .cfg_out68          (cfg_dout68            ),
      .cfg_out69          (cfg_dout69            ),
      .cfg_out70          (cfg_dout70            ),
      .cfg_out71          (cfg_dout71            ),
      .cfg_out72          (cfg_dout72            ),
      .cfg_out73          (cfg_dout73            ),
      .cfg_out74          (cfg_dout74            ),
      .cfg_out75          (cfg_dout75            ),
      .cfg_out76          (cfg_dout76            ),
      .cfg_out77          (cfg_dout77            ),
      .cfg_out78          (cfg_dout78            ),
      .cfg_out79          (cfg_dout79            ),
      .cfg_out80          (cfg_dout80            ),
      .cfg_out81          (cfg_dout81            ),
      .cfg_out82          (cfg_dout82            ),
      .cfg_out83          (cfg_dout83            ),
      .cfg_out84          (cfg_dout84            ),
      .cfg_out85          (cfg_dout85            ),
      .cfg_out86          (cfg_dout86            ),
      .cfg_out87          (cfg_dout87            ),
      .cfg_out88          (cfg_dout88            ),
      .cfg_out89          (cfg_dout89            ),
      .cfg_out90          (cfg_dout90            ),
      .cfg_out91          (cfg_dout91            ),
      .cfg_out92          (cfg_dout92            ),
      .cfg_out93          (cfg_dout93            ),
      .cfg_out94          (cfg_dout94            ),
      .cfg_out95          (cfg_dout95            ),
      .cfg_out96          (cfg_dout96            ),
      .cfg_out97          (cfg_dout97            ),
      .cfg_out98          (cfg_dout98            ),
      .cfg_out99          (cfg_dout99            ),
      .cfg_out100          (cfg_dout100            ),
      .cfg_out101          (cfg_dout101            ),
      .cfg_out102          (cfg_dout102            ),
      .cfg_out103          (cfg_dout103            ),
      .cfg_out104          (cfg_dout104            ),
      .cfg_out105          (cfg_dout105            ),
      .cfg_out106          (cfg_dout106            ),
      .cfg_out107          (cfg_dout107            ),
      .cfg_out108          (cfg_dout108            ),
      .cfg_out109          (cfg_dout109            ),
      .cfg_out110          (cfg_dout110            ),
      .cfg_out111          (cfg_dout111            ),
      .cfg_out112          (cfg_dout112            ),
      .cfg_out113          (cfg_dout113            ),
      .cfg_out114          (cfg_dout114            ),
      .cfg_out115          (cfg_dout115            ),
      .cfg_out116          (cfg_dout116            ),
      .cfg_out117          (cfg_dout117            ),
      .cfg_out118          (cfg_dout118            ),
      .cfg_out119          (cfg_dout119            ),
      .cfg_out120          (cfg_dout120            ),
      .cfg_out121          (cfg_dout121            ),
      .cfg_out122          (cfg_dout122            ),
      .cfg_out123          (cfg_dout123            ),
      .cfg_out124          (cfg_dout124            ),
      .cfg_out125          (cfg_dout125            ),
      .cfg_out126          (cfg_dout126            ),
      .cfg_out127          (cfg_dout127            ),
      .cfg_out128          (cfg_dout128            ),
      .cfg_out129          (cfg_dout129            ),
      .cfg_out130          (cfg_dout130            ),
      .cfg_out131          (cfg_dout131            ),
      .cfg_out132          (cfg_dout132            ),
      .cfg_out133          (cfg_dout133            ),
      .cfg_out134          (cfg_dout134            ),
      .cfg_out135          (cfg_dout135            ),
      .cfg_out136          (cfg_dout136            ),
      .cfg_out137          (cfg_dout137            ),
      .cfg_out138          (cfg_dout138            ),
      .cfg_out139          (cfg_dout139            ),
      .cfg_out140          (cfg_dout140            ),
      .cfg_out141          (cfg_dout141            ),
      .cfg_out142          (cfg_dout142            ),
      .cfg_out143          (cfg_dout143            ),
      .cfg_out144          (cfg_dout144            ),
      .cfg_out145          (cfg_dout145            ),
      .cfg_out146          (cfg_dout146            ),
      .cfg_out147          (cfg_dout147            ),
      .cfg_out148          (cfg_dout148            ),
      .cfg_out149          (cfg_dout149            ),
      .cfg_out150          (cfg_dout150            ),
      .cfg_out151          (cfg_dout151            ),
      .cfg_out152          (cfg_dout152            ),
      .cfg_out153          (cfg_dout153            ),
      .cfg_out154          (cfg_dout154            ),
      .cfg_out155          (cfg_dout155            ),
      .cfg_out156          (cfg_dout156            ),
      .cfg_out157          (cfg_dout157            ),
      .cfg_out158          (cfg_dout158            ),
      .cfg_out159          (cfg_dout159            ),
      .cfg_out160          (cfg_dout160            ),
      .cfg_out161          (cfg_dout161            ),
      .cfg_out162          (cfg_dout162            ),
      .cfg_out163          (cfg_dout163            ),
      .cfg_out164          (cfg_dout164            ),
      .cfg_out165          (cfg_dout165            ),
      .cfg_out166          (cfg_dout166            ),
      .cfg_out167          (cfg_dout167            ),
      .cfg_out168          (cfg_dout168            ),
      .cfg_out169          (cfg_dout169            ),
      .cfg_out170          (cfg_dout170            ),
      .cfg_out171          (cfg_dout171            ),
      .cfg_out172          (cfg_dout172            ),
      .cfg_out173          (cfg_dout173            ),
      .cfg_out174          (cfg_dout174            ),
      .cfg_out175          (cfg_dout175            ),
      .cfg_out176          (cfg_dout176            ),
      .cfg_out177          (cfg_dout177            ),
      .cfg_out178          (cfg_dout178            ),
      .cfg_out179          (cfg_dout179            ),
      .cfg_out180          (cfg_dout180            ),
      .cfg_out181          (cfg_dout181            ),
      .cfg_out182          (cfg_dout182            ),
      .cfg_out183          (cfg_dout183            ),
      .cfg_out184          (cfg_dout184            ),
      .cfg_out185          (cfg_dout185            ),
      .cfg_out186          (cfg_dout186            ),
      .cfg_out187          (cfg_dout187            ),
      .cfg_out188          (cfg_dout188            ),
      .cfg_out189          (cfg_dout189            ),
      .cfg_out190          (cfg_dout190            ),
      .cfg_out191          (cfg_dout191            ),
      .cfg_out192          (cfg_dout192            ),
      .cfg_out193          (cfg_dout193            ),
      .cfg_out194          (cfg_dout194            ),
      .cfg_out195          (cfg_dout195            ),
      .cfg_out196          (cfg_dout196            ),
      .cfg_out197          (cfg_dout197            ),
      .cfg_out198          (cfg_dout198            ),
      .cfg_out199          (cfg_dout199            ),
      .cfg_out200          (cfg_dout200            ),
      .cfg_out201          (cfg_dout201            ),
      .cfg_out202          (cfg_dout202            ),
      .cfg_out203          (cfg_dout203            ),
      .cfg_out204          (cfg_dout204            ),
      .cfg_out205          (cfg_dout205            ),
      .cfg_out206          (cfg_dout206            ),
      .cfg_out207          (cfg_dout207            ),
      .cfg_out208          (cfg_dout208            ),
      .cfg_out209          (cfg_dout209            ),
      .cfg_out210          (cfg_dout210            ),
      .cfg_out211          (cfg_dout211            ),
      .cfg_out212          (cfg_dout212            ),
      .cfg_out213          (cfg_dout213            ),
      .cfg_out214          (cfg_dout214            ),
      .cfg_out215          (cfg_dout215            ),
      .cfg_out216          (cfg_dout216            ),
      .cfg_out217          (cfg_dout217            ),
      .cfg_out218          (cfg_dout218            ),
      .cfg_out219          (cfg_dout219            ),
      .cfg_out220          (cfg_dout220            ),
      .cfg_out221          (cfg_dout221            ),
      .cfg_out222          (cfg_dout222            ),
      .cfg_out223          (cfg_dout223            ),
      .cfg_out224          (cfg_dout224            ),
      .cfg_out225          (cfg_dout225            ),
      .cfg_out226          (cfg_dout226            ),
      .cfg_out227          (cfg_dout227            ),
      .cfg_out228          (cfg_dout228            ),
      .cfg_out229          (cfg_dout229            ),
      .cfg_out230          (cfg_dout230            ),
      .cfg_out231          (cfg_dout231            ),
      .cfg_out232          (cfg_dout232            ),
      .cfg_out233          (cfg_dout233            ),
      .cfg_out234          (cfg_dout234            ),
      .cfg_out235          (cfg_dout235            ),
      .cfg_out236          (cfg_dout236            ),
      .cfg_out237          (cfg_dout237            ),
      .cfg_out238          (cfg_dout238            ),
      .cfg_out239          (cfg_dout239            ),
      .cfg_out240          (cfg_dout240            ),
      .cfg_out241          (cfg_dout241            ),
      .cfg_out242          (cfg_dout242            ),
      .cfg_out243          (cfg_dout243            ),
      .cfg_out244          (cfg_dout244            ),
      .cfg_out245          (cfg_dout245            ),
      .cfg_out246          (cfg_dout246            ),
      .cfg_out247          (cfg_dout247            ),
      .cfg_out248          (cfg_dout248            ),
      .cfg_out249          (cfg_dout249            ),
      .cfg_out250          (cfg_dout250            ),
      .cfg_out251          (cfg_dout251            ),
      .cfg_out252          (cfg_dout252            ),
      .cfg_out253          (cfg_dout253            ),
      .cfg_out254          (cfg_dout254            ),
      .cfg_out255          (cfg_dout255            ),
      .cfg_out256          (cfg_dout256            ),
      .cfg_out257          (cfg_dout257            ),
      .cfg_out258          (cfg_dout258            ),
      .cfg_out259          (cfg_dout259            ),
      .cfg_out260          (cfg_dout260            ),
      .cfg_out261          (cfg_dout261            ),
      .cfg_out262          (cfg_dout262            ),
      .cfg_out263          (cfg_dout263            ),
      .cfg_out264          (cfg_dout264            ),
      .cfg_out265          (cfg_dout265            ),
      .cfg_out266          (cfg_dout266            ),
      .cfg_out267          (cfg_dout267            ),
      .cfg_out268          (cfg_dout268            ),
      .cfg_out269          (cfg_dout269            ),
      .cfg_out270          (cfg_dout270            ),
      .cfg_out271          (cfg_dout271            ),
      .cfg_out272          (cfg_dout272            ),
      .cfg_out273          (cfg_dout273            ),
      .cfg_out274          (cfg_dout274            ),
      .cfg_out275          (cfg_dout275            ),
      .cfg_out276          (cfg_dout276            ),
      .cfg_out277          (cfg_dout277            ),
      .cfg_out278          (cfg_dout278            ),
      .cfg_out279          (cfg_dout279            ),
      .cfg_out280          (cfg_dout280            ),
      .cfg_out281          (cfg_dout281            ),
      .cfg_out282          (cfg_dout282            ),
      .cfg_out283          (cfg_dout283            ),
      .cfg_out284          (cfg_dout284            ),
      .cfg_out285          (cfg_dout285            ),
      .cfg_out286          (cfg_dout286            ),
      .cfg_out287          (cfg_dout287            ),
      .cfg_out288          (cfg_dout288            ),
      .cfg_out289          (cfg_dout289            ),
      .cfg_out290          (cfg_dout290            ),
      .cfg_out291          (cfg_dout291            ),
      .cfg_out292          (cfg_dout292            ),
      .cfg_out293          (cfg_dout293            ),
      .cfg_out294          (cfg_dout294            ),
      .cfg_out295          (cfg_dout295            ),
      .cfg_out296          (cfg_dout296            ),
      .cfg_out297          (cfg_dout297            ),
      .cfg_out298          (cfg_dout298            ),
      .cfg_out299          (cfg_dout299            ),
      .cfg_out300          (cfg_dout300            ),
      .cfg_out301          (cfg_dout301            ),
      .cfg_out302          (cfg_dout302            ),
      .cfg_out303          (cfg_dout303            ),
      .cfg_out304          (cfg_dout304            ),
      .cfg_out305          (cfg_dout305            ),
      .cfg_out306          (cfg_dout306            ),
      .cfg_out307          (cfg_dout307            ),
      .cfg_out308          (cfg_dout308            ),
      .cfg_out309          (cfg_dout309            ),
      .cfg_out310          (cfg_dout310            ),
      .cfg_out311          (cfg_dout311            ),
      .cfg_out312          (cfg_dout312            ),
      .cfg_out313          (cfg_dout313            ),
      .cfg_out314          (cfg_dout314            ),
      .cfg_out315          (cfg_dout315            ),
      .cfg_out316          (cfg_dout316            ),
      .cfg_out317          (cfg_dout317            ),
      .cfg_out318          (cfg_dout318            ),
      .cfg_out319          (cfg_dout319            ),
      .cfg_out320          (cfg_dout320            ),
      .cfg_out321          (cfg_dout321            ),
      .cfg_out322          (cfg_dout322            ),
      .cfg_out323          (cfg_dout323            ),
      .cfg_out324          (cfg_dout324            ),
      .cfg_out325          (cfg_dout325            ),
      .cfg_out326          (cfg_dout326            ),
      .cfg_out327          (cfg_dout327            ),
      .cfg_out328          (cfg_dout328            ),
      .cfg_out329          (cfg_dout329            ),
      .cfg_out330          (cfg_dout330            ),
      .cfg_out331          (cfg_dout331            ),
      .cfg_out332          (cfg_dout332            ),
      .cfg_out333          (cfg_dout333            ),
      .cfg_out334          (cfg_dout334            ),
      .cfg_out335          (cfg_dout335            ),
      .cfg_out336          (cfg_dout336            ),
      .cfg_out337          (cfg_dout337            ),
      .cfg_out338          (cfg_dout338            ),
      .cfg_out339          (cfg_dout339            ),
      .cfg_out340          (cfg_dout340            ),
      .cfg_out341          (cfg_dout341            ),
      .cfg_out342          (cfg_dout342            ),
      .cfg_out343          (cfg_dout343            ),
      .cfg_out344          (cfg_dout344            ),
      .cfg_out345          (cfg_dout345            ),
      .cfg_out346          (cfg_dout346            ),
      .cfg_out347          (cfg_dout347            ),
      .cfg_out348          (cfg_dout348            ),
      .cfg_out349          (cfg_dout349            ),
      .cfg_out350          (cfg_dout350            ),
      .cfg_out351          (cfg_dout351            ),
      .cfg_out352          (cfg_dout352            ),
      .cfg_out353          (cfg_dout353            ),
      .cfg_out354          (cfg_dout354            ),
      .cfg_out355          (cfg_dout355            ),
      .cfg_out356          (cfg_dout356            ),
      .cfg_out357          (cfg_dout357            ),
      .cfg_out358          (cfg_dout358            ),
      .cfg_out359          (cfg_dout359            ),
      .cfg_out360          (cfg_dout360            ),
      .cfg_out361          (cfg_dout361            ),
      .cfg_out362          (cfg_dout362            ),
      .cfg_out363          (cfg_dout363            ),
      .cfg_out364          (cfg_dout364            ),
      .cfg_out365          (cfg_dout365            ),
      .cfg_out366          (cfg_dout366            ),
      .cfg_out367          (cfg_dout367            ),
      .cfg_out368          (cfg_dout368            ),
      .cfg_out369          (cfg_dout369            ),
      .cfg_out370          (cfg_dout370            ),
      .cfg_out371          (cfg_dout371            ),
      .cfg_out372          (cfg_dout372            ),
      .cfg_out373          (cfg_dout373            ),
      .cfg_out374          (cfg_dout374            ),
      .cfg_out375          (cfg_dout375            ),
      .cfg_out376          (cfg_dout376            ),
      .cfg_out377          (cfg_dout377            ),
      .cfg_out378          (cfg_dout378            ),
      .cfg_out379          (cfg_dout379            ),
      .cfg_out380          (cfg_dout380            ),
      .cfg_out381          (cfg_dout381            ),
      .cfg_out382          (cfg_dout382            ),
      .cfg_out383          (cfg_dout383            ),
      .cfg_out384          (cfg_dout384            ),
      .cfg_out385          (cfg_dout385            ),
      .cfg_out386          (cfg_dout386            ),
      .cfg_out387          (cfg_dout387            ),
      .cfg_out388          (cfg_dout388            ),
      .cfg_out389          (cfg_dout389            ),
      .cfg_out390          (cfg_dout390            ),
      .cfg_out391          (cfg_dout391            ),
      .cfg_out392          (cfg_dout392            ),
      .cfg_out393          (cfg_dout393            ),
      .cfg_out394          (cfg_dout394            ),
      .cfg_out395          (cfg_dout395            ),
      .cfg_out396          (cfg_dout396            ),
      .cfg_out397          (cfg_dout397            ),
      .cfg_out398          (cfg_dout398            ),
      .cfg_out399          (cfg_dout399            ),
      .cfg_out400          (cfg_dout400            ),
      .cfg_out401          (cfg_dout401            ),
      .cfg_out402          (cfg_dout402            ),
      .cfg_out403          (cfg_dout403            ),
      .cfg_out404          (cfg_dout404            ),
      .cfg_out405          (cfg_dout405            ),
      .cfg_out406          (cfg_dout406            ),
      .cfg_out407          (cfg_dout407            ),
      .cfg_out408          (cfg_dout408            ),
      .cfg_out409          (cfg_dout409            ),
      .cfg_out410          (cfg_dout410            ),
      .cfg_out411          (cfg_dout411            ),
      .cfg_out412          (cfg_dout412            ),
      .cfg_out413          (cfg_dout413            ),
      .cfg_out414          (cfg_dout414            ),
      .cfg_out415          (cfg_dout415            ),
      .cfg_out416          (cfg_dout416            ),
      .cfg_out417          (cfg_dout417            ),
      .cfg_out418          (cfg_dout418            ),
      .cfg_out419          (cfg_dout419            ),
      .cfg_out420          (cfg_dout420            ),
      .cfg_out421          (cfg_dout421            ),
      .cfg_out422          (cfg_dout422            ),
      .cfg_out423          (cfg_dout423            ),
      .cfg_out424          (cfg_dout424            ),
      .cfg_out425          (cfg_dout425            ),
      .cfg_out426          (cfg_dout426            ),
      .cfg_out427          (cfg_dout427            ),
      .cfg_out428          (cfg_dout428            ),
      .cfg_out429          (cfg_dout429            ),
      .cfg_out430          (cfg_dout430            ),
      .cfg_out431          (cfg_dout431            ),
      .cfg_out432          (cfg_dout432            ),
      .cfg_out433          (cfg_dout433            ),
      .cfg_out434          (cfg_dout434            ),
      .cfg_out435          (cfg_dout435            ),
      .cfg_out436          (cfg_dout436            ),
      .cfg_out437          (cfg_dout437            ),
      .cfg_out438          (cfg_dout438            ),
      .cfg_out439          (cfg_dout439            ),
      .cfg_out440          (cfg_dout440            ),
      .cfg_out441          (cfg_dout441            ),
      .cfg_out442          (cfg_dout442            ),
      .cfg_out443          (cfg_dout443            ),
      .cfg_out444          (cfg_dout444            ),
      .cfg_out445          (cfg_dout445            ),
      .cfg_out446          (cfg_dout446            ),
      .cfg_out447          (cfg_dout447            ),
      .cfg_out448          (cfg_dout448            ),
      .cfg_out449          (cfg_dout449            ),
      .cfg_out450          (cfg_dout450            ),
      .cfg_out451          (cfg_dout451            ),
      .cfg_out452          (cfg_dout452            ),
      .cfg_out453          (cfg_dout453            ),
      .cfg_out454          (cfg_dout454            ),
      .cfg_out455          (cfg_dout455            ),
      .cfg_out456          (cfg_dout456            ),
      .cfg_out457          (cfg_dout457            ),
      .cfg_out458          (cfg_dout458            ),
      .cfg_out459          (cfg_dout459            ),
      .cfg_out460          (cfg_dout460            ),
      .cfg_out461          (cfg_dout461            ),
      .cfg_out462          (cfg_dout462            ),
      .cfg_out463          (cfg_dout463            ),
      .cfg_out464          (cfg_dout464            ),
      .cfg_out465          (cfg_dout465            ),
      .cfg_out466          (cfg_dout466            ),
      .cfg_out467          (cfg_dout467            ),
      .cfg_out468          (cfg_dout468            ),
      .cfg_out469          (cfg_dout469            ),
      .cfg_out470          (cfg_dout470            ),
      .cfg_out471          (cfg_dout471            ),
      .cfg_out472          (cfg_dout472            ),
      .cfg_out473          (cfg_dout473            ),
      .cfg_out474          (cfg_dout474            ),
      .cfg_out475          (cfg_dout475            ),
      .cfg_out476          (cfg_dout476            ),
      .cfg_out477          (cfg_dout477            ),
      .cfg_out478          (cfg_dout478            ),
      .cfg_out479          (cfg_dout479            ),
      .cfg_out480          (cfg_dout480            ),
      .cfg_out481          (cfg_dout481            ),
      .cfg_out482          (cfg_dout482            ),
      .cfg_out483          (cfg_dout483            ),
      .cfg_out484          (cfg_dout484            ),
      .cfg_out485          (cfg_dout485            ),
      .cfg_out486          (cfg_dout486            ),
      .cfg_out487          (cfg_dout487            ),
      .cfg_out488          (cfg_dout488            ),
      .cfg_out489          (cfg_dout489            ),
      .cfg_out490          (cfg_dout490            ),
      .cfg_out491          (cfg_dout491            ),
      .cfg_out492          (cfg_dout492            ),
      .cfg_out493          (cfg_dout493            ),
      .cfg_out494          (cfg_dout494            ),
      .cfg_out495          (cfg_dout495            ),
      .cfg_out496          (cfg_dout496            ),
      .cfg_out497          (cfg_dout497            ),
      .cfg_out498          (cfg_dout498            ),
      .cfg_out499          (cfg_dout499            ),
      .cfg_out500          (cfg_dout500            ),
      .cfg_out501          (cfg_dout501            ),
      .cfg_out502          (cfg_dout502            ),
      .cfg_out503          (cfg_dout503            ),
      .cfg_out504          (cfg_dout504            ),
      .cfg_out505          (cfg_dout505            ),
      .cfg_out506          (cfg_dout506            ),
      .cfg_out507          (cfg_dout507            ),
      .cfg_out508          (cfg_dout508            ),
      .cfg_out509          (cfg_dout509            ),
      .cfg_out510          (cfg_dout510            ),
      .cfg_out511          (cfg_dout511            ),
      .cfg_in0           (cfg_din0             ),
      .cfg_in1           (cfg_din1             ),
      .cfg_in2           (cfg_din2             ),
      .cfg_in3           (cfg_din3             ),
      .cfg_in4           (cfg_din4             ),
      .cfg_in5           (cfg_din5             ),
      .cfg_in6           (cfg_din6             ),
      .cfg_in7           (cfg_din7             ),
      .cfg_in8           (cfg_din8             ),
      .cfg_in9           (cfg_din9             ),
      .cfg_in10           (cfg_din10             ),
      .cfg_in11           (cfg_din11             ),
      .cfg_in12           (cfg_din12             ),
      .cfg_in13           (cfg_din13             ),
      .cfg_in14           (cfg_din14             ),
      .cfg_in15           (cfg_din15             ),
      .cfg_in16           (cfg_din16             ),
      .cfg_in17           (cfg_din17             ),
      .cfg_in18           (cfg_din18             ),
      .cfg_in19           (cfg_din19             ),
      .cfg_in20           (cfg_din20             ),
      .cfg_in21           (cfg_din21             ),
      .cfg_in22           (cfg_din22             ),
      .cfg_in23           (cfg_din23             ),
      .cfg_in24           (cfg_din24             ),
      .cfg_in25           (cfg_din25             ),
      .cfg_in26           (cfg_din26             ),
      .cfg_in27           (cfg_din27             ),
      .cfg_in28           (cfg_din28             ),
      .cfg_in29           (cfg_din29             ),
      .cfg_in30           (cfg_din30             ),
      .cfg_in31           (cfg_din31             ),
      .cfg_in32           (cfg_din32             ),
      .cfg_in33           (cfg_din33             ),
      .cfg_in34           (cfg_din34             ),
      .cfg_in35           (cfg_din35             ),
      .cfg_in36           (cfg_din36             ),
      .cfg_in37           (cfg_din37             ),
      .cfg_in38           (cfg_din38             ),
      .cfg_in39           (cfg_din39             ),
      .cfg_in40           (cfg_din40             ),
      .cfg_in41           (cfg_din41             ),
      .cfg_in42           (cfg_din42             ),
      .cfg_in43           (cfg_din43             ),
      .cfg_in44           (cfg_din44             ),
      .cfg_in45           (cfg_din45             ),
      .cfg_in46           (cfg_din46             ),
      .cfg_in47           (cfg_din47             ),
      .cfg_in48           (cfg_din48             ),
      .cfg_in49           (cfg_din49             ),
      .cfg_in50           (cfg_din50             ),
      .cfg_in51           (cfg_din51             ),
      .cfg_in52           (cfg_din52             ),
      .cfg_in53           (cfg_din53             ),
      .cfg_in54           (cfg_din54             ),
      .cfg_in55           (cfg_din55             ),
      .cfg_in56           (cfg_din56             ),
      .cfg_in57           (cfg_din57             ),
      .cfg_in58           (cfg_din58             ),
      .cfg_in59           (cfg_din59             ),
      .cfg_in60           (cfg_din60             ),
      .cfg_in61           (cfg_din61             ),
      .cfg_in62           (cfg_din62             ),
      .cfg_in63           (cfg_din63             ),
      .cfg_in64           (cfg_din64             ),
      .cfg_in65           (cfg_din65             ),
      .cfg_in66           (cfg_din66             ),
      .cfg_in67           (cfg_din67             ),
      .cfg_in68           (cfg_din68             ),
      .cfg_in69           (cfg_din69             ),
      .cfg_in70           (cfg_din70             ),
      .cfg_in71           (cfg_din71             ),
      .cfg_in72           (cfg_din72             ),
      .cfg_in73           (cfg_din73             ),
      .cfg_in74           (cfg_din74             ),
      .cfg_in75           (cfg_din75             ),
      .cfg_in76           (cfg_din76             ),
      .cfg_in77           (cfg_din77             ),
      .cfg_in78           (cfg_din78             ),
      .cfg_in79           (cfg_din79             ),
      .cfg_in80           (cfg_din80             ),
      .cfg_in81           (cfg_din81             ),
      .cfg_in82           (cfg_din82             ),
      .cfg_in83           (cfg_din83             ),
      .cfg_in84           (cfg_din84             ),
      .cfg_in85           (cfg_din85             ),
      .cfg_in86           (cfg_din86             ),
      .cfg_in87           (cfg_din87             ),
      .cfg_in88           (cfg_din88             ),
      .cfg_in89           (cfg_din89             ),
      .cfg_in90           (cfg_din90             ),
      .cfg_in91           (cfg_din91             ),
      .cfg_in92           (cfg_din92             ),
      .cfg_in93           (cfg_din93             ),
      .cfg_in94           (cfg_din94             ),
      .cfg_in95           (cfg_din95             ),
      .cfg_in96           (cfg_din96             ),
      .cfg_in97           (cfg_din97             ),
      .cfg_in98           (cfg_din98             ),
      .cfg_in99           (cfg_din99             ),
      .cfg_in100           (cfg_din100             ),
      .cfg_in101           (cfg_din101             ),
      .cfg_in102           (cfg_din102             ),
      .cfg_in103           (cfg_din103             ),
      .cfg_in104           (cfg_din104             ),
      .cfg_in105           (cfg_din105             ),
      .cfg_in106           (cfg_din106             ),
      .cfg_in107           (cfg_din107             ),
      .cfg_in108           (cfg_din108             ),
      .cfg_in109           (cfg_din109             ),
      .cfg_in110           (cfg_din110             ),
      .cfg_in111           (cfg_din111             ),
      .cfg_in112           (cfg_din112             ),
      .cfg_in113           (cfg_din113             ),
      .cfg_in114           (cfg_din114             ),
      .cfg_in115           (cfg_din115             ),
      .cfg_in116           (cfg_din116             ),
      .cfg_in117           (cfg_din117             ),
      .cfg_in118           (cfg_din118             ),
      .cfg_in119           (cfg_din119             ),
      .cfg_in120           (cfg_din120             ),
      .cfg_in121           (cfg_din121             ),
      .cfg_in122           (cfg_din122             ),
      .cfg_in123           (cfg_din123             ),
      .cfg_in124           (cfg_din124             ),
      .cfg_in125           (cfg_din125             ),
      .cfg_in126           (cfg_din126             ),
      .cfg_in127           (cfg_din127             ),
      .cfg_in128           (cfg_din128             ),
      .cfg_in129           (cfg_din129             ),
      .cfg_in130           (cfg_din130             ),
      .cfg_in131           (cfg_din131             ),
      .cfg_in132           (cfg_din132             ),
      .cfg_in133           (cfg_din133             ),
      .cfg_in134           (cfg_din134             ),
      .cfg_in135           (cfg_din135             ),
      .cfg_in136           (cfg_din136             ),
      .cfg_in137           (cfg_din137             ),
      .cfg_in138           (cfg_din138             ),
      .cfg_in139           (cfg_din139             ),
      .cfg_in140           (cfg_din140             ),
      .cfg_in141           (cfg_din141             ),
      .cfg_in142           (cfg_din142             ),
      .cfg_in143           (cfg_din143             ),
      .cfg_in144           (cfg_din144             ),
      .cfg_in145           (cfg_din145             ),
      .cfg_in146           (cfg_din146             ),
      .cfg_in147           (cfg_din147             ),
      .cfg_in148           (cfg_din148             ),
      .cfg_in149           (cfg_din149             ),
      .cfg_in150           (cfg_din150             ),
      .cfg_in151           (cfg_din151             ),
      .cfg_in152           (cfg_din152             ),
      .cfg_in153           (cfg_din153             ),
      .cfg_in154           (cfg_din154             ),
      .cfg_in155           (cfg_din155             ),
      .cfg_in156           (cfg_din156             ),
      .cfg_in157           (cfg_din157             ),
      .cfg_in158           (cfg_din158             ),
      .cfg_in159           (cfg_din159             ),
      .cfg_in160           (cfg_din160             ),
      .cfg_in161           (cfg_din161             ),
      .cfg_in162           (cfg_din162             ),
      .cfg_in163           (cfg_din163             ),
      .cfg_in164           (cfg_din164             ),
      .cfg_in165           (cfg_din165             ),
      .cfg_in166           (cfg_din166             ),
      .cfg_in167           (cfg_din167             ),
      .cfg_in168           (cfg_din168             ),
      .cfg_in169           (cfg_din169             ),
      .cfg_in170           (cfg_din170             ),
      .cfg_in171           (cfg_din171             ),
      .cfg_in172           (cfg_din172             ),
      .cfg_in173           (cfg_din173             ),
      .cfg_in174           (cfg_din174             ),
      .cfg_in175           (cfg_din175             ),
      .cfg_in176           (cfg_din176             ),
      .cfg_in177           (cfg_din177             ),
      .cfg_in178           (cfg_din178             ),
      .cfg_in179           (cfg_din179             ),
      .cfg_in180           (cfg_din180             ),
      .cfg_in181           (cfg_din181             ),
      .cfg_in182           (cfg_din182             ),
      .cfg_in183           (cfg_din183             ),
      .cfg_in184           (cfg_din184             ),
      .cfg_in185           (cfg_din185             ),
      .cfg_in186           (cfg_din186             ),
      .cfg_in187           (cfg_din187             ),
      .cfg_in188           (cfg_din188             ),
      .cfg_in189           (cfg_din189             ),
      .cfg_in190           (cfg_din190             ),
      .cfg_in191           (cfg_din191             ),
      .cfg_in192           (cfg_din192             ),
      .cfg_in193           (cfg_din193             ),
      .cfg_in194           (cfg_din194             ),
      .cfg_in195           (cfg_din195             ),
      .cfg_in196           (cfg_din196             ),
      .cfg_in197           (cfg_din197             ),
      .cfg_in198           (cfg_din198             ),
      .cfg_in199           (cfg_din199             ),
      .cfg_in200           (cfg_din200             ),
      .cfg_in201           (cfg_din201             ),
      .cfg_in202           (cfg_din202             ),
      .cfg_in203           (cfg_din203             ),
      .cfg_in204           (cfg_din204             ),
      .cfg_in205           (cfg_din205             ),
      .cfg_in206           (cfg_din206             ),
      .cfg_in207           (cfg_din207             ),
      .cfg_in208           (cfg_din208             ),
      .cfg_in209           (cfg_din209             ),
      .cfg_in210           (cfg_din210             ),
      .cfg_in211           (cfg_din211             ),
      .cfg_in212           (cfg_din212             ),
      .cfg_in213           (cfg_din213             ),
      .cfg_in214           (cfg_din214             ),
      .cfg_in215           (cfg_din215             ),
      .cfg_in216           (cfg_din216             ),
      .cfg_in217           (cfg_din217             ),
      .cfg_in218           (cfg_din218             ),
      .cfg_in219           (cfg_din219             ),
      .cfg_in220           (cfg_din220             ),
      .cfg_in221           (cfg_din221             ),
      .cfg_in222           (cfg_din222             ),
      .cfg_in223           (cfg_din223             ),
      .cfg_in224           (cfg_din224             ),
      .cfg_in225           (cfg_din225             ),
      .cfg_in226           (cfg_din226             ),
      .cfg_in227           (cfg_din227             ),
      .cfg_in228           (cfg_din228             ),
      .cfg_in229           (cfg_din229             ),
      .cfg_in230           (cfg_din230             ),
      .cfg_in231           (cfg_din231             ),
      .cfg_in232           (cfg_din232             ),
      .cfg_in233           (cfg_din233             ),
      .cfg_in234           (cfg_din234             ),
      .cfg_in235           (cfg_din235             ),
      .cfg_in236           (cfg_din236             ),
      .cfg_in237           (cfg_din237             ),
      .cfg_in238           (cfg_din238             ),
      .cfg_in239           (cfg_din239             ),
      .cfg_in240           (cfg_din240             ),
      .cfg_in241           (cfg_din241             ),
      .cfg_in242           (cfg_din242             ),
      .cfg_in243           (cfg_din243             ),
      .cfg_in244           (cfg_din244             ),
      .cfg_in245           (cfg_din245             ),
      .cfg_in246           (cfg_din246             ),
      .cfg_in247           (cfg_din247             ),
      .cfg_in248           (cfg_din248             ),
      .cfg_in249           (cfg_din249             ),
      .cfg_in250           (cfg_din250             ),
      .cfg_in251           (cfg_din251             ),
      .cfg_in252           (cfg_din252             ),
      .cfg_in253           (cfg_din253             ),
      .cfg_in254           (cfg_din254             ),
      .cfg_in255           (cfg_din255             ),
      .cfg_in256           (cfg_din256             ),
      .cfg_in257           (cfg_din257             ),
      .cfg_in258           (cfg_din258             ),
      .cfg_in259           (cfg_din259             ),
      .cfg_in260           (cfg_din260             ),
      .cfg_in261           (cfg_din261             ),
      .cfg_in262           (cfg_din262             ),
      .cfg_in263           (cfg_din263             ),
      .cfg_in264           (cfg_din264             ),
      .cfg_in265           (cfg_din265             ),
      .cfg_in266           (cfg_din266             ),
      .cfg_in267           (cfg_din267             ),
      .cfg_in268           (cfg_din268             ),
      .cfg_in269           (cfg_din269             ),
      .cfg_in270           (cfg_din270             ),
      .cfg_in271           (cfg_din271             ),
      .cfg_in272           (cfg_din272             ),
      .cfg_in273           (cfg_din273             ),
      .cfg_in274           (cfg_din274             ),
      .cfg_in275           (cfg_din275             ),
      .cfg_in276           (cfg_din276             ),
      .cfg_in277           (cfg_din277             ),
      .cfg_in278           (cfg_din278             ),
      .cfg_in279           (cfg_din279             ),
      .cfg_in280           (cfg_din280             ),
      .cfg_in281           (cfg_din281             ),
      .cfg_in282           (cfg_din282             ),
      .cfg_in283           (cfg_din283             ),
      .cfg_in284           (cfg_din284             ),
      .cfg_in285           (cfg_din285             ),
      .cfg_in286           (cfg_din286             ),
      .cfg_in287           (cfg_din287             ),
      .cfg_in288           (cfg_din288             ),
      .cfg_in289           (cfg_din289             ),
      .cfg_in290           (cfg_din290             ),
      .cfg_in291           (cfg_din291             ),
      .cfg_in292           (cfg_din292             ),
      .cfg_in293           (cfg_din293             ),
      .cfg_in294           (cfg_din294             ),
      .cfg_in295           (cfg_din295             ),
      .cfg_in296           (cfg_din296             ),
      .cfg_in297           (cfg_din297             ),
      .cfg_in298           (cfg_din298             ),
      .cfg_in299           (cfg_din299             ),
      .cfg_in300           (cfg_din300             ),
      .cfg_in301           (cfg_din301             ),
      .cfg_in302           (cfg_din302             ),
      .cfg_in303           (cfg_din303             ),
      .cfg_in304           (cfg_din304             ),
      .cfg_in305           (cfg_din305             ),
      .cfg_in306           (cfg_din306             ),
      .cfg_in307           (cfg_din307             ),
      .cfg_in308           (cfg_din308             ),
      .cfg_in309           (cfg_din309             ),
      .cfg_in310           (cfg_din310             ),
      .cfg_in311           (cfg_din311             ),
      .cfg_in312           (cfg_din312             ),
      .cfg_in313           (cfg_din313             ),
      .cfg_in314           (cfg_din314             ),
      .cfg_in315           (cfg_din315             ),
      .cfg_in316           (cfg_din316             ),
      .cfg_in317           (cfg_din317             ),
      .cfg_in318           (cfg_din318             ),
      .cfg_in319           (cfg_din319             ),
      .cfg_in320           (cfg_din320             ),
      .cfg_in321           (cfg_din321             ),
      .cfg_in322           (cfg_din322             ),
      .cfg_in323           (cfg_din323             ),
      .cfg_in324           (cfg_din324             ),
      .cfg_in325           (cfg_din325             ),
      .cfg_in326           (cfg_din326             ),
      .cfg_in327           (cfg_din327             ),
      .cfg_in328           (cfg_din328             ),
      .cfg_in329           (cfg_din329             ),
      .cfg_in330           (cfg_din330             ),
      .cfg_in331           (cfg_din331             ),
      .cfg_in332           (cfg_din332             ),
      .cfg_in333           (cfg_din333             ),
      .cfg_in334           (cfg_din334             ),
      .cfg_in335           (cfg_din335             ),
      .cfg_in336           (cfg_din336             ),
      .cfg_in337           (cfg_din337             ),
      .cfg_in338           (cfg_din338             ),
      .cfg_in339           (cfg_din339             ),
      .cfg_in340           (cfg_din340             ),
      .cfg_in341           (cfg_din341             ),
      .cfg_in342           (cfg_din342             ),
      .cfg_in343           (cfg_din343             ),
      .cfg_in344           (cfg_din344             ),
      .cfg_in345           (cfg_din345             ),
      .cfg_in346           (cfg_din346             ),
      .cfg_in347           (cfg_din347             ),
      .cfg_in348           (cfg_din348             ),
      .cfg_in349           (cfg_din349             ),
      .cfg_in350           (cfg_din350             ),
      .cfg_in351           (cfg_din351             ),
      .cfg_in352           (cfg_din352             ),
      .cfg_in353           (cfg_din353             ),
      .cfg_in354           (cfg_din354             ),
      .cfg_in355           (cfg_din355             ),
      .cfg_in356           (cfg_din356             ),
      .cfg_in357           (cfg_din357             ),
      .cfg_in358           (cfg_din358             ),
      .cfg_in359           (cfg_din359             ),
      .cfg_in360           (cfg_din360             ),
      .cfg_in361           (cfg_din361             ),
      .cfg_in362           (cfg_din362             ),
      .cfg_in363           (cfg_din363             ),
      .cfg_in364           (cfg_din364             ),
      .cfg_in365           (cfg_din365             ),
      .cfg_in366           (cfg_din366             ),
      .cfg_in367           (cfg_din367             ),
      .cfg_in368           (cfg_din368             ),
      .cfg_in369           (cfg_din369             ),
      .cfg_in370           (cfg_din370             ),
      .cfg_in371           (cfg_din371             ),
      .cfg_in372           (cfg_din372             ),
      .cfg_in373           (cfg_din373             ),
      .cfg_in374           (cfg_din374             ),
      .cfg_in375           (cfg_din375             ),
      .cfg_in376           (cfg_din376             ),
      .cfg_in377           (cfg_din377             ),
      .cfg_in378           (cfg_din378             ),
      .cfg_in379           (cfg_din379             ),
      .cfg_in380           (cfg_din380             ),
      .cfg_in381           (cfg_din381             ),
      .cfg_in382           (cfg_din382             ),
      .cfg_in383           (cfg_din383             ),
      .cfg_in384           (cfg_din384             ),
      .cfg_in385           (cfg_din385             ),
      .cfg_in386           (cfg_din386             ),
      .cfg_in387           (cfg_din387             ),
      .cfg_in388           (cfg_din388             ),
      .cfg_in389           (cfg_din389             ),
      .cfg_in390           (cfg_din390             ),
      .cfg_in391           (cfg_din391             ),
      .cfg_in392           (cfg_din392             ),
      .cfg_in393           (cfg_din393             ),
      .cfg_in394           (cfg_din394             ),
      .cfg_in395           (cfg_din395             ),
      .cfg_in396           (cfg_din396             ),
      .cfg_in397           (cfg_din397             ),
      .cfg_in398           (cfg_din398             ),
      .cfg_in399           (cfg_din399             ),
      .cfg_in400           (cfg_din400             ),
      .cfg_in401           (cfg_din401             ),
      .cfg_in402           (cfg_din402             ),
      .cfg_in403           (cfg_din403             ),
      .cfg_in404           (cfg_din404             ),
      .cfg_in405           (cfg_din405             ),
      .cfg_in406           (cfg_din406             ),
      .cfg_in407           (cfg_din407             ),
      .cfg_in408           (cfg_din408             ),
      .cfg_in409           (cfg_din409             ),
      .cfg_in410           (cfg_din410             ),
      .cfg_in411           (cfg_din411             ),
      .cfg_in412           (cfg_din412             ),
      .cfg_in413           (cfg_din413             ),
      .cfg_in414           (cfg_din414             ),
      .cfg_in415           (cfg_din415             ),
      .cfg_in416           (cfg_din416             ),
      .cfg_in417           (cfg_din417             ),
      .cfg_in418           (cfg_din418             ),
      .cfg_in419           (cfg_din419             ),
      .cfg_in420           (cfg_din420             ),
      .cfg_in421           (cfg_din421             ),
      .cfg_in422           (cfg_din422             ),
      .cfg_in423           (cfg_din423             ),
      .cfg_in424           (cfg_din424             ),
      .cfg_in425           (cfg_din425             ),
      .cfg_in426           (cfg_din426             ),
      .cfg_in427           (cfg_din427             ),
      .cfg_in428           (cfg_din428             ),
      .cfg_in429           (cfg_din429             ),
      .cfg_in430           (cfg_din430             ),
      .cfg_in431           (cfg_din431             ),
      .cfg_in432           (cfg_din432             ),
      .cfg_in433           (cfg_din433             ),
      .cfg_in434           (cfg_din434             ),
      .cfg_in435           (cfg_din435             ),
      .cfg_in436           (cfg_din436             ),
      .cfg_in437           (cfg_din437             ),
      .cfg_in438           (cfg_din438             ),
      .cfg_in439           (cfg_din439             ),
      .cfg_in440           (cfg_din440             ),
      .cfg_in441           (cfg_din441             ),
      .cfg_in442           (cfg_din442             ),
      .cfg_in443           (cfg_din443             ),
      .cfg_in444           (cfg_din444             ),
      .cfg_in445           (cfg_din445             ),
      .cfg_in446           (cfg_din446             ),
      .cfg_in447           (cfg_din447             ),
      .cfg_in448           (cfg_din448             ),
      .cfg_in449           (cfg_din449             ),
      .cfg_in450           (cfg_din450             ),
      .cfg_in451           (cfg_din451             ),
      .cfg_in452           (cfg_din452             ),
      .cfg_in453           (cfg_din453             ),
      .cfg_in454           (cfg_din454             ),
      .cfg_in455           (cfg_din455             ),
      .cfg_in456           (cfg_din456             ),
      .cfg_in457           (cfg_din457             ),
      .cfg_in458           (cfg_din458             ),
      .cfg_in459           (cfg_din459             ),
      .cfg_in460           (cfg_din460             ),
      .cfg_in461           (cfg_din461             ),
      .cfg_in462           (cfg_din462             ),
      .cfg_in463           (cfg_din463             ),
      .cfg_in464           (cfg_din464             ),
      .cfg_in465           (cfg_din465             ),
      .cfg_in466           (cfg_din466             ),
      .cfg_in467           (cfg_din467             ),
      .cfg_in468           (cfg_din468             ),
      .cfg_in469           (cfg_din469             ),
      .cfg_in470           (cfg_din470             ),
      .cfg_in471           (cfg_din471             ),
      .cfg_in472           (cfg_din472             ),
      .cfg_in473           (cfg_din473             ),
      .cfg_in474           (cfg_din474             ),
      .cfg_in475           (cfg_din475             ),
      .cfg_in476           (cfg_din476             ),
      .cfg_in477           (cfg_din477             ),
      .cfg_in478           (cfg_din478             ),
      .cfg_in479           (cfg_din479             ),
      .cfg_in480           (cfg_din480             ),
      .cfg_in481           (cfg_din481             ),
      .cfg_in482           (cfg_din482             ),
      .cfg_in483           (cfg_din483             ),
      .cfg_in484           (cfg_din484             ),
      .cfg_in485           (cfg_din485             ),
      .cfg_in486           (cfg_din486             ),
      .cfg_in487           (cfg_din487             ),
      .cfg_in488           (cfg_din488             ),
      .cfg_in489           (cfg_din489             ),
      .cfg_in490           (cfg_din490             ),
      .cfg_in491           (cfg_din491             ),
      .cfg_in492           (cfg_din492             ),
      .cfg_in493           (cfg_din493             ),
      .cfg_in494           (cfg_din494             ),
      .cfg_in495           (cfg_din495             ),
      .cfg_in496           (cfg_din496             ),
      .cfg_in497           (cfg_din497             ),
      .cfg_in498           (cfg_din498             ),
      .cfg_in499           (cfg_din499             ),
      .cfg_in500           (cfg_din500             ),
      .cfg_in501           (cfg_din501             ),
      .cfg_in502           (cfg_din502             ),
      .cfg_in503           (cfg_din503             ),
      .cfg_in504           (cfg_din504             ),
      .cfg_in505           (cfg_din505             ),
      .cfg_in506           (cfg_din506             ),
      .cfg_in507           (cfg_din507             ),
      .cfg_in508           (cfg_din508             ),
      .cfg_in509           (cfg_din509             ),
      .cfg_in510           (cfg_din510             ),
      .cfg_in511           (cfg_din511             ),
      .cfg_en0           (cfg_en0              ),
      .cfg_en1           (cfg_en1              ),
      .cfg_en2           (cfg_en2              ),
      .cfg_en3           (cfg_en3              ),
      .cfg_en4           (cfg_en4              ),
      .cfg_en5           (cfg_en5              ),
      .cfg_en6           (cfg_en6              ),
      .cfg_en7           (cfg_en7              ),
      .cfg_en8           (cfg_en8              ),
      .cfg_en9           (cfg_en9              ),
      .cfg_en10           (cfg_en10              ),
      .cfg_en11           (cfg_en11              ),
      .cfg_en12           (cfg_en12              ),
      .cfg_en13           (cfg_en13              ),
      .cfg_en14           (cfg_en14              ),
      .cfg_en15           (cfg_en15              ),
      .cfg_en16           (cfg_en16              ),
      .cfg_en17           (cfg_en17              ),
      .cfg_en18           (cfg_en18              ),
      .cfg_en19           (cfg_en19              ),
      .cfg_en20           (cfg_en20              ),
      .cfg_en21           (cfg_en21              ),
      .cfg_en22           (cfg_en22              ),
      .cfg_en23           (cfg_en23              ),
      .cfg_en24           (cfg_en24              ),
      .cfg_en25           (cfg_en25              ),
      .cfg_en26           (cfg_en26              ),
      .cfg_en27           (cfg_en27              ),
      .cfg_en28           (cfg_en28              ),
      .cfg_en29           (cfg_en29              ),
      .cfg_en30           (cfg_en30              ),
      .cfg_en31           (cfg_en31              ),
      .cfg_en32           (cfg_en32              ),
      .cfg_en33           (cfg_en33              ),
      .cfg_en34           (cfg_en34              ),
      .cfg_en35           (cfg_en35              ),
      .cfg_en36           (cfg_en36              ),
      .cfg_en37           (cfg_en37              ),
      .cfg_en38           (cfg_en38              ),
      .cfg_en39           (cfg_en39              ),
      .cfg_en40           (cfg_en40              ),
      .cfg_en41           (cfg_en41              ),
      .cfg_en42           (cfg_en42              ),
      .cfg_en43           (cfg_en43              ),
      .cfg_en44           (cfg_en44              ),
      .cfg_en45           (cfg_en45              ),
      .cfg_en46           (cfg_en46              ),
      .cfg_en47           (cfg_en47              ),
      .cfg_en48           (cfg_en48              ),
      .cfg_en49           (cfg_en49              ),
      .cfg_en50           (cfg_en50              ),
      .cfg_en51           (cfg_en51              ),
      .cfg_en52           (cfg_en52              ),
      .cfg_en53           (cfg_en53              ),
      .cfg_en54           (cfg_en54              ),
      .cfg_en55           (cfg_en55              ),
      .cfg_en56           (cfg_en56              ),
      .cfg_en57           (cfg_en57              ),
      .cfg_en58           (cfg_en58              ),
      .cfg_en59           (cfg_en59              ),
      .cfg_en60           (cfg_en60              ),
      .cfg_en61           (cfg_en61              ),
      .cfg_en62           (cfg_en62              ),
      .cfg_en63           (cfg_en63              ),
      .cfg_en64           (cfg_en64              ),
      .cfg_en65           (cfg_en65              ),
      .cfg_en66           (cfg_en66              ),
      .cfg_en67           (cfg_en67              ),
      .cfg_en68           (cfg_en68              ),
      .cfg_en69           (cfg_en69              ),
      .cfg_en70           (cfg_en70              ),
      .cfg_en71           (cfg_en71              ),
      .cfg_en72           (cfg_en72              ),
      .cfg_en73           (cfg_en73              ),
      .cfg_en74           (cfg_en74              ),
      .cfg_en75           (cfg_en75              ),
      .cfg_en76           (cfg_en76              ),
      .cfg_en77           (cfg_en77              ),
      .cfg_en78           (cfg_en78              ),
      .cfg_en79           (cfg_en79              ),
      .cfg_en80           (cfg_en80              ),
      .cfg_en81           (cfg_en81              ),
      .cfg_en82           (cfg_en82              ),
      .cfg_en83           (cfg_en83              ),
      .cfg_en84           (cfg_en84              ),
      .cfg_en85           (cfg_en85              ),
      .cfg_en86           (cfg_en86              ),
      .cfg_en87           (cfg_en87              ),
      .cfg_en88           (cfg_en88              ),
      .cfg_en89           (cfg_en89              ),
      .cfg_en90           (cfg_en90              ),
      .cfg_en91           (cfg_en91              ),
      .cfg_en92           (cfg_en92              ),
      .cfg_en93           (cfg_en93              ),
      .cfg_en94           (cfg_en94              ),
      .cfg_en95           (cfg_en95              ),
      .cfg_en96           (cfg_en96              ),
      .cfg_en97           (cfg_en97              ),
      .cfg_en98           (cfg_en98              ),
      .cfg_en99           (cfg_en99              ),
      .cfg_en100           (cfg_en100              ),
      .cfg_en101           (cfg_en101              ),
      .cfg_en102           (cfg_en102              ),
      .cfg_en103           (cfg_en103              ),
      .cfg_en104           (cfg_en104              ),
      .cfg_en105           (cfg_en105              ),
      .cfg_en106           (cfg_en106              ),
      .cfg_en107           (cfg_en107              ),
      .cfg_en108           (cfg_en108              ),
      .cfg_en109           (cfg_en109              ),
      .cfg_en110           (cfg_en110              ),
      .cfg_en111           (cfg_en111              ),
      .cfg_en112           (cfg_en112              ),
      .cfg_en113           (cfg_en113              ),
      .cfg_en114           (cfg_en114              ),
      .cfg_en115           (cfg_en115              ),
      .cfg_en116           (cfg_en116              ),
      .cfg_en117           (cfg_en117              ),
      .cfg_en118           (cfg_en118              ),
      .cfg_en119           (cfg_en119              ),
      .cfg_en120           (cfg_en120              ),
      .cfg_en121           (cfg_en121              ),
      .cfg_en122           (cfg_en122              ),
      .cfg_en123           (cfg_en123              ),
      .cfg_en124           (cfg_en124              ),
      .cfg_en125           (cfg_en125              ),
      .cfg_en126           (cfg_en126              ),
      .cfg_en127           (cfg_en127              ),
      .cfg_en128           (cfg_en128              ),
      .cfg_en129           (cfg_en129              ),
      .cfg_en130           (cfg_en130              ),
      .cfg_en131           (cfg_en131              ),
      .cfg_en132           (cfg_en132              ),
      .cfg_en133           (cfg_en133              ),
      .cfg_en134           (cfg_en134              ),
      .cfg_en135           (cfg_en135              ),
      .cfg_en136           (cfg_en136              ),
      .cfg_en137           (cfg_en137              ),
      .cfg_en138           (cfg_en138              ),
      .cfg_en139           (cfg_en139              ),
      .cfg_en140           (cfg_en140              ),
      .cfg_en141           (cfg_en141              ),
      .cfg_en142           (cfg_en142              ),
      .cfg_en143           (cfg_en143              ),
      .cfg_en144           (cfg_en144              ),
      .cfg_en145           (cfg_en145              ),
      .cfg_en146           (cfg_en146              ),
      .cfg_en147           (cfg_en147              ),
      .cfg_en148           (cfg_en148              ),
      .cfg_en149           (cfg_en149              ),
      .cfg_en150           (cfg_en150              ),
      .cfg_en151           (cfg_en151              ),
      .cfg_en152           (cfg_en152              ),
      .cfg_en153           (cfg_en153              ),
      .cfg_en154           (cfg_en154              ),
      .cfg_en155           (cfg_en155              ),
      .cfg_en156           (cfg_en156              ),
      .cfg_en157           (cfg_en157              ),
      .cfg_en158           (cfg_en158              ),
      .cfg_en159           (cfg_en159              ),
      .cfg_en160           (cfg_en160              ),
      .cfg_en161           (cfg_en161              ),
      .cfg_en162           (cfg_en162              ),
      .cfg_en163           (cfg_en163              ),
      .cfg_en164           (cfg_en164              ),
      .cfg_en165           (cfg_en165              ),
      .cfg_en166           (cfg_en166              ),
      .cfg_en167           (cfg_en167              ),
      .cfg_en168           (cfg_en168              ),
      .cfg_en169           (cfg_en169              ),
      .cfg_en170           (cfg_en170              ),
      .cfg_en171           (cfg_en171              ),
      .cfg_en172           (cfg_en172              ),
      .cfg_en173           (cfg_en173              ),
      .cfg_en174           (cfg_en174              ),
      .cfg_en175           (cfg_en175              ),
      .cfg_en176           (cfg_en176              ),
      .cfg_en177           (cfg_en177              ),
      .cfg_en178           (cfg_en178              ),
      .cfg_en179           (cfg_en179              ),
      .cfg_en180           (cfg_en180              ),
      .cfg_en181           (cfg_en181              ),
      .cfg_en182           (cfg_en182              ),
      .cfg_en183           (cfg_en183              ),
      .cfg_en184           (cfg_en184              ),
      .cfg_en185           (cfg_en185              ),
      .cfg_en186           (cfg_en186              ),
      .cfg_en187           (cfg_en187              ),
      .cfg_en188           (cfg_en188              ),
      .cfg_en189           (cfg_en189              ),
      .cfg_en190           (cfg_en190              ),
      .cfg_en191           (cfg_en191              ),
      .cfg_en192           (cfg_en192              ),
      .cfg_en193           (cfg_en193              ),
      .cfg_en194           (cfg_en194              ),
      .cfg_en195           (cfg_en195              ),
      .cfg_en196           (cfg_en196              ),
      .cfg_en197           (cfg_en197              ),
      .cfg_en198           (cfg_en198              ),
      .cfg_en199           (cfg_en199              ),
      .cfg_en200           (cfg_en200              ),
      .cfg_en201           (cfg_en201              ),
      .cfg_en202           (cfg_en202              ),
      .cfg_en203           (cfg_en203              ),
      .cfg_en204           (cfg_en204              ),
      .cfg_en205           (cfg_en205              ),
      .cfg_en206           (cfg_en206              ),
      .cfg_en207           (cfg_en207              ),
      .cfg_en208           (cfg_en208              ),
      .cfg_en209           (cfg_en209              ),
      .cfg_en210           (cfg_en210              ),
      .cfg_en211           (cfg_en211              ),
      .cfg_en212           (cfg_en212              ),
      .cfg_en213           (cfg_en213              ),
      .cfg_en214           (cfg_en214              ),
      .cfg_en215           (cfg_en215              ),
      .cfg_en216           (cfg_en216              ),
      .cfg_en217           (cfg_en217              ),
      .cfg_en218           (cfg_en218              ),
      .cfg_en219           (cfg_en219              ),
      .cfg_en220           (cfg_en220              ),
      .cfg_en221           (cfg_en221              ),
      .cfg_en222           (cfg_en222              ),
      .cfg_en223           (cfg_en223              ),
      .cfg_en224           (cfg_en224              ),
      .cfg_en225           (cfg_en225              ),
      .cfg_en226           (cfg_en226              ),
      .cfg_en227           (cfg_en227              ),
      .cfg_en228           (cfg_en228              ),
      .cfg_en229           (cfg_en229              ),
      .cfg_en230           (cfg_en230              ),
      .cfg_en231           (cfg_en231              ),
      .cfg_en232           (cfg_en232              ),
      .cfg_en233           (cfg_en233              ),
      .cfg_en234           (cfg_en234              ),
      .cfg_en235           (cfg_en235              ),
      .cfg_en236           (cfg_en236              ),
      .cfg_en237           (cfg_en237              ),
      .cfg_en238           (cfg_en238              ),
      .cfg_en239           (cfg_en239              ),
      .cfg_en240           (cfg_en240              ),
      .cfg_en241           (cfg_en241              ),
      .cfg_en242           (cfg_en242              ),
      .cfg_en243           (cfg_en243              ),
      .cfg_en244           (cfg_en244              ),
      .cfg_en245           (cfg_en245              ),
      .cfg_en246           (cfg_en246              ),
      .cfg_en247           (cfg_en247              ),
      .cfg_en248           (cfg_en248              ),
      .cfg_en249           (cfg_en249              ),
      .cfg_en250           (cfg_en250              ),
      .cfg_en251           (cfg_en251              ),
      .cfg_en252           (cfg_en252              ),
      .cfg_en253           (cfg_en253              ),
      .cfg_en254           (cfg_en254              ),
      .cfg_en255           (cfg_en255              ),
      .cfg_en256           (cfg_en256              ),
      .cfg_en257           (cfg_en257              ),
      .cfg_en258           (cfg_en258              ),
      .cfg_en259           (cfg_en259              ),
      .cfg_en260           (cfg_en260              ),
      .cfg_en261           (cfg_en261              ),
      .cfg_en262           (cfg_en262              ),
      .cfg_en263           (cfg_en263              ),
      .cfg_en264           (cfg_en264              ),
      .cfg_en265           (cfg_en265              ),
      .cfg_en266           (cfg_en266              ),
      .cfg_en267           (cfg_en267              ),
      .cfg_en268           (cfg_en268              ),
      .cfg_en269           (cfg_en269              ),
      .cfg_en270           (cfg_en270              ),
      .cfg_en271           (cfg_en271              ),
      .cfg_en272           (cfg_en272              ),
      .cfg_en273           (cfg_en273              ),
      .cfg_en274           (cfg_en274              ),
      .cfg_en275           (cfg_en275              ),
      .cfg_en276           (cfg_en276              ),
      .cfg_en277           (cfg_en277              ),
      .cfg_en278           (cfg_en278              ),
      .cfg_en279           (cfg_en279              ),
      .cfg_en280           (cfg_en280              ),
      .cfg_en281           (cfg_en281              ),
      .cfg_en282           (cfg_en282              ),
      .cfg_en283           (cfg_en283              ),
      .cfg_en284           (cfg_en284              ),
      .cfg_en285           (cfg_en285              ),
      .cfg_en286           (cfg_en286              ),
      .cfg_en287           (cfg_en287              ),
      .cfg_en288           (cfg_en288              ),
      .cfg_en289           (cfg_en289              ),
      .cfg_en290           (cfg_en290              ),
      .cfg_en291           (cfg_en291              ),
      .cfg_en292           (cfg_en292              ),
      .cfg_en293           (cfg_en293              ),
      .cfg_en294           (cfg_en294              ),
      .cfg_en295           (cfg_en295              ),
      .cfg_en296           (cfg_en296              ),
      .cfg_en297           (cfg_en297              ),
      .cfg_en298           (cfg_en298              ),
      .cfg_en299           (cfg_en299              ),
      .cfg_en300           (cfg_en300              ),
      .cfg_en301           (cfg_en301              ),
      .cfg_en302           (cfg_en302              ),
      .cfg_en303           (cfg_en303              ),
      .cfg_en304           (cfg_en304              ),
      .cfg_en305           (cfg_en305              ),
      .cfg_en306           (cfg_en306              ),
      .cfg_en307           (cfg_en307              ),
      .cfg_en308           (cfg_en308              ),
      .cfg_en309           (cfg_en309              ),
      .cfg_en310           (cfg_en310              ),
      .cfg_en311           (cfg_en311              ),
      .cfg_en312           (cfg_en312              ),
      .cfg_en313           (cfg_en313              ),
      .cfg_en314           (cfg_en314              ),
      .cfg_en315           (cfg_en315              ),
      .cfg_en316           (cfg_en316              ),
      .cfg_en317           (cfg_en317              ),
      .cfg_en318           (cfg_en318              ),
      .cfg_en319           (cfg_en319              ),
      .cfg_en320           (cfg_en320              ),
      .cfg_en321           (cfg_en321              ),
      .cfg_en322           (cfg_en322              ),
      .cfg_en323           (cfg_en323              ),
      .cfg_en324           (cfg_en324              ),
      .cfg_en325           (cfg_en325              ),
      .cfg_en326           (cfg_en326              ),
      .cfg_en327           (cfg_en327              ),
      .cfg_en328           (cfg_en328              ),
      .cfg_en329           (cfg_en329              ),
      .cfg_en330           (cfg_en330              ),
      .cfg_en331           (cfg_en331              ),
      .cfg_en332           (cfg_en332              ),
      .cfg_en333           (cfg_en333              ),
      .cfg_en334           (cfg_en334              ),
      .cfg_en335           (cfg_en335              ),
      .cfg_en336           (cfg_en336              ),
      .cfg_en337           (cfg_en337              ),
      .cfg_en338           (cfg_en338              ),
      .cfg_en339           (cfg_en339              ),
      .cfg_en340           (cfg_en340              ),
      .cfg_en341           (cfg_en341              ),
      .cfg_en342           (cfg_en342              ),
      .cfg_en343           (cfg_en343              ),
      .cfg_en344           (cfg_en344              ),
      .cfg_en345           (cfg_en345              ),
      .cfg_en346           (cfg_en346              ),
      .cfg_en347           (cfg_en347              ),
      .cfg_en348           (cfg_en348              ),
      .cfg_en349           (cfg_en349              ),
      .cfg_en350           (cfg_en350              ),
      .cfg_en351           (cfg_en351              ),
      .cfg_en352           (cfg_en352              ),
      .cfg_en353           (cfg_en353              ),
      .cfg_en354           (cfg_en354              ),
      .cfg_en355           (cfg_en355              ),
      .cfg_en356           (cfg_en356              ),
      .cfg_en357           (cfg_en357              ),
      .cfg_en358           (cfg_en358              ),
      .cfg_en359           (cfg_en359              ),
      .cfg_en360           (cfg_en360              ),
      .cfg_en361           (cfg_en361              ),
      .cfg_en362           (cfg_en362              ),
      .cfg_en363           (cfg_en363              ),
      .cfg_en364           (cfg_en364              ),
      .cfg_en365           (cfg_en365              ),
      .cfg_en366           (cfg_en366              ),
      .cfg_en367           (cfg_en367              ),
      .cfg_en368           (cfg_en368              ),
      .cfg_en369           (cfg_en369              ),
      .cfg_en370           (cfg_en370              ),
      .cfg_en371           (cfg_en371              ),
      .cfg_en372           (cfg_en372              ),
      .cfg_en373           (cfg_en373              ),
      .cfg_en374           (cfg_en374              ),
      .cfg_en375           (cfg_en375              ),
      .cfg_en376           (cfg_en376              ),
      .cfg_en377           (cfg_en377              ),
      .cfg_en378           (cfg_en378              ),
      .cfg_en379           (cfg_en379              ),
      .cfg_en380           (cfg_en380              ),
      .cfg_en381           (cfg_en381              ),
      .cfg_en382           (cfg_en382              ),
      .cfg_en383           (cfg_en383              ),
      .cfg_en384           (cfg_en384              ),
      .cfg_en385           (cfg_en385              ),
      .cfg_en386           (cfg_en386              ),
      .cfg_en387           (cfg_en387              ),
      .cfg_en388           (cfg_en388              ),
      .cfg_en389           (cfg_en389              ),
      .cfg_en390           (cfg_en390              ),
      .cfg_en391           (cfg_en391              ),
      .cfg_en392           (cfg_en392              ),
      .cfg_en393           (cfg_en393              ),
      .cfg_en394           (cfg_en394              ),
      .cfg_en395           (cfg_en395              ),
      .cfg_en396           (cfg_en396              ),
      .cfg_en397           (cfg_en397              ),
      .cfg_en398           (cfg_en398              ),
      .cfg_en399           (cfg_en399              ),
      .cfg_en400           (cfg_en400              ),
      .cfg_en401           (cfg_en401              ),
      .cfg_en402           (cfg_en402              ),
      .cfg_en403           (cfg_en403              ),
      .cfg_en404           (cfg_en404              ),
      .cfg_en405           (cfg_en405              ),
      .cfg_en406           (cfg_en406              ),
      .cfg_en407           (cfg_en407              ),
      .cfg_en408           (cfg_en408              ),
      .cfg_en409           (cfg_en409              ),
      .cfg_en410           (cfg_en410              ),
      .cfg_en411           (cfg_en411              ),
      .cfg_en412           (cfg_en412              ),
      .cfg_en413           (cfg_en413              ),
      .cfg_en414           (cfg_en414              ),
      .cfg_en415           (cfg_en415              ),
      .cfg_en416           (cfg_en416              ),
      .cfg_en417           (cfg_en417              ),
      .cfg_en418           (cfg_en418              ),
      .cfg_en419           (cfg_en419              ),
      .cfg_en420           (cfg_en420              ),
      .cfg_en421           (cfg_en421              ),
      .cfg_en422           (cfg_en422              ),
      .cfg_en423           (cfg_en423              ),
      .cfg_en424           (cfg_en424              ),
      .cfg_en425           (cfg_en425              ),
      .cfg_en426           (cfg_en426              ),
      .cfg_en427           (cfg_en427              ),
      .cfg_en428           (cfg_en428              ),
      .cfg_en429           (cfg_en429              ),
      .cfg_en430           (cfg_en430              ),
      .cfg_en431           (cfg_en431              ),
      .cfg_en432           (cfg_en432              ),
      .cfg_en433           (cfg_en433              ),
      .cfg_en434           (cfg_en434              ),
      .cfg_en435           (cfg_en435              ),
      .cfg_en436           (cfg_en436              ),
      .cfg_en437           (cfg_en437              ),
      .cfg_en438           (cfg_en438              ),
      .cfg_en439           (cfg_en439              ),
      .cfg_en440           (cfg_en440              ),
      .cfg_en441           (cfg_en441              ),
      .cfg_en442           (cfg_en442              ),
      .cfg_en443           (cfg_en443              ),
      .cfg_en444           (cfg_en444              ),
      .cfg_en445           (cfg_en445              ),
      .cfg_en446           (cfg_en446              ),
      .cfg_en447           (cfg_en447              ),
      .cfg_en448           (cfg_en448              ),
      .cfg_en449           (cfg_en449              ),
      .cfg_en450           (cfg_en450              ),
      .cfg_en451           (cfg_en451              ),
      .cfg_en452           (cfg_en452              ),
      .cfg_en453           (cfg_en453              ),
      .cfg_en454           (cfg_en454              ),
      .cfg_en455           (cfg_en455              ),
      .cfg_en456           (cfg_en456              ),
      .cfg_en457           (cfg_en457              ),
      .cfg_en458           (cfg_en458              ),
      .cfg_en459           (cfg_en459              ),
      .cfg_en460           (cfg_en460              ),
      .cfg_en461           (cfg_en461              ),
      .cfg_en462           (cfg_en462              ),
      .cfg_en463           (cfg_en463              ),
      .cfg_en464           (cfg_en464              ),
      .cfg_en465           (cfg_en465              ),
      .cfg_en466           (cfg_en466              ),
      .cfg_en467           (cfg_en467              ),
      .cfg_en468           (cfg_en468              ),
      .cfg_en469           (cfg_en469              ),
      .cfg_en470           (cfg_en470              ),
      .cfg_en471           (cfg_en471              ),
      .cfg_en472           (cfg_en472              ),
      .cfg_en473           (cfg_en473              ),
      .cfg_en474           (cfg_en474              ),
      .cfg_en475           (cfg_en475              ),
      .cfg_en476           (cfg_en476              ),
      .cfg_en477           (cfg_en477              ),
      .cfg_en478           (cfg_en478              ),
      .cfg_en479           (cfg_en479              ),
      .cfg_en480           (cfg_en480              ),
      .cfg_en481           (cfg_en481              ),
      .cfg_en482           (cfg_en482              ),
      .cfg_en483           (cfg_en483              ),
      .cfg_en484           (cfg_en484              ),
      .cfg_en485           (cfg_en485              ),
      .cfg_en486           (cfg_en486              ),
      .cfg_en487           (cfg_en487              ),
      .cfg_en488           (cfg_en488              ),
      .cfg_en489           (cfg_en489              ),
      .cfg_en490           (cfg_en490              ),
      .cfg_en491           (cfg_en491              ),
      .cfg_en492           (cfg_en492              ),
      .cfg_en493           (cfg_en493              ),
      .cfg_en494           (cfg_en494              ),
      .cfg_en495           (cfg_en495              ),
      .cfg_en496           (cfg_en496              ),
      .cfg_en497           (cfg_en497              ),
      .cfg_en498           (cfg_en498              ),
      .cfg_en499           (cfg_en499              ),
      .cfg_en500           (cfg_en500              ),
      .cfg_en501           (cfg_en501              ),
      .cfg_en502           (cfg_en502              ),
      .cfg_en503           (cfg_en503              ),
      .cfg_en504           (cfg_en504              ),
      .cfg_en505           (cfg_en505              ),
      .cfg_en506           (cfg_en506              ),
      .cfg_en507           (cfg_en507              ),
      .cfg_en508           (cfg_en508              ),
      .cfg_en509           (cfg_en509              ),
      .cfg_en510           (cfg_en510              ),
      .cfg_en511           (cfg_en511              ),
      .match_out0        (match_out0           ),
      .match_out1        (match_out1           ),
      .match_out2        (match_out2           ),
      .match_out3        (match_out3           ),
      .match_out4        (match_out4           ),
      .match_out5        (match_out5           ),
      .match_out6        (match_out6           ),
      .match_out7        (match_out7           ),
      .match_out8        (match_out8           ),
      .match_out9        (match_out9           ),
      .match_out10        (match_out10           ),
      .match_out11        (match_out11           ),
      .match_out12        (match_out12           ),
      .match_out13        (match_out13           ),
      .match_out14        (match_out14           ),
      .match_out15        (match_out15           ),
      .match_out16        (match_out16           ),
      .match_out17        (match_out17           ),
      .match_out18        (match_out18           ),
      .match_out19        (match_out19           ),
      .match_out20        (match_out20           ),
      .match_out21        (match_out21           ),
      .match_out22        (match_out22           ),
      .match_out23        (match_out23           ),
      .match_out24        (match_out24           ),
      .match_out25        (match_out25           ),
      .match_out26        (match_out26           ),
      .match_out27        (match_out27           ),
      .match_out28        (match_out28           ),
      .match_out29        (match_out29           ),
      .match_out30        (match_out30           ),
      .match_out31        (match_out31           ),
      .match_out32        (match_out32           ),
      .match_out33        (match_out33           ),
      .match_out34        (match_out34           ),
      .match_out35        (match_out35           ),
      .match_out36        (match_out36           ),
      .match_out37        (match_out37           ),
      .match_out38        (match_out38           ),
      .match_out39        (match_out39           ),
      .match_out40        (match_out40           ),
      .match_out41        (match_out41           ),
      .match_out42        (match_out42           ),
      .match_out43        (match_out43           ),
      .match_out44        (match_out44           ),
      .match_out45        (match_out45           ),
      .match_out46        (match_out46           ),
      .match_out47        (match_out47           ),
      .match_out48        (match_out48           ),
      .match_out49        (match_out49           ),
      .match_out50        (match_out50           ),
      .match_out51        (match_out51           ),
      .match_out52        (match_out52           ),
      .match_out53        (match_out53           ),
      .match_out54        (match_out54           ),
      .match_out55        (match_out55           ),
      .match_out56        (match_out56           ),
      .match_out57        (match_out57           ),
      .match_out58        (match_out58           ),
      .match_out59        (match_out59           ),
      .match_out60        (match_out60           ),
      .match_out61        (match_out61           ),
      .match_out62        (match_out62           ),
      .match_out63        (match_out63           ),
      .match_out64        (match_out64           ),
      .match_out65        (match_out65           ),
      .match_out66        (match_out66           ),
      .match_out67        (match_out67           ),
      .match_out68        (match_out68           ),
      .match_out69        (match_out69           ),
      .match_out70        (match_out70           ),
      .match_out71        (match_out71           ),
      .match_out72        (match_out72           ),
      .match_out73        (match_out73           ),
      .match_out74        (match_out74           ),
      .match_out75        (match_out75           ),
      .match_out76        (match_out76           ),
      .match_out77        (match_out77           ),
      .match_out78        (match_out78           ),
      .match_out79        (match_out79           ),
      .match_out80        (match_out80           ),
      .match_out81        (match_out81           ),
      .match_out82        (match_out82           ),
      .match_out83        (match_out83           ),
      .match_out84        (match_out84           ),
      .match_out85        (match_out85           ),
      .match_out86        (match_out86           ),
      .match_out87        (match_out87           ),
      .match_out88        (match_out88           ),
      .match_out89        (match_out89           ),
      .match_out90        (match_out90           ),
      .match_out91        (match_out91           ),
      .match_out92        (match_out92           ),
      .match_out93        (match_out93           ),
      .match_out94        (match_out94           ),
      .match_out95        (match_out95           ),
      .match_out96        (match_out96           ),
      .match_out97        (match_out97           ),
      .match_out98        (match_out98           ),
      .match_out99        (match_out99           ),
      .match_out100        (match_out100           ),
      .match_out101        (match_out101           ),
      .match_out102        (match_out102           ),
      .match_out103        (match_out103           ),
      .match_out104        (match_out104           ),
      .match_out105        (match_out105           ),
      .match_out106        (match_out106           ),
      .match_out107        (match_out107           ),
      .match_out108        (match_out108           ),
      .match_out109        (match_out109           ),
      .match_out110        (match_out110           ),
      .match_out111        (match_out111           ),
      .match_out112        (match_out112           ),
      .match_out113        (match_out113           ),
      .match_out114        (match_out114           ),
      .match_out115        (match_out115           ),
      .match_out116        (match_out116           ),
      .match_out117        (match_out117           ),
      .match_out118        (match_out118           ),
      .match_out119        (match_out119           ),
      .match_out120        (match_out120           ),
      .match_out121        (match_out121           ),
      .match_out122        (match_out122           ),
      .match_out123        (match_out123           ),
      .match_out124        (match_out124           ),
      .match_out125        (match_out125           ),
      .match_out126        (match_out126           ),
      .match_out127        (match_out127           ),
      .match_out128        (match_out128           ),
      .match_out129        (match_out129           ),
      .match_out130        (match_out130           ),
      .match_out131        (match_out131           ),
      .match_out132        (match_out132           ),
      .match_out133        (match_out133           ),
      .match_out134        (match_out134           ),
      .match_out135        (match_out135           ),
      .match_out136        (match_out136           ),
      .match_out137        (match_out137           ),
      .match_out138        (match_out138           ),
      .match_out139        (match_out139           ),
      .match_out140        (match_out140           ),
      .match_out141        (match_out141           ),
      .match_out142        (match_out142           ),
      .match_out143        (match_out143           ),
      .match_out144        (match_out144           ),
      .match_out145        (match_out145           ),
      .match_out146        (match_out146           ),
      .match_out147        (match_out147           ),
      .match_out148        (match_out148           ),
      .match_out149        (match_out149           ),
      .match_out150        (match_out150           ),
      .match_out151        (match_out151           ),
      .match_out152        (match_out152           ),
      .match_out153        (match_out153           ),
      .match_out154        (match_out154           ),
      .match_out155        (match_out155           ),
      .match_out156        (match_out156           ),
      .match_out157        (match_out157           ),
      .match_out158        (match_out158           ),
      .match_out159        (match_out159           ),
      .match_out160        (match_out160           ),
      .match_out161        (match_out161           ),
      .match_out162        (match_out162           ),
      .match_out163        (match_out163           ),
      .match_out164        (match_out164           ),
      .match_out165        (match_out165           ),
      .match_out166        (match_out166           ),
      .match_out167        (match_out167           ),
      .match_out168        (match_out168           ),
      .match_out169        (match_out169           ),
      .match_out170        (match_out170           ),
      .match_out171        (match_out171           ),
      .match_out172        (match_out172           ),
      .match_out173        (match_out173           ),
      .match_out174        (match_out174           ),
      .match_out175        (match_out175           ),
      .match_out176        (match_out176           ),
      .match_out177        (match_out177           ),
      .match_out178        (match_out178           ),
      .match_out179        (match_out179           ),
      .match_out180        (match_out180           ),
      .match_out181        (match_out181           ),
      .match_out182        (match_out182           ),
      .match_out183        (match_out183           ),
      .match_out184        (match_out184           ),
      .match_out185        (match_out185           ),
      .match_out186        (match_out186           ),
      .match_out187        (match_out187           ),
      .match_out188        (match_out188           ),
      .match_out189        (match_out189           ),
      .match_out190        (match_out190           ),
      .match_out191        (match_out191           ),
      .match_out192        (match_out192           ),
      .match_out193        (match_out193           ),
      .match_out194        (match_out194           ),
      .match_out195        (match_out195           ),
      .match_out196        (match_out196           ),
      .match_out197        (match_out197           ),
      .match_out198        (match_out198           ),
      .match_out199        (match_out199           ),
      .match_out200        (match_out200           ),
      .match_out201        (match_out201           ),
      .match_out202        (match_out202           ),
      .match_out203        (match_out203           ),
      .match_out204        (match_out204           ),
      .match_out205        (match_out205           ),
      .match_out206        (match_out206           ),
      .match_out207        (match_out207           ),
      .match_out208        (match_out208           ),
      .match_out209        (match_out209           ),
      .match_out210        (match_out210           ),
      .match_out211        (match_out211           ),
      .match_out212        (match_out212           ),
      .match_out213        (match_out213           ),
      .match_out214        (match_out214           ),
      .match_out215        (match_out215           ),
      .match_out216        (match_out216           ),
      .match_out217        (match_out217           ),
      .match_out218        (match_out218           ),
      .match_out219        (match_out219           ),
      .match_out220        (match_out220           ),
      .match_out221        (match_out221           ),
      .match_out222        (match_out222           ),
      .match_out223        (match_out223           ),
      .match_out224        (match_out224           ),
      .match_out225        (match_out225           ),
      .match_out226        (match_out226           ),
      .match_out227        (match_out227           ),
      .match_out228        (match_out228           ),
      .match_out229        (match_out229           ),
      .match_out230        (match_out230           ),
      .match_out231        (match_out231           ),
      .match_out232        (match_out232           ),
      .match_out233        (match_out233           ),
      .match_out234        (match_out234           ),
      .match_out235        (match_out235           ),
      .match_out236        (match_out236           ),
      .match_out237        (match_out237           ),
      .match_out238        (match_out238           ),
      .match_out239        (match_out239           ),
      .match_out240        (match_out240           ),
      .match_out241        (match_out241           ),
      .match_out242        (match_out242           ),
      .match_out243        (match_out243           ),
      .match_out244        (match_out244           ),
      .match_out245        (match_out245           ),
      .match_out246        (match_out246           ),
      .match_out247        (match_out247           ),
      .match_out248        (match_out248           ),
      .match_out249        (match_out249           ),
      .match_out250        (match_out250           ),
      .match_out251        (match_out251           ),
      .match_out252        (match_out252           ),
      .match_out253        (match_out253           ),
      .match_out254        (match_out254           ),
      .match_out255        (match_out255           ),
      .match_out256        (match_out256           ),
      .match_out257        (match_out257           ),
      .match_out258        (match_out258           ),
      .match_out259        (match_out259           ),
      .match_out260        (match_out260           ),
      .match_out261        (match_out261           ),
      .match_out262        (match_out262           ),
      .match_out263        (match_out263           ),
      .match_out264        (match_out264           ),
      .match_out265        (match_out265           ),
      .match_out266        (match_out266           ),
      .match_out267        (match_out267           ),
      .match_out268        (match_out268           ),
      .match_out269        (match_out269           ),
      .match_out270        (match_out270           ),
      .match_out271        (match_out271           ),
      .match_out272        (match_out272           ),
      .match_out273        (match_out273           ),
      .match_out274        (match_out274           ),
      .match_out275        (match_out275           ),
      .match_out276        (match_out276           ),
      .match_out277        (match_out277           ),
      .match_out278        (match_out278           ),
      .match_out279        (match_out279           ),
      .match_out280        (match_out280           ),
      .match_out281        (match_out281           ),
      .match_out282        (match_out282           ),
      .match_out283        (match_out283           ),
      .match_out284        (match_out284           ),
      .match_out285        (match_out285           ),
      .match_out286        (match_out286           ),
      .match_out287        (match_out287           ),
      .match_out288        (match_out288           ),
      .match_out289        (match_out289           ),
      .match_out290        (match_out290           ),
      .match_out291        (match_out291           ),
      .match_out292        (match_out292           ),
      .match_out293        (match_out293           ),
      .match_out294        (match_out294           ),
      .match_out295        (match_out295           ),
      .match_out296        (match_out296           ),
      .match_out297        (match_out297           ),
      .match_out298        (match_out298           ),
      .match_out299        (match_out299           ),
      .match_out300        (match_out300           ),
      .match_out301        (match_out301           ),
      .match_out302        (match_out302           ),
      .match_out303        (match_out303           ),
      .match_out304        (match_out304           ),
      .match_out305        (match_out305           ),
      .match_out306        (match_out306           ),
      .match_out307        (match_out307           ),
      .match_out308        (match_out308           ),
      .match_out309        (match_out309           ),
      .match_out310        (match_out310           ),
      .match_out311        (match_out311           ),
      .match_out312        (match_out312           ),
      .match_out313        (match_out313           ),
      .match_out314        (match_out314           ),
      .match_out315        (match_out315           ),
      .match_out316        (match_out316           ),
      .match_out317        (match_out317           ),
      .match_out318        (match_out318           ),
      .match_out319        (match_out319           ),
      .match_out320        (match_out320           ),
      .match_out321        (match_out321           ),
      .match_out322        (match_out322           ),
      .match_out323        (match_out323           ),
      .match_out324        (match_out324           ),
      .match_out325        (match_out325           ),
      .match_out326        (match_out326           ),
      .match_out327        (match_out327           ),
      .match_out328        (match_out328           ),
      .match_out329        (match_out329           ),
      .match_out330        (match_out330           ),
      .match_out331        (match_out331           ),
      .match_out332        (match_out332           ),
      .match_out333        (match_out333           ),
      .match_out334        (match_out334           ),
      .match_out335        (match_out335           ),
      .match_out336        (match_out336           ),
      .match_out337        (match_out337           ),
      .match_out338        (match_out338           ),
      .match_out339        (match_out339           ),
      .match_out340        (match_out340           ),
      .match_out341        (match_out341           ),
      .match_out342        (match_out342           ),
      .match_out343        (match_out343           ),
      .match_out344        (match_out344           ),
      .match_out345        (match_out345           ),
      .match_out346        (match_out346           ),
      .match_out347        (match_out347           ),
      .match_out348        (match_out348           ),
      .match_out349        (match_out349           ),
      .match_out350        (match_out350           ),
      .match_out351        (match_out351           ),
      .match_out352        (match_out352           ),
      .match_out353        (match_out353           ),
      .match_out354        (match_out354           ),
      .match_out355        (match_out355           ),
      .match_out356        (match_out356           ),
      .match_out357        (match_out357           ),
      .match_out358        (match_out358           ),
      .match_out359        (match_out359           ),
      .match_out360        (match_out360           ),
      .match_out361        (match_out361           ),
      .match_out362        (match_out362           ),
      .match_out363        (match_out363           ),
      .match_out364        (match_out364           ),
      .match_out365        (match_out365           ),
      .match_out366        (match_out366           ),
      .match_out367        (match_out367           ),
      .match_out368        (match_out368           ),
      .match_out369        (match_out369           ),
      .match_out370        (match_out370           ),
      .match_out371        (match_out371           ),
      .match_out372        (match_out372           ),
      .match_out373        (match_out373           ),
      .match_out374        (match_out374           ),
      .match_out375        (match_out375           ),
      .match_out376        (match_out376           ),
      .match_out377        (match_out377           ),
      .match_out378        (match_out378           ),
      .match_out379        (match_out379           ),
      .match_out380        (match_out380           ),
      .match_out381        (match_out381           ),
      .match_out382        (match_out382           ),
      .match_out383        (match_out383           ),
      .match_out384        (match_out384           ),
      .match_out385        (match_out385           ),
      .match_out386        (match_out386           ),
      .match_out387        (match_out387           ),
      .match_out388        (match_out388           ),
      .match_out389        (match_out389           ),
      .match_out390        (match_out390           ),
      .match_out391        (match_out391           ),
      .match_out392        (match_out392           ),
      .match_out393        (match_out393           ),
      .match_out394        (match_out394           ),
      .match_out395        (match_out395           ),
      .match_out396        (match_out396           ),
      .match_out397        (match_out397           ),
      .match_out398        (match_out398           ),
      .match_out399        (match_out399           ),
      .match_out400        (match_out400           ),
      .match_out401        (match_out401           ),
      .match_out402        (match_out402           ),
      .match_out403        (match_out403           ),
      .match_out404        (match_out404           ),
      .match_out405        (match_out405           ),
      .match_out406        (match_out406           ),
      .match_out407        (match_out407           ),
      .match_out408        (match_out408           ),
      .match_out409        (match_out409           ),
      .match_out410        (match_out410           ),
      .match_out411        (match_out411           ),
      .match_out412        (match_out412           ),
      .match_out413        (match_out413           ),
      .match_out414        (match_out414           ),
      .match_out415        (match_out415           ),
      .match_out416        (match_out416           ),
      .match_out417        (match_out417           ),
      .match_out418        (match_out418           ),
      .match_out419        (match_out419           ),
      .match_out420        (match_out420           ),
      .match_out421        (match_out421           ),
      .match_out422        (match_out422           ),
      .match_out423        (match_out423           ),
      .match_out424        (match_out424           ),
      .match_out425        (match_out425           ),
      .match_out426        (match_out426           ),
      .match_out427        (match_out427           ),
      .match_out428        (match_out428           ),
      .match_out429        (match_out429           ),
      .match_out430        (match_out430           ),
      .match_out431        (match_out431           ),
      .match_out432        (match_out432           ),
      .match_out433        (match_out433           ),
      .match_out434        (match_out434           ),
      .match_out435        (match_out435           ),
      .match_out436        (match_out436           ),
      .match_out437        (match_out437           ),
      .match_out438        (match_out438           ),
      .match_out439        (match_out439           ),
      .match_out440        (match_out440           ),
      .match_out441        (match_out441           ),
      .match_out442        (match_out442           ),
      .match_out443        (match_out443           ),
      .match_out444        (match_out444           ),
      .match_out445        (match_out445           ),
      .match_out446        (match_out446           ),
      .match_out447        (match_out447           ),
      .match_out448        (match_out448           ),
      .match_out449        (match_out449           ),
      .match_out450        (match_out450           ),
      .match_out451        (match_out451           ),
      .match_out452        (match_out452           ),
      .match_out453        (match_out453           ),
      .match_out454        (match_out454           ),
      .match_out455        (match_out455           ),
      .match_out456        (match_out456           ),
      .match_out457        (match_out457           ),
      .match_out458        (match_out458           ),
      .match_out459        (match_out459           ),
      .match_out460        (match_out460           ),
      .match_out461        (match_out461           ),
      .match_out462        (match_out462           ),
      .match_out463        (match_out463           ),
      .match_out464        (match_out464           ),
      .match_out465        (match_out465           ),
      .match_out466        (match_out466           ),
      .match_out467        (match_out467           ),
      .match_out468        (match_out468           ),
      .match_out469        (match_out469           ),
      .match_out470        (match_out470           ),
      .match_out471        (match_out471           ),
      .match_out472        (match_out472           ),
      .match_out473        (match_out473           ),
      .match_out474        (match_out474           ),
      .match_out475        (match_out475           ),
      .match_out476        (match_out476           ),
      .match_out477        (match_out477           ),
      .match_out478        (match_out478           ),
      .match_out479        (match_out479           ),
      .match_out480        (match_out480           ),
      .match_out481        (match_out481           ),
      .match_out482        (match_out482           ),
      .match_out483        (match_out483           ),
      .match_out484        (match_out484           ),
      .match_out485        (match_out485           ),
      .match_out486        (match_out486           ),
      .match_out487        (match_out487           ),
      .match_out488        (match_out488           ),
      .match_out489        (match_out489           ),
      .match_out490        (match_out490           ),
      .match_out491        (match_out491           ),
      .match_out492        (match_out492           ),
      .match_out493        (match_out493           ),
      .match_out494        (match_out494           ),
      .match_out495        (match_out495           ),
      .match_out496        (match_out496           ),
      .match_out497        (match_out497           ),
      .match_out498        (match_out498           ),
      .match_out499        (match_out499           ),
      .match_out500        (match_out500           ),
      .match_out501        (match_out501           ),
      .match_out502        (match_out502           ),
      .match_out503        (match_out503           ),
      .match_out504        (match_out504           ),
      .match_out505        (match_out505           ),
      .match_out506        (match_out506           ),
      .match_out507        (match_out507           ),
      .match_out508        (match_out508           ),
      .match_out509        (match_out509           ),
      .match_out510        (match_out510           ),
      .match_out511        (match_out511           ),
      .match_out              (trigger_din               )
     );


