      input  [C_PROBE0_WIDTH-1:0]             probe0,
      input  [C_PROBE1_WIDTH-1:0]             probe1,
      input  [C_PROBE2_WIDTH-1:0]             probe2,
      input  [C_PROBE3_WIDTH-1:0]             probe3,
      input  [C_PROBE4_WIDTH-1:0]             probe4,
      input  [C_PROBE5_WIDTH-1:0]             probe5,
      input  [C_PROBE6_WIDTH-1:0]             probe6,
      input  [C_PROBE7_WIDTH-1:0]             probe7,
      input  [C_PROBE8_WIDTH-1:0]             probe8,
      input  [C_PROBE9_WIDTH-1:0]             probe9,
      input  [C_PROBE10_WIDTH-1:0]            probe10,
      input  [C_PROBE11_WIDTH-1:0]            probe11,
      input  [C_PROBE12_WIDTH-1:0]            probe12,
      input  [C_PROBE13_WIDTH-1:0]            probe13,
      input  [C_PROBE14_WIDTH-1:0]            probe14,
      input  [C_PROBE15_WIDTH-1:0]            probe15,
      input  [C_PROBE16_WIDTH-1:0]            probe16,
      input  [C_PROBE17_WIDTH-1:0]            probe17,
      input  [C_PROBE18_WIDTH-1:0]            probe18,
      input  [C_PROBE19_WIDTH-1:0]            probe19,
      input  [C_PROBE20_WIDTH-1:0]            probe20,
      input  [C_PROBE21_WIDTH-1:0]            probe21,
      input  [C_PROBE22_WIDTH-1:0]            probe22,
      input  [C_PROBE23_WIDTH-1:0]            probe23,
      input  [C_PROBE24_WIDTH-1:0]            probe24,
      input  [C_PROBE25_WIDTH-1:0]            probe25,
      input  [C_PROBE26_WIDTH-1:0]            probe26,
      input  [C_PROBE27_WIDTH-1:0]            probe27,
      input  [C_PROBE28_WIDTH-1:0]            probe28,
      input  [C_PROBE29_WIDTH-1:0]            probe29,
      input  [C_PROBE30_WIDTH-1:0]            probe30,
      input  [C_PROBE31_WIDTH-1:0]            probe31,
      input  [C_PROBE32_WIDTH-1:0]            probe32,
      input  [C_PROBE33_WIDTH-1:0]            probe33,
      input  [C_PROBE34_WIDTH-1:0]            probe34,
      input  [C_PROBE35_WIDTH-1:0]            probe35,
      input  [C_PROBE36_WIDTH-1:0]            probe36,
      input  [C_PROBE37_WIDTH-1:0]            probe37,
      input  [C_PROBE38_WIDTH-1:0]            probe38,
      input  [C_PROBE39_WIDTH-1:0]            probe39,
      input  [C_PROBE40_WIDTH-1:0]            probe40,
      input  [C_PROBE41_WIDTH-1:0]            probe41,
      input  [C_PROBE42_WIDTH-1:0]            probe42,
      input  [C_PROBE43_WIDTH-1:0]            probe43,
      input  [C_PROBE44_WIDTH-1:0]            probe44,
      input  [C_PROBE45_WIDTH-1:0]            probe45,
      input  [C_PROBE46_WIDTH-1:0]            probe46,
      input  [C_PROBE47_WIDTH-1:0]            probe47,
      input  [C_PROBE48_WIDTH-1:0]            probe48,
      input  [C_PROBE49_WIDTH-1:0]            probe49,
      input  [C_PROBE50_WIDTH-1:0]            probe50,
      input  [C_PROBE51_WIDTH-1:0]            probe51,
      input  [C_PROBE52_WIDTH-1:0]            probe52,
      input  [C_PROBE53_WIDTH-1:0]            probe53,
      input  [C_PROBE54_WIDTH-1:0]            probe54,
      input  [C_PROBE55_WIDTH-1:0]            probe55,
      input  [C_PROBE56_WIDTH-1:0]            probe56,
      input  [C_PROBE57_WIDTH-1:0]            probe57,
      input  [C_PROBE58_WIDTH-1:0]            probe58,
      input  [C_PROBE59_WIDTH-1:0]            probe59,
      input  [C_PROBE60_WIDTH-1:0]            probe60,
      input  [C_PROBE61_WIDTH-1:0]            probe61,
      input  [C_PROBE62_WIDTH-1:0]            probe62,
      input  [C_PROBE63_WIDTH-1:0]            probe63,
      input  [C_PROBE64_WIDTH-1:0]            probe64,
      input  [C_PROBE65_WIDTH-1:0]            probe65,
      input  [C_PROBE66_WIDTH-1:0]            probe66,
      input  [C_PROBE67_WIDTH-1:0]            probe67,
      input  [C_PROBE68_WIDTH-1:0]            probe68,
      input  [C_PROBE69_WIDTH-1:0]            probe69,
      input  [C_PROBE70_WIDTH-1:0]            probe70,
      input  [C_PROBE71_WIDTH-1:0]            probe71,
      input  [C_PROBE72_WIDTH-1:0]            probe72,
      input  [C_PROBE73_WIDTH-1:0]            probe73,
      input  [C_PROBE74_WIDTH-1:0]            probe74,
      input  [C_PROBE75_WIDTH-1:0]            probe75,
      input  [C_PROBE76_WIDTH-1:0]            probe76,
      input  [C_PROBE77_WIDTH-1:0]            probe77,
      input  [C_PROBE78_WIDTH-1:0]            probe78,
      input  [C_PROBE79_WIDTH-1:0]            probe79,
      input  [C_PROBE80_WIDTH-1:0]            probe80,
      input  [C_PROBE81_WIDTH-1:0]            probe81,
      input  [C_PROBE82_WIDTH-1:0]            probe82,
      input  [C_PROBE83_WIDTH-1:0]            probe83,
      input  [C_PROBE84_WIDTH-1:0]            probe84,
      input  [C_PROBE85_WIDTH-1:0]            probe85,
      input  [C_PROBE86_WIDTH-1:0]            probe86,
      input  [C_PROBE87_WIDTH-1:0]            probe87,
      input  [C_PROBE88_WIDTH-1:0]            probe88,
      input  [C_PROBE89_WIDTH-1:0]            probe89,
      input  [C_PROBE90_WIDTH-1:0]            probe90,
      input  [C_PROBE91_WIDTH-1:0]            probe91,
      input  [C_PROBE92_WIDTH-1:0]            probe92,
      input  [C_PROBE93_WIDTH-1:0]            probe93,
      input  [C_PROBE94_WIDTH-1:0]            probe94,
      input  [C_PROBE95_WIDTH-1:0]            probe95,
      input  [C_PROBE96_WIDTH-1:0]            probe96,
      input  [C_PROBE97_WIDTH-1:0]            probe97,
      input  [C_PROBE98_WIDTH-1:0]            probe98,
      input  [C_PROBE99_WIDTH-1:0]            probe99,
      input  [C_PROBE100_WIDTH-1:0]           probe100,
      input  [C_PROBE101_WIDTH-1:0]           probe101,
      input  [C_PROBE102_WIDTH-1:0]           probe102,
      input  [C_PROBE103_WIDTH-1:0]           probe103,
      input  [C_PROBE104_WIDTH-1:0]           probe104,
      input  [C_PROBE105_WIDTH-1:0]           probe105,
      input  [C_PROBE106_WIDTH-1:0]           probe106,
      input  [C_PROBE107_WIDTH-1:0]           probe107,
      input  [C_PROBE108_WIDTH-1:0]           probe108,
      input  [C_PROBE109_WIDTH-1:0]           probe109,
      input  [C_PROBE110_WIDTH-1:0]           probe110,
      input  [C_PROBE111_WIDTH-1:0]           probe111,
      input  [C_PROBE112_WIDTH-1:0]           probe112,
      input  [C_PROBE113_WIDTH-1:0]           probe113,
      input  [C_PROBE114_WIDTH-1:0]           probe114,
      input  [C_PROBE115_WIDTH-1:0]           probe115,
      input  [C_PROBE116_WIDTH-1:0]           probe116,
      input  [C_PROBE117_WIDTH-1:0]           probe117,
      input  [C_PROBE118_WIDTH-1:0]           probe118,
      input  [C_PROBE119_WIDTH-1:0]           probe119,
      input  [C_PROBE120_WIDTH-1:0]           probe120,
      input  [C_PROBE121_WIDTH-1:0]           probe121,
      input  [C_PROBE122_WIDTH-1:0]           probe122,
      input  [C_PROBE123_WIDTH-1:0]           probe123,
      input  [C_PROBE124_WIDTH-1:0]           probe124,
      input  [C_PROBE125_WIDTH-1:0]           probe125,
      input  [C_PROBE126_WIDTH-1:0]           probe126,
      input  [C_PROBE127_WIDTH-1:0]           probe127,
      input  [C_PROBE128_WIDTH-1:0]           probe128,
      input  [C_PROBE129_WIDTH-1:0]           probe129,
      input  [C_PROBE130_WIDTH-1:0]           probe130,
      input  [C_PROBE131_WIDTH-1:0]           probe131,
      input  [C_PROBE132_WIDTH-1:0]           probe132,
      input  [C_PROBE133_WIDTH-1:0]           probe133,
      input  [C_PROBE134_WIDTH-1:0]           probe134,
      input  [C_PROBE135_WIDTH-1:0]           probe135,
      input  [C_PROBE136_WIDTH-1:0]           probe136,
      input  [C_PROBE137_WIDTH-1:0]           probe137,
      input  [C_PROBE138_WIDTH-1:0]           probe138,
      input  [C_PROBE139_WIDTH-1:0]           probe139,
      input  [C_PROBE140_WIDTH-1:0]           probe140,
      input  [C_PROBE141_WIDTH-1:0]           probe141,
      input  [C_PROBE142_WIDTH-1:0]           probe142,
      input  [C_PROBE143_WIDTH-1:0]           probe143,
      input  [C_PROBE144_WIDTH-1:0]           probe144,
      input  [C_PROBE145_WIDTH-1:0]           probe145,
      input  [C_PROBE146_WIDTH-1:0]           probe146,
      input  [C_PROBE147_WIDTH-1:0]           probe147,
      input  [C_PROBE148_WIDTH-1:0]           probe148,
      input  [C_PROBE149_WIDTH-1:0]           probe149,
      input  [C_PROBE150_WIDTH-1:0]           probe150,
      input  [C_PROBE151_WIDTH-1:0]           probe151,
      input  [C_PROBE152_WIDTH-1:0]           probe152,
      input  [C_PROBE153_WIDTH-1:0]           probe153,
      input  [C_PROBE154_WIDTH-1:0]           probe154,
      input  [C_PROBE155_WIDTH-1:0]           probe155,
      input  [C_PROBE156_WIDTH-1:0]           probe156,
      input  [C_PROBE157_WIDTH-1:0]           probe157,
      input  [C_PROBE158_WIDTH-1:0]           probe158,
      input  [C_PROBE159_WIDTH-1:0]           probe159,
      input  [C_PROBE160_WIDTH-1:0]           probe160,
      input  [C_PROBE161_WIDTH-1:0]           probe161,
      input  [C_PROBE162_WIDTH-1:0]           probe162,
      input  [C_PROBE163_WIDTH-1:0]           probe163,
      input  [C_PROBE164_WIDTH-1:0]           probe164,
      input  [C_PROBE165_WIDTH-1:0]           probe165,
      input  [C_PROBE166_WIDTH-1:0]           probe166,
      input  [C_PROBE167_WIDTH-1:0]           probe167,
      input  [C_PROBE168_WIDTH-1:0]           probe168,
      input  [C_PROBE169_WIDTH-1:0]           probe169,
      input  [C_PROBE170_WIDTH-1:0]           probe170,
      input  [C_PROBE171_WIDTH-1:0]           probe171,
      input  [C_PROBE172_WIDTH-1:0]           probe172,
      input  [C_PROBE173_WIDTH-1:0]           probe173,
      input  [C_PROBE174_WIDTH-1:0]           probe174,
      input  [C_PROBE175_WIDTH-1:0]           probe175,
      input  [C_PROBE176_WIDTH-1:0]           probe176,
      input  [C_PROBE177_WIDTH-1:0]           probe177,
      input  [C_PROBE178_WIDTH-1:0]           probe178,
      input  [C_PROBE179_WIDTH-1:0]           probe179,
      input  [C_PROBE180_WIDTH-1:0]           probe180,
      input  [C_PROBE181_WIDTH-1:0]           probe181,
      input  [C_PROBE182_WIDTH-1:0]           probe182,
      input  [C_PROBE183_WIDTH-1:0]           probe183,
      input  [C_PROBE184_WIDTH-1:0]           probe184,
      input  [C_PROBE185_WIDTH-1:0]           probe185,
      input  [C_PROBE186_WIDTH-1:0]           probe186,
      input  [C_PROBE187_WIDTH-1:0]           probe187,
      input  [C_PROBE188_WIDTH-1:0]           probe188,
      input  [C_PROBE189_WIDTH-1:0]           probe189,
      input  [C_PROBE190_WIDTH-1:0]           probe190,
      input  [C_PROBE191_WIDTH-1:0]           probe191,
      input  [C_PROBE192_WIDTH-1:0]           probe192,
      input  [C_PROBE193_WIDTH-1:0]           probe193,
      input  [C_PROBE194_WIDTH-1:0]           probe194,
      input  [C_PROBE195_WIDTH-1:0]           probe195,
      input  [C_PROBE196_WIDTH-1:0]           probe196,
      input  [C_PROBE197_WIDTH-1:0]           probe197,
      input  [C_PROBE198_WIDTH-1:0]           probe198,
      input  [C_PROBE199_WIDTH-1:0]           probe199,
      input  [C_PROBE200_WIDTH-1:0]           probe200,
      input  [C_PROBE201_WIDTH-1:0]           probe201,
      input  [C_PROBE202_WIDTH-1:0]           probe202,
      input  [C_PROBE203_WIDTH-1:0]           probe203,
      input  [C_PROBE204_WIDTH-1:0]           probe204,
      input  [C_PROBE205_WIDTH-1:0]           probe205,
      input  [C_PROBE206_WIDTH-1:0]           probe206,
      input  [C_PROBE207_WIDTH-1:0]           probe207,
      input  [C_PROBE208_WIDTH-1:0]           probe208,
      input  [C_PROBE209_WIDTH-1:0]           probe209,
      input  [C_PROBE210_WIDTH-1:0]           probe210,
      input  [C_PROBE211_WIDTH-1:0]           probe211,
      input  [C_PROBE212_WIDTH-1:0]           probe212,
      input  [C_PROBE213_WIDTH-1:0]           probe213,
      input  [C_PROBE214_WIDTH-1:0]           probe214,
      input  [C_PROBE215_WIDTH-1:0]           probe215,
      input  [C_PROBE216_WIDTH-1:0]           probe216,
      input  [C_PROBE217_WIDTH-1:0]           probe217,
      input  [C_PROBE218_WIDTH-1:0]           probe218,
      input  [C_PROBE219_WIDTH-1:0]           probe219,
      input  [C_PROBE220_WIDTH-1:0]           probe220,
      input  [C_PROBE221_WIDTH-1:0]           probe221,
      input  [C_PROBE222_WIDTH-1:0]           probe222,
      input  [C_PROBE223_WIDTH-1:0]           probe223,
      input  [C_PROBE224_WIDTH-1:0]           probe224,
      input  [C_PROBE225_WIDTH-1:0]           probe225,
      input  [C_PROBE226_WIDTH-1:0]           probe226,
      input  [C_PROBE227_WIDTH-1:0]           probe227,
      input  [C_PROBE228_WIDTH-1:0]           probe228,
      input  [C_PROBE229_WIDTH-1:0]           probe229,
      input  [C_PROBE230_WIDTH-1:0]           probe230,
      input  [C_PROBE231_WIDTH-1:0]           probe231,
      input  [C_PROBE232_WIDTH-1:0]           probe232,
      input  [C_PROBE233_WIDTH-1:0]           probe233,
      input  [C_PROBE234_WIDTH-1:0]           probe234,
      input  [C_PROBE235_WIDTH-1:0]           probe235,
      input  [C_PROBE236_WIDTH-1:0]           probe236,
      input  [C_PROBE237_WIDTH-1:0]           probe237,
      input  [C_PROBE238_WIDTH-1:0]           probe238,
      input  [C_PROBE239_WIDTH-1:0]           probe239,
      input  [C_PROBE240_WIDTH-1:0]           probe240,
      input  [C_PROBE241_WIDTH-1:0]           probe241,
      input  [C_PROBE242_WIDTH-1:0]           probe242,
      input  [C_PROBE243_WIDTH-1:0]           probe243,
      input  [C_PROBE244_WIDTH-1:0]           probe244,
      input  [C_PROBE245_WIDTH-1:0]           probe245,
      input  [C_PROBE246_WIDTH-1:0]           probe246,
      input  [C_PROBE247_WIDTH-1:0]           probe247,
      input  [C_PROBE248_WIDTH-1:0]           probe248,
      input  [C_PROBE249_WIDTH-1:0]           probe249,
      input  [C_PROBE250_WIDTH-1:0]           probe250,
      input  [C_PROBE251_WIDTH-1:0]           probe251,
      input  [C_PROBE252_WIDTH-1:0]           probe252,
      input  [C_PROBE253_WIDTH-1:0]           probe253,
      input  [C_PROBE254_WIDTH-1:0]           probe254,
      input  [C_PROBE255_WIDTH-1:0]           probe255,
      input  [C_PROBE256_WIDTH-1:0]           probe256,
      input  [C_PROBE257_WIDTH-1:0]           probe257,
      input  [C_PROBE258_WIDTH-1:0]           probe258,
      input  [C_PROBE259_WIDTH-1:0]           probe259,
      input  [C_PROBE260_WIDTH-1:0]           probe260,
      input  [C_PROBE261_WIDTH-1:0]           probe261,
      input  [C_PROBE262_WIDTH-1:0]           probe262,
      input  [C_PROBE263_WIDTH-1:0]           probe263,
      input  [C_PROBE264_WIDTH-1:0]           probe264,
      input  [C_PROBE265_WIDTH-1:0]           probe265,
      input  [C_PROBE266_WIDTH-1:0]           probe266,
      input  [C_PROBE267_WIDTH-1:0]           probe267,
      input  [C_PROBE268_WIDTH-1:0]           probe268,
      input  [C_PROBE269_WIDTH-1:0]           probe269,
      input  [C_PROBE270_WIDTH-1:0]           probe270,
      input  [C_PROBE271_WIDTH-1:0]           probe271,
      input  [C_PROBE272_WIDTH-1:0]           probe272,
      input  [C_PROBE273_WIDTH-1:0]           probe273,
      input  [C_PROBE274_WIDTH-1:0]           probe274,
      input  [C_PROBE275_WIDTH-1:0]           probe275,
      input  [C_PROBE276_WIDTH-1:0]           probe276,
      input  [C_PROBE277_WIDTH-1:0]           probe277,
      input  [C_PROBE278_WIDTH-1:0]           probe278,
      input  [C_PROBE279_WIDTH-1:0]           probe279,
      input  [C_PROBE280_WIDTH-1:0]           probe280,
      input  [C_PROBE281_WIDTH-1:0]           probe281,
      input  [C_PROBE282_WIDTH-1:0]           probe282,
      input  [C_PROBE283_WIDTH-1:0]           probe283,
      input  [C_PROBE284_WIDTH-1:0]           probe284,
      input  [C_PROBE285_WIDTH-1:0]           probe285,
      input  [C_PROBE286_WIDTH-1:0]           probe286,
      input  [C_PROBE287_WIDTH-1:0]           probe287,
      input  [C_PROBE288_WIDTH-1:0]           probe288,
      input  [C_PROBE289_WIDTH-1:0]           probe289,
      input  [C_PROBE290_WIDTH-1:0]           probe290,
      input  [C_PROBE291_WIDTH-1:0]           probe291,
      input  [C_PROBE292_WIDTH-1:0]           probe292,
      input  [C_PROBE293_WIDTH-1:0]           probe293,
      input  [C_PROBE294_WIDTH-1:0]           probe294,
      input  [C_PROBE295_WIDTH-1:0]           probe295,
      input  [C_PROBE296_WIDTH-1:0]           probe296,
      input  [C_PROBE297_WIDTH-1:0]           probe297,
      input  [C_PROBE298_WIDTH-1:0]           probe298,
      input  [C_PROBE299_WIDTH-1:0]           probe299,
      input  [C_PROBE300_WIDTH-1:0]           probe300,
      input  [C_PROBE301_WIDTH-1:0]           probe301,
      input  [C_PROBE302_WIDTH-1:0]           probe302,
      input  [C_PROBE303_WIDTH-1:0]           probe303,
      input  [C_PROBE304_WIDTH-1:0]           probe304,
      input  [C_PROBE305_WIDTH-1:0]           probe305,
      input  [C_PROBE306_WIDTH-1:0]           probe306,
      input  [C_PROBE307_WIDTH-1:0]           probe307,
      input  [C_PROBE308_WIDTH-1:0]           probe308,
      input  [C_PROBE309_WIDTH-1:0]           probe309,
      input  [C_PROBE310_WIDTH-1:0]           probe310,
      input  [C_PROBE311_WIDTH-1:0]           probe311,
      input  [C_PROBE312_WIDTH-1:0]           probe312,
      input  [C_PROBE313_WIDTH-1:0]           probe313,
      input  [C_PROBE314_WIDTH-1:0]           probe314,
      input  [C_PROBE315_WIDTH-1:0]           probe315,
      input  [C_PROBE316_WIDTH-1:0]           probe316,
      input  [C_PROBE317_WIDTH-1:0]           probe317,
      input  [C_PROBE318_WIDTH-1:0]           probe318,
      input  [C_PROBE319_WIDTH-1:0]           probe319,
      input  [C_PROBE320_WIDTH-1:0]           probe320,
      input  [C_PROBE321_WIDTH-1:0]           probe321,
      input  [C_PROBE322_WIDTH-1:0]           probe322,
      input  [C_PROBE323_WIDTH-1:0]           probe323,
      input  [C_PROBE324_WIDTH-1:0]           probe324,
      input  [C_PROBE325_WIDTH-1:0]           probe325,
      input  [C_PROBE326_WIDTH-1:0]           probe326,
      input  [C_PROBE327_WIDTH-1:0]           probe327,
      input  [C_PROBE328_WIDTH-1:0]           probe328,
      input  [C_PROBE329_WIDTH-1:0]           probe329,
      input  [C_PROBE330_WIDTH-1:0]           probe330,
      input  [C_PROBE331_WIDTH-1:0]           probe331,
      input  [C_PROBE332_WIDTH-1:0]           probe332,
      input  [C_PROBE333_WIDTH-1:0]           probe333,
      input  [C_PROBE334_WIDTH-1:0]           probe334,
      input  [C_PROBE335_WIDTH-1:0]           probe335,
      input  [C_PROBE336_WIDTH-1:0]           probe336,
      input  [C_PROBE337_WIDTH-1:0]           probe337,
      input  [C_PROBE338_WIDTH-1:0]           probe338,
      input  [C_PROBE339_WIDTH-1:0]           probe339,
      input  [C_PROBE340_WIDTH-1:0]           probe340,
      input  [C_PROBE341_WIDTH-1:0]           probe341,
      input  [C_PROBE342_WIDTH-1:0]           probe342,
      input  [C_PROBE343_WIDTH-1:0]           probe343,
      input  [C_PROBE344_WIDTH-1:0]           probe344,
      input  [C_PROBE345_WIDTH-1:0]           probe345,
      input  [C_PROBE346_WIDTH-1:0]           probe346,
      input  [C_PROBE347_WIDTH-1:0]           probe347,
      input  [C_PROBE348_WIDTH-1:0]           probe348,
      input  [C_PROBE349_WIDTH-1:0]           probe349,
      input  [C_PROBE350_WIDTH-1:0]           probe350,
      input  [C_PROBE351_WIDTH-1:0]           probe351,
      input  [C_PROBE352_WIDTH-1:0]           probe352,
      input  [C_PROBE353_WIDTH-1:0]           probe353,
      input  [C_PROBE354_WIDTH-1:0]           probe354,
      input  [C_PROBE355_WIDTH-1:0]           probe355,
      input  [C_PROBE356_WIDTH-1:0]           probe356,
      input  [C_PROBE357_WIDTH-1:0]           probe357,
      input  [C_PROBE358_WIDTH-1:0]           probe358,
      input  [C_PROBE359_WIDTH-1:0]           probe359,
      input  [C_PROBE360_WIDTH-1:0]           probe360,
      input  [C_PROBE361_WIDTH-1:0]           probe361,
      input  [C_PROBE362_WIDTH-1:0]           probe362,
      input  [C_PROBE363_WIDTH-1:0]           probe363,
      input  [C_PROBE364_WIDTH-1:0]           probe364,
      input  [C_PROBE365_WIDTH-1:0]           probe365,
      input  [C_PROBE366_WIDTH-1:0]           probe366,
      input  [C_PROBE367_WIDTH-1:0]           probe367,
      input  [C_PROBE368_WIDTH-1:0]           probe368,
      input  [C_PROBE369_WIDTH-1:0]           probe369,
      input  [C_PROBE370_WIDTH-1:0]           probe370,
      input  [C_PROBE371_WIDTH-1:0]           probe371,
      input  [C_PROBE372_WIDTH-1:0]           probe372,
      input  [C_PROBE373_WIDTH-1:0]           probe373,
      input  [C_PROBE374_WIDTH-1:0]           probe374,
      input  [C_PROBE375_WIDTH-1:0]           probe375,
      input  [C_PROBE376_WIDTH-1:0]           probe376,
      input  [C_PROBE377_WIDTH-1:0]           probe377,
      input  [C_PROBE378_WIDTH-1:0]           probe378,
      input  [C_PROBE379_WIDTH-1:0]           probe379,
      input  [C_PROBE380_WIDTH-1:0]           probe380,
      input  [C_PROBE381_WIDTH-1:0]           probe381,
      input  [C_PROBE382_WIDTH-1:0]           probe382,
      input  [C_PROBE383_WIDTH-1:0]           probe383,
      input  [C_PROBE384_WIDTH-1:0]           probe384,
      input  [C_PROBE385_WIDTH-1:0]           probe385,
      input  [C_PROBE386_WIDTH-1:0]           probe386,
      input  [C_PROBE387_WIDTH-1:0]           probe387,
      input  [C_PROBE388_WIDTH-1:0]           probe388,
      input  [C_PROBE389_WIDTH-1:0]           probe389,
      input  [C_PROBE390_WIDTH-1:0]           probe390,
      input  [C_PROBE391_WIDTH-1:0]           probe391,
      input  [C_PROBE392_WIDTH-1:0]           probe392,
      input  [C_PROBE393_WIDTH-1:0]           probe393,
      input  [C_PROBE394_WIDTH-1:0]           probe394,
      input  [C_PROBE395_WIDTH-1:0]           probe395,
      input  [C_PROBE396_WIDTH-1:0]           probe396,
      input  [C_PROBE397_WIDTH-1:0]           probe397,
      input  [C_PROBE398_WIDTH-1:0]           probe398,
      input  [C_PROBE399_WIDTH-1:0]           probe399,
      input  [C_PROBE400_WIDTH-1:0]           probe400,
      input  [C_PROBE401_WIDTH-1:0]           probe401,
      input  [C_PROBE402_WIDTH-1:0]           probe402,
      input  [C_PROBE403_WIDTH-1:0]           probe403,
      input  [C_PROBE404_WIDTH-1:0]           probe404,
      input  [C_PROBE405_WIDTH-1:0]           probe405,
      input  [C_PROBE406_WIDTH-1:0]           probe406,
      input  [C_PROBE407_WIDTH-1:0]           probe407,
      input  [C_PROBE408_WIDTH-1:0]           probe408,
      input  [C_PROBE409_WIDTH-1:0]           probe409,
      input  [C_PROBE410_WIDTH-1:0]           probe410,
      input  [C_PROBE411_WIDTH-1:0]           probe411,
      input  [C_PROBE412_WIDTH-1:0]           probe412,
      input  [C_PROBE413_WIDTH-1:0]           probe413,
      input  [C_PROBE414_WIDTH-1:0]           probe414,
      input  [C_PROBE415_WIDTH-1:0]           probe415,
      input  [C_PROBE416_WIDTH-1:0]           probe416,
      input  [C_PROBE417_WIDTH-1:0]           probe417,
      input  [C_PROBE418_WIDTH-1:0]           probe418,
      input  [C_PROBE419_WIDTH-1:0]           probe419,
      input  [C_PROBE420_WIDTH-1:0]           probe420,
      input  [C_PROBE421_WIDTH-1:0]           probe421,
      input  [C_PROBE422_WIDTH-1:0]           probe422,
      input  [C_PROBE423_WIDTH-1:0]           probe423,
      input  [C_PROBE424_WIDTH-1:0]           probe424,
      input  [C_PROBE425_WIDTH-1:0]           probe425,
      input  [C_PROBE426_WIDTH-1:0]           probe426,
      input  [C_PROBE427_WIDTH-1:0]           probe427,
      input  [C_PROBE428_WIDTH-1:0]           probe428,
      input  [C_PROBE429_WIDTH-1:0]           probe429,
      input  [C_PROBE430_WIDTH-1:0]           probe430,
      input  [C_PROBE431_WIDTH-1:0]           probe431,
      input  [C_PROBE432_WIDTH-1:0]           probe432,
      input  [C_PROBE433_WIDTH-1:0]           probe433,
      input  [C_PROBE434_WIDTH-1:0]           probe434,
      input  [C_PROBE435_WIDTH-1:0]           probe435,
      input  [C_PROBE436_WIDTH-1:0]           probe436,
      input  [C_PROBE437_WIDTH-1:0]           probe437,
      input  [C_PROBE438_WIDTH-1:0]           probe438,
      input  [C_PROBE439_WIDTH-1:0]           probe439,
      input  [C_PROBE440_WIDTH-1:0]           probe440,
      input  [C_PROBE441_WIDTH-1:0]           probe441,
      input  [C_PROBE442_WIDTH-1:0]           probe442,
      input  [C_PROBE443_WIDTH-1:0]           probe443,
      input  [C_PROBE444_WIDTH-1:0]           probe444,
      input  [C_PROBE445_WIDTH-1:0]           probe445,
      input  [C_PROBE446_WIDTH-1:0]           probe446,
      input  [C_PROBE447_WIDTH-1:0]           probe447,
      input  [C_PROBE448_WIDTH-1:0]           probe448,
      input  [C_PROBE449_WIDTH-1:0]           probe449,
      input  [C_PROBE450_WIDTH-1:0]           probe450,
      input  [C_PROBE451_WIDTH-1:0]           probe451,
      input  [C_PROBE452_WIDTH-1:0]           probe452,
      input  [C_PROBE453_WIDTH-1:0]           probe453,
      input  [C_PROBE454_WIDTH-1:0]           probe454,
      input  [C_PROBE455_WIDTH-1:0]           probe455,
      input  [C_PROBE456_WIDTH-1:0]           probe456,
      input  [C_PROBE457_WIDTH-1:0]           probe457,
      input  [C_PROBE458_WIDTH-1:0]           probe458,
      input  [C_PROBE459_WIDTH-1:0]           probe459,
      input  [C_PROBE460_WIDTH-1:0]           probe460,
      input  [C_PROBE461_WIDTH-1:0]           probe461,
      input  [C_PROBE462_WIDTH-1:0]           probe462,
      input  [C_PROBE463_WIDTH-1:0]           probe463,
      input  [C_PROBE464_WIDTH-1:0]           probe464,
      input  [C_PROBE465_WIDTH-1:0]           probe465,
      input  [C_PROBE466_WIDTH-1:0]           probe466,
      input  [C_PROBE467_WIDTH-1:0]           probe467,
      input  [C_PROBE468_WIDTH-1:0]           probe468,
      input  [C_PROBE469_WIDTH-1:0]           probe469,
      input  [C_PROBE470_WIDTH-1:0]           probe470,
      input  [C_PROBE471_WIDTH-1:0]           probe471,
      input  [C_PROBE472_WIDTH-1:0]           probe472,
      input  [C_PROBE473_WIDTH-1:0]           probe473,
      input  [C_PROBE474_WIDTH-1:0]           probe474,
      input  [C_PROBE475_WIDTH-1:0]           probe475,
      input  [C_PROBE476_WIDTH-1:0]           probe476,
      input  [C_PROBE477_WIDTH-1:0]           probe477,
      input  [C_PROBE478_WIDTH-1:0]           probe478,
      input  [C_PROBE479_WIDTH-1:0]           probe479,
      input  [C_PROBE480_WIDTH-1:0]           probe480,
      input  [C_PROBE481_WIDTH-1:0]           probe481,
      input  [C_PROBE482_WIDTH-1:0]           probe482,
      input  [C_PROBE483_WIDTH-1:0]           probe483,
      input  [C_PROBE484_WIDTH-1:0]           probe484,
      input  [C_PROBE485_WIDTH-1:0]           probe485,
      input  [C_PROBE486_WIDTH-1:0]           probe486,
      input  [C_PROBE487_WIDTH-1:0]           probe487,
      input  [C_PROBE488_WIDTH-1:0]           probe488,
      input  [C_PROBE489_WIDTH-1:0]           probe489,
      input  [C_PROBE490_WIDTH-1:0]           probe490,
      input  [C_PROBE491_WIDTH-1:0]           probe491,
      input  [C_PROBE492_WIDTH-1:0]           probe492,
      input  [C_PROBE493_WIDTH-1:0]           probe493,
      input  [C_PROBE494_WIDTH-1:0]           probe494,
      input  [C_PROBE495_WIDTH-1:0]           probe495,
      input  [C_PROBE496_WIDTH-1:0]           probe496,
      input  [C_PROBE497_WIDTH-1:0]           probe497,
      input  [C_PROBE498_WIDTH-1:0]           probe498,
      input  [C_PROBE499_WIDTH-1:0]           probe499,
      input  [C_PROBE500_WIDTH-1:0]           probe500,
      input  [C_PROBE501_WIDTH-1:0]           probe501,
      input  [C_PROBE502_WIDTH-1:0]           probe502,
      input  [C_PROBE503_WIDTH-1:0]           probe503,
      input  [C_PROBE504_WIDTH-1:0]           probe504,
      input  [C_PROBE505_WIDTH-1:0]           probe505,
      input  [C_PROBE506_WIDTH-1:0]           probe506,
      input  [C_PROBE507_WIDTH-1:0]           probe507,
      input  [C_PROBE508_WIDTH-1:0]           probe508,
      input  [C_PROBE509_WIDTH-1:0]           probe509,
      input  [C_PROBE510_WIDTH-1:0]           probe510,
      input  [C_PROBE511_WIDTH-1:0]           probe511,
