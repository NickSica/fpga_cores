`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 19696)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5DWIWhnhqhOGvj3OuNtw9qgJrBWHcT4pImUXhQTKfS1z43z7L8LEU1Ox
TZ+rBsr1aIUeqHr1CDCqJ+ZIZNBQ/pbfpjcxZSWykq7cnQSgJ/QQIiusolc4Wv3PjqlTr4De0AJG
3MfFNGbFAoMn2qM28c3MPLVwJBXeotwSU1RFSDY7Vf7UD6HsKqRLGB8J6tKWNpwPHuxgjXcYpToq
phs753YOKTNNIPJdSfx5snBkGdTpDdkxHYURjbPO5+1dGZq6OINuLejxrTV747JN/NP92YXn71aq
qo/bgfLUFwt1oxqe9Z0ugjYZKvEOiUgkPwNj+TnU/ApKvjI+GHME+F6voP18k1w0zjbYYeozaklD
ar/JKu1I8yJYQSqOSDaybp9njVFNhimKy+a0gwaRZ5pHDrwNQQcnjxTxEscPr4CASTHubgitzCrU
eSB17CaaxsalgBIMeAhR4Yp4ExnLQp5jCegXfbFvHgLrK9Fey18A8ZZ/PguU4xWi/nirtCOLKCak
Np2F/xCESnse5QlgcVTSAnzhAYU5TbFgLsIAXivqUBAONZIRoeYR17Q/1XH1sBWwfcaM2egglFey
b9ofwMzQVY8pC7v63Ed6NiIb2zk10YqMWNgd4OXhJolM2Vnl/O8xIXOWmJWx9N4NRiq2b08BjJRG
f++aWbC9qw3iJp/pZK73hnwuopzXM9o4DtLUa1qhmPZBeEKEI5WadHuSO8ylMzbW617DthGH0ux/
jI4ULf1KMwOJ2iS7m75Q3jHBureKaX+k82y7HYTF88B/2swGUFewKBKfWYqBaK18ra1OWSWTwYff
IIf3wcfq4wUNUuGFYhI7e+NhRiHDPft2EW3yUM2gLdElcVv4y1aUKYxPht9dEyQeXfDh8zwX0Pa6
I9XoNJ/5ninSLSQCEQhe6QaJq95lLANC7vey/xg1rep+t6NloydwVyddBTVnwB7Hx5jSDb4QJzGG
z7g7QrWsgu+MM6/2NtGrr7ZA8Aj2M1zixtyYq2tJiZJ5QiqeKbPmgHHdjRnEkFg6Q6vgYrTvjF2+
2jFXsQPjkZDeiG/vVNpKHi7BHt9qoJa7cRxENkDyPuGMAj7eoEI+9vuSnSlZuz5MXUV8eexLn+p4
CaekvtscCTj9tMqUkOzAXCJD5nrCbsNQV7oyK2TIzLWDYQ22JqFXh3SGR/Ez61U/yTv9M2buPS6q
/F7Zd3JH6Yw2fPnk5UT+O1fvHVugP1CFOjHqpm+Vs1cTIQkNEf7EAfi80/qaqzZprC4emb7TP89R
5ZrWIxDVc/+ZaDAUtb6QjAI3kfQTc8X6pUpi3EsgJOAcslbGWJwaS+cSDue+NeeSQT9zpCec8vFP
BfTHFIa0t2W1FKe3wwm2cCQgPOPFh8Vp4M6gPGiEcUQ33mFaqvJRIQiWxj5XsagDXQxkS/Iu6D5k
KPCBmE9ixG3rxK0N49aI87GAAlEmAZbyJKQZ0H6sdjtOJfcwmmB+qXVW90Ae/jpgDTg2qWjvftFq
yjllQyJtPJVODtSXB94ZiAcZBhqNvKMIg64pBCUR04EPAqQQXS9E+W64gdNnzTiCBUYJPVwUG8i+
qwCn0j6/1uKJwiGA+4dGMyxoperCHuWsLm8lfTgQzdzCunXYClN54sXYC8GppDTbdhDXm8RUw4ai
dsBMF8636k1p/3d1D7f7UE2PKG0e9c2zMe5B/+A97O1ZxlsIEwbZ7GTWWVRajXtrGdWmA5QQRNR0
c6OlWMRbicOtmDBYqoPavUyTVlZPmGa1V/sy2xgWJ5c1Mz7DIe+EgmZflI8Rf/E3O0nYYmrvUZo0
yxEDi3pwJYUyDqDUBxoAkuzD00OfcqVTjTmELyJKFqF2Otfyx7GKI3+sF3LJda9wOwRl7wzbYhhM
pCC+8RB6+E46Pp4xjJSGjr5MGbCvBC+lk4pLIn9/uGChCHuqnZTM3Gac/O8fUdVfE8Gid2GJ+mAO
fZUotpwGDNHlzViQgpqvQrCXLXgMG+uK+R4qLYlijl9xJWSRxTs7tBJZ/JbtanNwgav7BYzbTVLG
DTsNVz6AD2JjZf6wLVq9Kd/mA2vgRvwDLlBRApfOzVBarlAa03jA/HzopdiCLphv3vhODhm/hKcY
VNonu/tcy/bf7r5kWMuZXV3XbcZowavPtBbtYr+/UZbhUvun372g0bSwor6tiLDikCj5dC8iYFLp
uu0oMFVwOWRJk3ylAR47Sx5HXXeZMEr/UvTpRx7Jby+tJ2rHePbdh/LoT91zT4TmMyMKCH4b9w02
mnGnG0ez94S30vKBTPT05BGb4G1TQyUDIMp+gYHiWKkrddhdGZVjUxX0j8d+BkllDMLDG8odUOwo
LqpMmNBLoXxEtMVO3tILZc7LjSatMN/IThJgmVo/rvb+iaAkLmrGgJKCjUQWGu0rf5wY8ojzMdEh
AE/pGwCjOF/r68af0plEpW80UH+df4nysP61tdWXiyMAza8ZGaAYxRWqNgo/6e2V/jGZ53LR+xWY
mzek6vvo60nSvikjJpwA3SXecnLKI5ReXVbkjIIY5lp/9AqPQXlbtl97+hbWO4oUDCoOOXLuzEAh
qOaiK8yAVWfcwi2bqbjXymDMMyivJG0sdI5LcQnqwGSImYr3lHOSkeFAnghUZ02IxbRYHmbuL4IG
Ugf3nNiem29I4eXVXcGusOnuKGvRij4AOfjPD2i8Rwj8XYulhusBvPilyEWFNgJdbG1ngLwSbt4z
4RXM652KKBstJQMjkzbzdFWMCfvmOCiZOoSRZxv0puYE1WGX1dcO9Qdtfq1M6+VvP4ygN9PYU7yy
TeV2SQnNpQqPEhSt+pg5FgR3IVXnmSSBUZpucfKKUE9KGNATqs4g6Y8mnkjHBNiU3vOPYF5Cpo6o
a4IFur2N7dhZjcd4NhpXtKnImZ8iO6PQLuuTxXAJ1LC0c3+4tH/VunZ5G0lWUUJNrCOGcyjisgY1
/Fi0cBoZ5l5X8Hs+yrX/MlPJefsclIaOc2K3WnhVpb1yO1g06K9TcbIIx8/Ltjxq4sDj9xVrMwNv
tqMiMVdYbRm6zNjEzVcGQS1MFfJ06enb6KPJ3c2ravYKYXeHO/1JxNG85YDyhGqisBk5I5Gvdh3I
oIDmEryGjap3+R8zYpMeboA+J/5KhRU3v5Jl1iB6LRu59sQjHWJnLffbk3ORH4k8FDsgs9+qL8z+
gPvDqHM7/zOK8ai+0LOirQyousvg6PXUVW3zmuPzN6wpeKGFuEDwi5SpSdRk5H0miG4M7NME/uOW
pZkvcGNflMvJzOGzRDnsgDMuuQ+T34N/kRhutiv5x5FcePfyav/bxOeTltHH/snBNmiHdASFJCIs
DmdGsG8N+JhQBqWhkRv5ltpA7LYmiMLxlx5B6odIq48ts6670v2LMsZsSbUGWQ21ztM6CO3OwC+Q
rY4httu2fxmQ/Yh3qTkgElh3+doLI/9+UVdZrf9fHRSAcBJR/y9jqO359pBlGTGOP7sROkUpY+iN
vhtQRJ+p2iyhMehfOvWMbZWh1TrK9Ip0zySKTYnwHMUOtR4DDDyE8hoD76Me1L/SVwHxc4qbxpoF
sVsDe21dh9cXGNZR+Ac9Vdg3Tk2tgwEM8/SlDuMgCF+ZWxCLbTiZrFZPfLvggHDgWv/Vb2Uz19YI
T6UmfFLdYHGU6CDNpDJ1hmtC95VEvw+vHOHooZiSxMhAxDvbeYbtIErB/lKhPEI5OM9gzryGzvqz
uNdvDGHCOGAX3xBaVR5ioJ1THYQg6BxUawCBP5DeZd6dnDmpVI7bd4+rWuCNccb/K6Y3B4efgzo6
rJid7EuqdlrFHO6EPr+FwjoDBLzhU8WRrqturIyXOFDQpltDYCPfJHYSRguXDfgPM+n8ZMAyB6ej
7wiYz8bu/A0bvF9bSG6g6lL5D9swwZYsj3DPT+VmGTJquO+0X1TAQIgBge35P6dkNqy/WsdTCdGE
IScIfyljxU3UBFa7OckvwjVwBXjNOl1ssM3FYl0vsx9/ovXsxhZGVNX7nNw4phbnHLAYI2UBd/b6
DUuv9afRDLDPH0EOrp4zEzFggtIz7wP0mZZRNcicsUkGc6cNPrz0/l44vEQ7cCxUSCDYpdyPtZnx
TVw4rpacsyXqyu6J4BRcr4whn3i8n5pe419JM2EQko4Je/eFAFuJhfHiXy8EyDXRQv8WKlpikrYP
fjnM31h5iXOtVys9VLfSSymLup8zf2XBE4sCelW2zAZ+cuhkDw7pjKHxX6i80/TQnGwHl24ZlTJM
5MZ6hkwLyGv14F3UunzLESxnlf2EFItyGTOgXp+B6P8ZYkaSM17zUpCAzNLW6nlGMlS1lpaKkmwS
XX2q2ICyohPpx6dr7UHw/7w7yf/gz+vCLYwj/bRpcPCOtkUWlx4fK56LzhyEJ4Zt/N2XSQc5Xoj7
82SbXb/aEOjl+2mesthKABqPebpzcR7LzQ99sIpZzxETBgfSFsO8EJm90eGGioGPwYpEeMdKzVWm
xVN9z7Dh312D3TBJo199chiiVQCMzRMToSAICK27P/SOW5swyWKDKfCoMO9h0+AWRQ53n9p67AbI
B/v71/SD2nfPuYjsV4r/3sQ1iRf8smI8rLXZay7ZK3fpCLzK5QL0+zrYQImkfRMC9uqah+6/kTmJ
0RhPX8/xhrIA5A4NHP0yRbVXFu7OIDAxd6cw7BQGFTFuAZ2HQj5doRIqaQEJFmAHM6gmh4dBGf+k
bxvsS1JOfYL610pxEUVHTjKAAuEUStym7J2cMcJJUL9UvXg1QP6CbNg6ZzKYy3nIRp8CmzctRe5s
1Pq2GdOCTYtJ2+I+8iWVVf8L+LJ9/9jVpfpj+gFWkYkBAZV85AChdeKdyHjQbdYCpoQP6Uwq0Rzj
xdVYE7TR4Jw1Nwir9S/KnPGmy9xpQhpnu7mFYjLdKHDOrpDCjaA/V/GJOW7XuhcsVhCYPNLCt5D7
7mI8rigUmez4EbXz5I3KCseEcututtXP1Pyhr99n76QvzE03QegQqIRdr3i4F1+0icSPB+bB0rEf
Rhox/x/tIIE85c9X7mD/KqCDVKVjotQAnj+71//SfvfvFkKyDhJp4N4BrUF3eLJl69qus3oNZdhp
nXL+bS/baBa1qTfoDf7cLFyXV6IkuSQNZxQmS+XsZ6z3ZgZCKjRvXCrzOQvlj+kIw9TQTdsBV2UB
bW0ViXwhixH/OtCL0+a/LqCbwSNeoWCHhO1i98CAp2AShfXJAT/AnO7ihmv6fLnv9olR2BxEmnzV
mjojien7vCUAXHjY8TSe0gDiQFKVl1Yq4IDvAAcmWVTjWl8XnmHzvNR9vzdhT9OB/n5tHNyRxwVt
sB/Fneho1P4kvnkQFHkm/wzrTgsaJVFR4AOsMAX0K7zw+sO+uZ7hyhPKRTPfoLtp2X3rzrq9+qZQ
zByHlCIR5dbXEBM/raMV3lAShX5/NVI8UFeTSUaVzPaZV+yUSW0K0cCkooLp5uSIwyGN+a+guOjT
yt0Gjx5Y8HyVLcZ065FGaUTZvdKS06P9/T29IQ+hina/n7Minw8Hd+ZS9ERFZw5iT6fcU7tugasi
idn/IwobBhxSOuNE4YuBzaiz+6Am5OXO2Rfu3PGyglnZ6iyeT0q9Fb1HGLbLUZ4b5FS9yGrqZv8W
kHQpNDUtWDEOYrD+uMcRdaD3PhXD1e/se0I1GIsTCmGKhlq6PsSoCn0z0Pxuz+OqW37qM1hazRhG
ZWXcNSCf+MshVMYsackHMc6jVedKLTq9+h1mElYlZgpkphCqK1YxX3n+7pRmRYuZW0ej0WlwrRlq
bA/CgT+AEKjsIUXXW0ZttzPkdsvBymKaVin2YeORnFbCCw+q/fR7fTbNyzODW860Jbo227bb1uM+
CaMvfvIp0UpFgPLy8AnYoJ78I+oTBEDtlHFn81kGEdRKQ6mdlE8hcgxLLFRiv6p+Qy8+nr32UnJ3
ymxuYvMKit72eQK1B4ykCwIIGm7ZSvE/+qRdVUNNtswjxzEZGnpQB1za0Rz3xTFQ534SMSxLd5j+
lqPa+OI6c4mhGoqP5TKwwWYTOz66bu4Lo5js70bRt8J4OF/sBHvpByt/IRAx7QfxOHVhkYctjlc3
LvCO03yWGaHlWwa8nK7PAtW9e9fKfY9kgpXAYyr7sISEEbD5t8KMGG0zHiO003o33kGsy9ZO5Obv
ryK6nKHxp8TF1ujIHRJSRW6QQQitJlIx+Y0fB0vaHEtn0LCVkzXhovSpP7O+ph+D7upIf8Z0/yKv
Dwqr9H4LEJhU3GI+n2SXH1yZxI0ioGW0tSgV2u0Rh52Cjpe4fRnlH6akRH0lMI4Ahb7NyRww2sbW
uTH/douH5JILTSZ4SlXrurt9rmj8TG0W8ridliXFTUfc5Gboo00m+7shxpqw4uC3W9ySHrI+wRrt
GhYtE4FGnil2xuoRY+PVrPJd9dZw3F8eXH4kE/5niANus15vQvr8PJ9wGrA8ku99HRRfwE66bggS
6IdHu02I3bcGXw9eieKfqNdxW0rTTbs9Rr+/srvVOImoFwtAORQ3ptFKBtF3foFUiBEWjR38JJvS
AMSjf7mqeSr3hQpLPJXk7Dob91matIHzJ+vw7gbJ/wXHLJL7HpYr4dFM5u0P3JG0T94nb6HJz7t2
GbmbOEvPB9J34KadBnKaGzRgHXZsEn5lR3yCFB8QGgfThpzTkqa8syQEbnttCGivTQKkz10m4sx3
lenh2NEgRlNO1NvJ1iGPh6AGKFM4MAAasbSR/K6g6G1JF/SaYDBTIM6UH4JwFaND7XPphe+CqWJn
nME87KSxfhlFbPnoiP7JYJFpw75/U3hB/IY5mXTqxsDQLpGPFEvIxyTJlmFqkIxAHAzrkSjFffns
10iwWoE2oqvtnfqcj88zAnobZ3JS3KztvG6i6LASlj+AXhvjAqZ/0brHuSZKeCCwid9W2YeJp1sS
ufua/pvVazpcSnaiIKFluaB+J7XJKPvRMdZV9D66ZoKG8yFESnugMcBSKqSviIWAnGD7vmSe7D4B
hfl4ojpRK0K0evftlml7weL5QSiW5YxI+rkGQn7O3zGryYAVfPECrUF5yPS6/eseZFdcd29QLtQE
//q+McZEz6mQA518sQRxQZEB2clpTMc+fjlGtZJcGcvBePcNKV3trMiKVoZQ7N6i2ekyzSCgffWC
MkA8qicsBLatnh0qowiaVZwqgD/fxLNHOJhiLRI2qpsc/Vpg5ZlyF6zqglfJm//lW/qXphIyZKSe
nd1S5dm8/iJGHZEpBrl671PbRs5ZH5/VNuvMgVrKbWFkkUXQliz42pEMLw+mKiDWYpbznN9Dwbj4
PKaP6rRRbl4bKiot7EIYFjqz4e8FhHdMbeIjYOQC/+Ey4BZS6yJs/Dx8MLB3ENJuBn/S6gEU2/h7
h9im1AQ6lHfrGMnslfIydUp9P4yUuoY6mjK1BpjrV0kmWMtKviU2t7OGu6OJVX61vgCYC1T9uN9j
oyYceRaeg35xbJx48s+l5oVTG4n+IYxbYCIx/7QVS8jGyurQa4oX8hlc6EfBATtWAPzODSP5l1dk
xAX1fCMreJXiaT/Jn8yIvtiYEDOAB0LPOneC+7nwOam/smHfZsV2f4Qik5eh9NBJzb0yYPbVUbf9
oC1hEKQbANoST6Heso+f4h807oy9a8yim8QWrxHlelBFFSLQPfCiGKye+M302cvfPkx3SSCF5nXG
511ag95qoN8Bywp744okXJ0DnoKEDaVJFFmo8t+5Fc3qq6ycKJynH/Tt9QocuLE9pI8zheQtFUhc
0slrxEO9sEXSqib+eZZxmFNVXUL7SAedI3TxBqXOcl1Lu/+H7sLmcmxJi8MjHIYvXL1Y+NoSshrd
C7syMqUKQLl9WUL6V7i9em1HWnKkn1asnPk7cSBNxxO4UmCSa2UgqD3OpafSlEZTHQWOoMRFK74b
7Bcug4hibKdC1OxwndYZo74h4vbB25O+99RN3KdRXORmtNHkQZasaZgweLsvzAova5nMHwaot0/X
L/80kjvB6nm7dN7jsWhI4Fg6ue7sDER41DPb2PU1pUiqPXd+ZKpDvWsszv5azwTqLbKB+2KOtnuG
WG7/hLVcLGOcK66Jk1OvI8NM9Yrr7XFUCZWKerxh6g8lvsi7fxgeEncyB8uCLgZek2FJHCEek4ek
nEl8jEed/rtsSbuc6zdoirCUrMJDdI2TcBmbbNYBkehJPkBjUt0V0OGtFLovNi0OzOJtAmffDdyh
+G53DcEmQI9JDknCsCXKNr78b84cfxrf1PZ3LPsxMRg7bn23ybp/jtdwW1TLcpBTaA73yAVoIsqN
KRoMy8JeywUAg7k6PRcdYw66bqdZsqH3zFHV3dAYebFCuo8Fcw1D38Qf7f/gHW0K6Egb/5VRpjBu
jj6HALL0dDYvQNygsUmtqr/4uGILgWd3jU3n/TLxO8USrPABEfvnh5DwKNgu3lhsKtWfh6LTFfgt
yptVo8GKkwqSqdF7sMIurq0Xynt+Y+Yg9qZf6BzqalRBMuollEc2eKcKj1TWbO1sGwVsSWtPcugg
iVBIN9M/5Vlc02HOJWlfZzeCFHUPcEYXsWp9uBrBsfFs8//Qf+pSTZjJSYdWHBScOxnF0Oq2x2lC
jgHFAxey0u/lOGAGICRDmYljGp9NWBCdl8ojkO6N5DKRec9LJ3U6+S1DpdkvLhGP1ut+9f8xxreh
nNV5Lz89qxGRggZzrTnOyYF0y0j75gP3G1tzdSYsiy97KVpCGS4jsCochRdRqD0MpH/hvvnZw1Bm
RNOwVQuAwHRQ2DdLlpXVZ8ye4N0HMlkQAq0odc8dNud2set3lZbZPKSzE5pzvQPSZhFrkztkzZse
EJST7JtECx/fyKVVeCaAc7/ZxrBFtTTxI+ft3eqQZj0t+rCRTnGo80N3rcuuez5bmz5g8eTf6O6x
XwoHxP8+NyBln5woe6UYeOzBdHyDWYEbufI9ALnZ8/w210mAzc0TkWHalA7QKbrghWohfJye1WKh
EdpdUIkgbmLKW8xtkJ1M6VvHN17UxueTH9f70wciHORefOSyyrNs+EPiYcTqVynYc8U1lqS2+836
Qt0+aJ1vXn/mbcRTqHXdiKsZcKl3DBCRqjV4oT1BjuC++JmdyqLzdB5I5DY4OP35IBfM1p5BBC39
mFx/9oixhxGIwuFoRgyel3p2aRZTSZcNxPipgMo6foAB/5p9Upv3VTw5ltbLkbVtWe5M75Lr+ZiL
FcaHJhGc2UtC6HPBu+Z1UXe+TrFxWOIi6kwlkE+kJicXlszbIy/QceDZdhnLj3BVBr/txv6ig6SL
40EYeIsnVW9sz0/j3O3jesclLoNQZr4vGpDalA9IOeuUi+f+kxG/9csxCifolkXrlNZ7HPQ/lYaf
AnsxBIqhRLrGOL2TFnbn/A2dw1mCiC5WTU4K2ZYqfDaSNcNRUSq09KlJTOfuxBMHQ9xTHIaZU8cC
WtCrfqO4SmFXvDYEjqfaQfLf4hviEAn567Fy+6pdrOlzJBetDvvRPFnpTo9nS+7NXIVPn9/a9iNl
GeIEsQ3D78y4Bwk7KhGJbF57XLOi/rUr6F+FiTGJRctympaltxNV6MaMD5IB5AAhUMUqYbR85jyv
enodPrZL8CFiehb8nJuWG3j8ARcv1fWIpAdo6hCnngfUB41NUd+tDjAeg37cdROuLzKAXdg6Lvjh
hpUjgqPA41KG2iEghKfB/wv62y0wxtD62ZBwG14QcRuURnS2qwMj0+CbpPpk4XyRj1O5ADFHFHy8
6DOqmhYBgBuVI6RUXGsXorfTuiMPhAOcCVMSnX+v2CLAY42U1RCvjh+aQ5lNxmvDqfqcqTBc2ZYI
N2hC5PANQWCvXU580qfKLqKGwlaBYmfc8H+WeqazvZYcVAKopAzJMst3DPmxvipYDOAp91zdcMzt
UzJlqkOsZ6XE6DmiXxgUMgIQK80bYg3xYTAhHZ3UluWHdN7iIXJ4tsEGtlN8gxsuiRh/+MPdD8Q5
hhmB9XVhUO+FpMaH5FrmdSQINNs/8NE2UB1S8Qy/qN9+w68WdJNW9ys/tLtp8iyVNa7EzxDRhpyl
iRH0vpvJ60Zt6EYHjcAfa1wLV1sfU50VaO6fia7wSYjjJp7BMCJnbSTuLHQB9+aszi/oTJnXx5Qr
e0dIQpVdLNnaKxdUFDrNCyUvGG7KAq3P47940xDVvPfWzjtRusaokiZDh2tQ3w6EreihzRodXkOd
q8RVxAgF34iyvesgbQEIWVa4k57yfkWiJccNc9gyQ+doyQFzDKVGZaEbyVHCsh5Ei1hy93NHfkTy
Z6/YcMJNNi7o7XOsGcpPtZTZyL8vVh64ZcbtPCjsmALf3QG4NkLHkfNJzjMUERryHAeuDJcCmNbK
qz6U8D55i/gnODC1bZaX7m8R3i7CBBngMaMDC4AAlq9Lb3FgSlEthxgFIV8CQ2LKXbLJvBSVXW0J
mAsoNoy0M7JNKFQtfL1knD4Tu0BhlEbhU5FisJRZkaIw7ktTXASmNUuxb1g+wG5DXQUJsTPrceWE
1DG2feKg8GwGg8bGIiM1eFF1CsGPa/7/WN0NPDDiDmaob7yAB4ixBSoHcTBVW2tmgZtqpzp/QC5A
LrbMTY2j8aUao0rp9EfzGKr4+h+qW7+ijizdNEUigVOYzyGXOBOw6HL6V2Oh6sQInzvbBFW+2YdD
u56YwCi/Fmh09dQ7h/VJvqbrZtlIcM0AgzA0fNOg5Q8pcdnqLxBpyV9BQMKTn5DUmAZYDBW7dRfW
q0FKNeqopNZ/IlG4lTt87t/V4dsNNNW4jjDjJen9drOjHROFln+Lmzc+MkV4Ta0T9/Nrf8y9i14W
y2lZflbGCP8Vis/HTIhy1TNuiBET1MBR5am474geUnccjvmSaeBDfa9JwpFYDfAuuT0Wm8s5uAhx
R1QBkocJmCAMinF7BoN3mFMxNc9P1ziDy2pEj/zHr8424XW6teOiVs/r4RZ0co9Je10lBbKPvVJU
2QOwXClQ68GLMWJ2NzpCUfFDodbySyYsIwQyJ9Re5lyInwpUPCaoDcbC6q/TjfXFwYdHRLuVafNl
gU1/GMl9UQvFALxr2IcHkJqfqx5vkf+nrHVOHnQaJbi3Q7hBpLBMB6REKrp23I0IIIzhA1tLrCoB
TChLz0DMjsYDywg3on3h9STpwKKBCPVM+/fKZku5GMLg1+VuU299JqD5MBfPQgwP5XMlClD/5iLo
j9++y81QjwJ14ucqOBRZSn0CPvd6CMBIyd8bv0tptmuV5o0nnxS7ajiNdM4Qes0cG66gIsxkJjvx
TM+fA1XHkfy32fiXGoxLMs/6jTUuKR1yFNXr3fwXZ/OzQ3uyK1ouHRVM5Sj0w98vTmOsC1Df+fVh
uYc2WtRsLetrTGCBjxKP0peaek17CIv2aN8v8yaO3S76CNfTIjju7f1PInDvSjCvXnXJB2mQkNy8
6p55mZWfSuRLPh6WeKGN5TqIHz7Lzf8qHOdjJnkf+7BjknfeyGAM6FLRo+kI152S8bR5cLK/3x8G
ruhcAIe2z+o4lqiqPM+OUDB30UcbBMKlBMEmBTSSnn+FwTgABmu/8PZjeVq6zTtq08yhxYJwehAl
oXub1NjtwXieidPFPUSHguz0akG/+3Lmz22WGosdTDBprPK+0wdkhadKEeHnOpvrnYcBsBzmDFQX
qpruY9NHinQ84+bPBCrM9B6oczQ7qH1tDlRQEyCqqjNT9FE9eWoxLFPI7h03ChmPHHk5ZN2lrQWZ
o4CBeqzx1Wqw29tODJwyBrLWkUlhi8aBPYh5Wc3mx75QKZuNynK4l1kDDYKPEN/8HXLCQ12/Fi66
zhSnicP/UPmdZzYVwVqFulzT4A6oj7yd7Drur07BtZy5UZHtVK9tNnBqxtF4lMOCqAuJzCBulfwB
q214Opu8/Hb7+yv1ZdC2NLF/KJNqk9BJxkp7PyWcausGVuIqGlR5iMC/AYADe1gkWtyR2hfZmH0j
/NRMXxxNwzujwNdo0GAtnpoZvlnscsZYh/HFikL0encmRNXf0UkbN20E7oc91FIDpzOnttF6j8aG
+sJmugjN5jytJl72AWeYbfE3G4oir7LwW8JNC35zWq5ZWWG8g7nyTg2a222sxczlVvhuR3hYP39o
3zxMJAzziSnMR9He6MrL07NCzDTN9zODdMFeqzT32AYFWsrJcO7aoQlrOX1ewDnp50KLXy3dbc93
ExYnNyhxmTKYDYNnSuWn16ak+r9cr72h4BQgZ8KvpOvcAO5rrfohX/cdX/ZGn5BbfWo9itooxQR3
j67aSOJIwC7TrTSGvK7Ln/J4wjIjE73cc5F/bTJceXwtOQK0sY0pS+ola0R5Y66+xmA6BoJULt5b
U0w6sLqz99AKFr1IY5qtwwnEt65xp8zr2PAot0YGyMFSRRueCnLRF9wSDHvA0z+uFEnaTND1AMbf
iMV+5kszJeDh4mDxOXp6RzG2YmIRXx7OnxSMwjg98BH3E5VUeK0BEy73wASAH8KCTXhIq/u/xmi4
Ij9GMctXmKn0NDnXMOC8D8hibWVXZYn8qOtggKLOuRpOd1CckEBD0NFBMEg69kaft7KZVFC+hjq1
xnIsjeVT09lFqklYmTA0No148/IOSn3kegpWgEq/1nsRcRXM4DD0x11CHrN7SnyirQ5S73GMOd4x
T/DB9HbTGpo4FnwlVBAR65BjnAL413KW9UREjRT6A1sd+PEt3BIrAGyn4IOnYkyfLFHscNaOMjwT
BhSwWecZbCr3jJmmA3f7lW33/vR30wjwIV+Auruiu7Kbar7QE2HtFHYwxW2esK/YErVBD0EhMVR8
3vh9PXtvmxf+2Q6OSefPIBZtojMikNCWtDrETMVW/H3vJn9KMmCIxVCNHZ3r6WBWQouMoQCBMsjY
QRsG1aaIHWEGR8aIYBwAS/Ws6ZiqIlC17DmxrGJibz3ixyBVLzv7QEw068YrvUbRRoN6p9VZy6hc
hOMu9GaZHq9zv1v1Jb0AMvJMVWABLP48UDtchmGQ1bqLk5Bd7jypr9rGWqtluCSpz+ZkE5cGWs7p
imCOd/TRwH9ilz/h+nBt3UV9FkxWtQMvZVUz/2H/eqBYQR9YvwBgWkSy9yVAk0qfq3AYZYs5YFjk
1G/mHWKSis/KPHLD8BbkyON3KK/ctrf/srAF/9ktjH7UsCsVxXjZf52GCVxCR0X9cEEYpPgUpRnm
BvuYDK1eDudD9RuRgkLAEd6cWjhx9+sb4ewR+WurFzjS/ExPVH2lkJnJFubFYvbo4PlbYInMyVOX
iB3Q2DDjA5f3wmJqoz9FpE8x/bGGP8jDgLCTz6JTE95SDNXad7sfCQ8DXPbq9BHWYp/sCOBjOFwK
yMYn3x1KOhyesUgxfo6PVLBkqmrGQbMtnAx17/KtkpNl19k31VvnCeJ6XQDUSXPmMtj3KBJnuk13
W8VMA7UAtLFPgy9mBfvGoFaKdWNLvYkXBCMcVOwKodvHFOyq47cBh8tq0/KgcMNjF4z7ta2s6MCg
NhCs6pyIVabMnxcXnu32zm4gmzEx/bMs5RCj3aFRkiozkwIL1OfOP3TQu5NU7aomWE2x7aHsuLaL
Y6jfBoFFkU3gPb4c+ryJ/TcpuRcom6gVKlZUUSezFawUPjl38huacHoQ89dNcXf5Mamxgl/BXgnE
NL+iEYPl8fwA5LVSDG6GtWpy8SepBgfbJN8MOCk9p8WQPkZfVk9x+3ofBqBQG4Ltw5byoVKC1/jK
L4ZxUwnC/2jbUCy3fLirmuP6YNxJJTxMsMdWAznjoX9U3TKi+SkUFTaZA35qA5XMdTyGHi1lgSEl
cYwAyQpKMiRp7e1bRvNo7WtUGdRacyKRhrdm9U3HPSWNI46fGNNOM57Dlzzp2gRSBZYD5zAO0KCc
D3OtwPX/Iv/UlYAn0jLjMagE3Xf+HY5RZSUHWDXGDcxg7F2jcpO6S905IFmghOJzqRrJQiNFo21e
wovi34H9OMxMPQETdCWbkZGf/2tmPCRCoMO6oHPCKIdWcRleNC+0LvHgpTL6b9DMtWhGqAGHOCFu
xCy8f6+TwDeLeHAyyaLWkE7r2A66HvVo0Kzhb/1DxDmQO0EEMUuNRnBBqWdevYapVMb8zLFLXU6d
3xQd6vqSlu01yw3cvML47dXRE63ycjIehBj6K1e3KQOVVGQHkZc5J/5atqIR+A45moB6Gdo78HlS
dpC8EKeWqdEsLS48xoe24jcmyxEZLfL6rmNAeHsoM35tqLzNR91mUsEtyTZcUuXs8qtYaVmwah6I
YBy/mg/h9aFqgKg1zdbZ0xyex05O4Jrxz266hzEPBgqV9/LF3Cnf/R98HUjCcJ8zDBiRmoEKvjIX
6ky3f37WuS6N5j/EZjiF4J4+yUUdrD4aEqToJxhOQJqpK7/Tq1k+Wi38bVZ2HZ2TEPi1qZSaiwxs
FvfY5YP5NNm+iU0RhECx1g9W6H+TykVRMSezpz1fYqL3vYmxFPPBzNDmEiTagAvB57/XGFB7mFd+
4k8mQQDycHB7HUjxWXkha2EZX8zM8qZ/s5HOIJdCJ10zRg9J3wmtCyIElNl1sRXVKH/6Z8hTyNLo
fP8Eepmfc1LIc/YFOarNQrlL/B2LLiD24rwdrj8qyrhmPQiCQxsGZjJqcFC8lqIB0UpVLb4po8eS
J35NgQCCNMH8IP2Vbu4TXrZUlWSa1W1jUKgmn4SuhfSLlCbRO8cgcm5mg2zYB+0demRYHVqgoHQs
QW/pRKelufqWqSjoC6M0w13LuYI8aMSwc/4jceutxh/4znbwlj+3JLPXhRqU17XgnbaQGL3lIsE0
nvVDu2/9VeODc9XiUbTEFLejDywmbnuF6NTBEEyhGtJJ4AJDpqYx7m+WNyaZXMrRqiALUjqax0/n
C+OIVxAZiDVnPOa3sihP8/yBM0F9Hl8QlJG0CjwAmSgV87cgz29aTTv+X82pauFFgMMkw2i8grni
aQbPiSqDACglN6ubImlZLOj1Kwy14yWJcU1vyUvO3IfP4zl0+ig15azBhUot1UFYOQendTwxXPGU
qm9kz6AQ6oE4MH9x24ftcvguc5f1NhKMmPNnOYGXLlWtJiawcM7aPFxg1dXEuyoAgdnTnaKkC8vd
TB1X1+dtzM88O6sm66QylZYJzttNAaRTm5+aIgiBztvzll//fhQg0cdDVEstYTNGblyCj+iV/07I
wN06SIAeZJGOGD7je0y0siWsLCGA7Uqz3oUS25prExhf1b+bs3RId1TMpcD5sXlmv9C9yRFnlnva
ju21q0HFOjFbAVi6t0+TbY5iDgJYMinVoTOJ7qKSmygQP9nuEUPtUAnllhkJcKdMG5QxnNsqYQpn
/tPSMdUxM7cvLV5WVy6r9IEHJJHF0YWjqxlF15nLyGmvhLN07Tj80A5pBEh5BLPGzrn8wRNr0Uor
c8w+LBzeCpkY2Qsfkn1fQxNAip6q7xaE2cNU3roINuYRfsba/uqO5vsK66i9PIEEFG99hZc4az8P
zTXhQSjs8UliyxQpJ2kheshhC0DFcj7IJhlkd8cpda9rHWcNrZENHKT++lQ6hH+DO7mAo0s9AeB6
jGKGqzx03mHHxP368TaptMgVX94Z8iV73bH0ZsJtj6/T+Viasvta/2yzpztWzIi9dmsxqbayiDzj
vPtsfZkaHbh/HOSPnHjI2JXhLvnK4ki1VapwMT/f1cUy/3pd65EAbrq7HVp4i7u2JA31ebhy7HKz
xBqmfuzuYrs4Jc0g9LKQaKxx3HzEhffKWeD2aVVO3Uq8EZGZsfSIxWkCAt4QXRIB8E8VxcPly32o
5fwNp+zBD92HYh5uTZx6JHEFmVXHz/5WLleQgZe2lmlxadkXtnczH8hzuceX91gnZDvOTN5JRjMj
wO9Pv21j6UeTyPsVuFOqobH2WsaZeVv1l+UlM0XiugTUPHO78M065FhujDFTenoDsBY0q15e4A5I
UF5PFr8mq8EgjP41WzKLfQV0kaNDRvRzObaP7MWKg6gZ7zU8BgjAuUTMpHFKTutQsSUvKKwaoYN3
+hD7pq/wfZad4jBTo+lZW4W9OSQk496ai0rjWc5c+tTCqydcezVdFqr4+fUHQpsdDa8ecemVHgET
iGEIUiIe3rSHG/9EbJobZ9a6UnWc6AY57bxCxd3VFF9RTl7l3MLFvRaT36FYy3T+Rb16DIVotCxz
b2r4JPIeWcsHtukL63iSgwiyKGt1u2o8tTqqg8XSKJqUg0TAheY57zrbik1AIgOZN39jSvMxiXe4
yvWXvKUnrT6EcNC0x2KvG0/iCFWZmmZrbMZcRcaTH7Vfw899aLZe1RuJMywnuEo+bRYAz32LO0Gp
AtK6t9DnyG1R5xzkD4pg6u4/A6knizwqs1EUIQiBf8O1PcrbGsOgoVUZhy2I52uXi3NXZu2xasod
ihPYCWyZ2wSbyuVohp6U+pyj+yNN0HWez38ACuXOmMeROxEkRYB909GvWqQbjt7YVM195hwAVGZ4
XjgR9Vrk1UKsYQ17WscXr9NL+rWsj8hJWkXZsT0XKs03dkkm+rHmj96hwMcaRXX/oKA0sVx6QSEB
+V148/QYhCPFOadpuUhozy3EMqLdMxTijbRS4nrsaSCT/UsJqRyDBzmwFtbv8kwW5BtEr997F345
jjgMhq/pzEHuzeuo9KCpjGIA4MYH/8y7a4qIQ1xE5RzwwIDA0Q5rhfVHipePlbxVRp9eLkqMiETT
VAVWeyR+25fDF+3feNw/wJpZdHNctAz37tJSyFOO/L95QCCJ1ImZLMBadE6CE1xLvjDRfdH4riBq
zxqVMT7bJLgLoWHof3tSUFDT+5BGwJxsnEQEqo+JTGF5YlpRTA8XuO+aV5+oP1RvM7eYk6Vzdlbo
v56Pt1iB3I0lYJsBUpHL/CkZUqCFHNRuyNu2VmDq2W6AEIg822bQqQOu2OTma8IroA6sceP8zuIk
Tc4RTvps11P1cLmB7yq69uU3HLXw6jzIpz8zNwnEm9VegaDBQG57wnJxSktKVhk+JEa0GiXFKYcp
KiqRCZzd0GFDgQ1ET4q2SMpAUDq0l/LydvCHRT2G8BIynD+2l9NcUo5TN4Kso83IucEH4F6yzLLy
AuCFauXTZVOLc//kAStzx7ixV08SIvnz87yq9rZJox5a087bbKuZtGr+jsI2rhNz5HD1lBgfk4om
WMIPQUL9XlIxNW7IfgXZcLZL+F0gGvVRewJskiaXMRnUaUS0Fg3pJ9fLOhSndEGf5h1Nhf2bw8BD
q/H/sjQpFHR2DPjgwp1I+7DKdJgSwfkY0MSxvIXKcPVP0cElK898AZlxCBk5ZXOEUCUsvX1T6AQm
NOtdMdBd3KB1wEMmyHiFaaGTT5fOtLdOs+WAjEsMECMzXQ9Beo88ktADc7z596kwr0UX6THaBwiJ
GS9a1Slipye3dHSUJAKTQYcJnybeJZnJTthEDOLJOqt9LLmU/iBWvAZ9GlsZLIVQFTUlBZeb9IrW
Z/oW9Vqiokerr8EzE0iAFacIK048PhIDMkws14l1HG8A4e4oJjOLPoORf7hzpjD7jmXGySRqhDtr
FU7vsq7WMZUhKHUYdkoqr93th79dpWWncZkXqAOr32TsjqZYrF1xvaAEQ6DNc0yCvqfJzkF6+qki
wXUJuScKGLy1TfaV2/kwTdq62vkFhMXpYh88rpxOlZIsz/5mSzDqFvrc/nS3Sw/RyrWQGN7rV3Ow
o5s09ODPvG/TQa2EUcljnWgS5pR5LXfPxRlUW3ecS1vfUIbbOTSw6IBMFEAOXIN3bluBJHe+nLCt
MaRV9nAAL97w5JFAtMJU8CCq7bmksHcaXSPG77CZPpuoVrTtmW6usPD4VGoTYSjDcCqjjM0VaeUj
tvNL+q8MKh8DrVMz+Fq1TCPgaAuav02SlYL1IIP6JbVpaGRVfhAV4Iu39xXhYDh0Z6vBVJ/2O9QP
ILMdRWmqA5vxHef6R/L4+IjwZUtjLVB+ZoCJ3ZHva7q5WRPWljmuXwbcssdD8/QOqkWj+lMi+YOC
SjvGT8893MXaX8aPbCc+L7VLDTkG/IoyYsIv9uUnyeTGCd9lbJV+bj3byGDS1WkHtTADvnM4Z1K6
JzPxeGatKrkedKN7JBhMitI44QJxyGOGJcvcWS3tZewWvEOe9BJbXbXobO9KwMFKqpUkVcAFpWku
SybZ3H7FHdNypsieWP7jdZ0+m7dPYy++epoB50mF6panlVGR3hT+CiPPPtx8y2FPHH3ufWRk7h82
uEo/1/Hq4Avy3oWfOEJd7TkiHZBf/fmoiGl/AoCiGM7KiD44tZT7/pUFtsCBK0kq9LdpXsL84SDU
fskYAcXJUkYIgclBWZ6jG0WWuMztA0pZdlc1zeAdirmWv1gyUmUCgm2oJRMIfW0y5KiSWuQBCuXq
3SvnjA6k+cf1nnghEB9ZhTJjr2TGk03Oon7wgy97/z4UrMW4JeDbMyVwEzXPZhCkCcyl8vKKs/At
aVGKcjnLPMyehKvbarWiwAcwAm4sGo02MCHcLsKzgIDml9joFVpy5IGKreGqNO6yyZzQZzsHhkoG
Qb8wsgzXkamlsgYZqc5zsJt89bd4CtA6hsqzQWV49sIYmSUAK7cyibQ87PxWaMu8UQb3zEZTKuB4
0Jh2de6C6CTX6RIDlhBkyJhKp6ow8MWPg26i7s5mCROHmn/DlaVA7cLElKPYBpznfPHtYGnd0wKa
dVE6r04s7oZjgndd6VVeuxC5Okh2hZ3yWGavBCPPhedWrbcV5KcHOBOyO9R1+VI7BLLdTPsqkN9m
txSB5ndsog9GRj01LejF9hmTi+zcx3KXyjxCdcWUxiGl4+NTgZCmpRXlbRLBbCzICJvjLn133/FT
N99Px1qpnFxhYvY49XoPeqxSDZUMyjc0z3bQ0rhpWqaeu81Qu4gLkvlgBbnvHEX8PQ1INB7t1rr5
PGC24/+Ct8jxwGMddoZkZjLBblczGkaMg4h122PXAVIzG3AJYXVWs2e/82E+VX05q+WwrQrA6YVa
X8/g1KY4acoYSYYaD1jh9w3kFovUQrfsIxq0FMolzEomgJH//d005ZOyaSEQoExh/B7hXaxq01fQ
Sq+6OY/7RyXYQ11KNS2j4x0oZ8JoMk/nWcUtB8AfxDPj3H4FnZwxCocfl3PvjAv8RRrVY+XXepOp
ac05XL9niWWVCQRVEEGXl5tr6S4NVwmitBnwuJN7zmzljPcrJBzwSUBXqqxyp0bG5srVxnffAdWt
87uRqv3ioy+lFHeEEvNHPu/fMfkAIqMPMPZV5HGdfzscA2b51NdM5gQuSvjMLnxC803pNi3zWVF8
MVcCwt75fOXTMyxBGGHi+IEk1+8G6sQz0lO6GzJZKZz56Xw88rXbvbKcJ621olSH7g0g+sAX/Yt9
Z7RCff6sNkon21zXk7LNl1g1OUUmsL871tb6Dr2HHyfNyarDWFxpXJ/0YviKryhD46Y/Gfs8Zu/2
HENylHorP7y1lPpzykej+rPKFYPcehnSRTWpi7oaK+Y4NZ3/xNnvPUnCyXDEcbYSJJsaRf1DmOIJ
RY9hxILTEXuIedZUOYdmIEGnYCEuu5eCagOCZ3t3xMR9lRQ7Zml9FRJ0hfh/n8napzNijfwXofUI
5rVp/KU2LttyqwnMeSQt8pkzwAlqwAHQg6D6Ub8mWRrUlrK9ya9W/GRzhLVdtc7YIlw+PjE7SRNy
KGFjBXgqFpstxmg3IN+Y15Fwxu1kR/SLElT4aR6t8d4fqxfEHscrC94v/DJn8Lmn4+jyu33JdC9r
3odB+7opadLAsRdM4kjvU4/1JUNKPtAyHqPj4UoMh4x3pvhWWfeQAnRroBwj/eDIqWQ8VD7cPhpE
dRBoa4bdrSXOHRazb2qh66Wce/SQJ8P6C5IRxg1qRDfiZhqBqLB5MMNGtcbWHvHpt54HIxdeXWIA
4yH8Zk9d1T0lHLCvjIkMsLeo04RDuiTxd4OEDZS5+DO9aJghXk93stTKWklfStDeinVPU4jbTiyN
J7zOXnAaSIrgF1y/laL4FWeKBVYPxq5MN3hAT3U9KIr8a2oihu5Vdg9g6XIuNUivkTkOHSnwsskJ
2oC2bxJpjjwR/mGGcNO8/5x9cPaVbXLliygHFIcmvdK13PtyCJyS1M+PNkUrVjERZ1pKHJwEveIf
DC+fY5PX3zyG6WklxqKugHux7+PSuESMFHxsEcZTZyVV6bCoLQeZo/MX5ED/dNDHVXjzbycIkap/
kZ79COoYRtvyV+Dx6Q4PMrYLNtpbqrwpWPbBnAG9+ukLHQWcF4b4OYVkNxmsspg1E7efhNJ52NCj
Tw26rwuHPcVMXMG32DPd09RIA8j1vRQLAm/tgSziRElMWHx/lYc/yP8IRVg38tEb7QySxabacl1E
9dzFUYMjEj0GYTgOILiOL4fqTN3N9SRbfuAFt0LYrcA1lgyCG84hcmq7UfgpW1bp5mW5Iy4yuTtc
izCW0L+Zo7+QPwczADUa07Gb/9UjJu/FD15eqiJz6L5R/nR3bNvHLzHg6Hjyb+STK/frgnIEJyu7
rTFW0kn1PMsF22X2Gew04LxOy/kHrIPktH0KMO6Q4TA27/bq3PDwkxnI9NXVfCzgQkFqX0kZxeFs
F4MUMm3g7HjdO9yw3pkwPCkbBqfJPRt6aGxooGNIJlPysXnuPnFuBf2QCzNgfQcuw4bpEM+ika04
9WeMRjT2PC1fx+bVQ6lwzzcqWiy4nL1OI3LaX6RB/DGPUOwJcs0lUafsL58EpmEo53iDQlfqw1zM
aVIcK3Cgp7ubJbMkTnnL1vy5+VeRtWNPmuL4DlOxYCsOsmwIkJxHxK7UdujldsztjyPz0UpZufDu
K5SCFgidSLfmKKGzKRLGihOs9NgqGRMIikWDMm95xmaiLVCkzzC/7To88RcB3E4CGueMlY5zFMDa
jQP7Y1opSo0t/iXeuVS369hS/cRN4/DPvn29GZLiZwKIyGD33jbQHYLqPG0RM1ClwDSRsglGUFgk
a7cyl1WUxBr2D3aTPJPMQQs0ISMAgwyfayG/EOokktNWIZJVLX2lQ35L8H6lsE7nziwuH4BrD8j+
Qd3xk+GHJ55chqTbjZXazeXiUryMGtZ+3ZM+Hj6dmdjiBBROULGDLSFpdY8diSwM123AZiElDf3r
+wDRuZYykeSLyZJbqFKUzdnPAVZI39m/Bzo/dZfrN00TCddqetYZ/fzCJ1gcZB0ZpAVX82c+vw+N
mBKpUv1KygwNdpasaU6CyAFMjKMCdW6wkUK9Tir9yoUzAsHMBy8/4CT2DKR5ZNPU3XkMmq2qgfGT
V4OGucjgmeDjR+I4ale1QdZ42KF89i0/BUecaA1P4CQwT9i454Ti3k7n+cnxPXkoVf6MfYk7879X
0bAfYy6+nDq+GqAsn3iCd2HCucKG9rTmzpNNK+qWTTUXT47L464GiBDpYCha1UyvBJYdQmyV4hia
sgf8Xv3hEeATCxBZtIGeDMrusgGsuqfiRzxdhWUIgYCCblEVZc5lgMSyPb2RhUzsMkHiUH3zk3u3
J12GwYkcVpyRDRbSAtYCHMajS3oHIP9RiJ7667qECDaoLuds3OQtsvLh7WH7c3zpG23ejlklFo0f
MdtBbpckOhPWrh4XPbkS2BjGh+X1NW7klQhDmkmYbdMCzoDoNZFcA4svJhyP5nsxc8dvMRJ9SzQE
StU4t0vStD5sbUPvM/OtINq19UQIKaeZjjLSg8XHZ5lA1j8zynowGf7mE/6DHT19VBDsycDpeeHU
wGf+3ODTcHJr3tZ0nyC3yDBt9bk172GvNbFW/fQ4S9cS5W98Dpfxp3ZWt7uuoMFpbslQVjCv/AtE
VfGTqnakPudu17a37kKRQ1Xco91qbPjy28kWSjDzmJeRmNoa9lsITU+SkxldnmzCUUekCwItFsyL
tHQdBN/VKDy6vqOMyIddUuqP75s684o4kSSiaOzuVrGXG4y5ftcjbZUw9ucAMVoXnsqaNXhweKmu
+nsI5kIUI0nQ4LwQBgoCkzqVWHHJplgG0ZSK83p2IPfBTD+z09rAWA+2Tz0EfIoW5w78FEWZNBae
YWCybvsycxgfSfIAVDa4gSPsEeAs57hms/Fv1luk1GOTd+Skr5ZhOEP3IwSIfGgGnH1Vc7UcCsyD
d6VnoNEVIMax41nQE+uEUHJHu2YjMxUWSxoCPqsaaxKteo7qJrojXP0rUSCfmnDCtj8xmoVWlqdf
V1KlgUWfaZCrFvfNifqrCaJTgjsz0+KxAezKhBGbMUOn8pLKytzTkqKqLACZqiLIGHZ7ZWXwNLaU
067jkICZ5F5tziQqBMFAR4dn5sZfQDDAfYPFxNblddHLForaYcLpFpGw+X7u9ssYjiZ5/aw2XX+0
f+aWlclZd3LVux1cwrN76Tbt7l0/Q7aA0FIiRqZtWYoTBUq+jUkkWrIiHcg1XWTEm0WH+gnwxvbU
DDhSFQsBOSOfqdflbDbaFkEM/MLXxF2ns6ARVMrxLBqhxbAixOZYuCpVWFFPu7/8jHDtDxfpOPvt
vW7W++qScaYUVtf0lMKz+h4//h0YjZwcOSIdqymw57Otv9uuRX83nQM5qsQvQw6XqFhgUL9Vls26
Pe3dvKIapQ4tn2EebToQOH/6pVmOcfbw7AepXqz6h3oJTarpkZSQR9XeDqsR+O4kddhbL2Y0I0lY
P4/KhKUHx22SLNA9qz+9LWg58xRyRR/17m3bE5wZGizbbchCxXHHDZDC6qH1XJDfaESjTWcXG4Aw
YjLFW6lImT8YaxHIjfmgBGub1dE/6jZsDyLtthD33qaBfnxMoqYPFyzJuCoet7cdLPRfdoySCQus
Lwm3TK//ejNrM+fxT1BgrMmYBju1xSFaCOrKKqxFoVzJY4X5sGQk64EFxMePbYrc1EIkD2eE8wb3
Lrq5lo9VmDh769l13Gu3qevwttb3BS3gOYByBTo7EP/ba7VZDu2AQYY9zsMwt/AWTvnGoKoQOk9/
nU+bzjSHPUnlP7Vgx58/TzIFYtwUGbeZgLAVhhfmqksexjQohyz3K6oZFmxyLCzgzQPBB+1kdnOa
ew3yXpbhzzjqTZp8aOLk4Yaim5FgGT7JmkI5ykZIP2sxPn5x3E7aLnS3yznKDSt66Zt7UvRAKfvz
uoj0O2M7Qf1FzwI2bTUpYM2ZuEKD5zLMSD81Q8jG1hpLuxkGLJa416Hg7a9cCRWHs7DhixZ/6LbE
dC1KU1GoKSkcWrBsw9+CuEWNc8IAhEaKLQ1Y5OMsOZdp5F7vrJ2rL9tJsKyDx/S6mPBtWY8m/6bp
drFb+DLi9L4WUcg1qZEZEkzx74tiiO+nQeGg1dMYYKeZ/PAgfm4K0lEUyH5kL4jD7DZq1P2XU0bK
S3KAk9ebcq3ASWsceooLgguvBiCCOUK6pC8yfbp0Q3Ot1MH6TO6HVvOrZePMScfMYwio/7AvGqWL
hyUVcujDpGWZFGCnrSCgSyskq3tWFAc4lM+xreZL4OOd3f68hefbfXfoxsoW6H04lhnoKHc0tUu5
HGgQt8pgUc08L0TCJRwOKm7KAIu3o51KnlniyCKI508eJnAyrospCUan4tIGRUCIn3c/wKCw0PtA
2Xu6yME55mqCZfEG2y1TpOOgyt9h+JTdthodATbY2lONSUngpmwF2Kv4KV1ZJoEBWkGGi2FtYHu9
J/Lk17T92oZdpNLTIa9jiIIwJe5nqjLeIAvrKHS9+poSbNlY1uEYz1E+ntIg4XSt550W2J7FNxIi
sY3hm+5yNafebKMrz0xsvJgTIvCvre+s4OE7nGAyaIh0JzZiAUH0BmIEk7aHQHWptUYUfKCT6euE
yjP1m1XRaLQe2TLzmPR4i4iMaI8gBxYivRq/Z+WRcO+9X0Gv1VV4qU48eICfiTkDRdlDCu+NVSSY
DmUv0POAClZAryZr2Viv4Bgj8Cii+ahfgVlv79xkPmdHzFfWeuhxEEzM5nx2BT1CX625z4NMFRNJ
G3oOxEoeAQo3YG3FoXR3GoNHAz7FTs6ZjKYaKvLw9FSt7Cw7RD5niumMLvRw6iQFt/2tsck6X6Zx
YEWSVhBpLNW/phbiJ4dpVNJLJ7Ic+xUFmcL7U1smZtV8qTm8FfboMYNmekneSs/aYfgaUbJ53RXV
+dzDcpfiXmaPKYn4alwCG9hRDekh6DJrHelm1yFDnFXqE7lXdEyKNDuZEHMehZ8FBIjJA9Edn/nK
3oGPwVrL6lry1aTri7UWMYHfre1tYlKutmW4YUUj4aY5u0p66moUHbwybHANnDJrW28BXVyG0eig
2/1Ki6j0dXxEJDJDTJOYwD7+1qbPhNNv+PIRqvvwj/Hbn2XWFhku7deVvRStzLqc+Kimf464AW6r
QJ7b3DNAl08BKeG2PENqvK5CClJ4vwels2kI94KpKzrAqVRAPh5za7W5Z36DpzvZ/xOlHdkZGfHw
1w6EawVluQzIcM+VlowxZ8Eg2qxFjjh1QmeU8Vr74wuVT8nNLZxdby3ywOuDK7JxPW23+9hL8aYI
Zi28Tpq/3Q1pv3XUODNmyx6MBnxJwuTHaJ+Y1UYjRCADZbuD157a1sC6fZZzeRFBxoa0voNHytEa
zx694HdU1kBhKw2Qe7Z+tW26s3qgdVsMRwPW1TUVVyQXynpPOe0cEEdjqM+YiejjrElWji7KUybi
M89IABBTe/f5TUe9ncZMZtGKds5LYHch3XBOXzyF/VUu3pHLkAeTvv+twVfbo2XirWW8R2mChIp5
miJFJNWqxQFijK9EM8fmf24jcDUebBWBOzpIhy91dOURxNuRY9G7/nJlgGJ+ORQeJJECIEJ+GGOY
A2/4szpp9eMSd5ik/OZKzrWzaeM0CXlPmiwLTIAI8yAAJBxogtiQ2/fBH+Bw9CtRZGi/9hcdprLn
0QOlF26M7st9G3u2IlZZBAbi/2dfNGRoVy+b+cBhES4tVVPzf1bX5X6YMYSIuticLlYyQCWkOOaa
2nUt8OzbGNmjF5wAok3W6wODzspUGR7KhE7vDMSOyzMAghjAIH5s8iCxeNE9rb0MQF1QqKPP2Ngd
56Isa8XkwlDQwpGRZGuI+BB+sDVWGHaTDnoo79knzwaUFsr4/zdU6oWFMsOZuaf5llsgG4xalS4O
W5A9jgPn8hPMU0h/eF+p59QF7Q8y87mxxoJQbIekViT37/B38HxaVt1espiJRC2ErmTrN58vtney
KN/uKRnt/SzgaF/PkJnpN6SKpYOTxGNKuMiXwsxDnmkl0bMKULGx1OhSXPy1XG+aFrG4McrqEey5
S3YSoNH1ihPdyVh/L+h5v3qDLfThcNwBVHM5ow6pzAljeaEpzFtdAw54drmmXqothPw6CAMBdHmZ
RAa/cSU1P8pooWw5qJPxCtUqI2aC6opzMI12pwJuGrxHa/UQT+FaVsC+wEQqzDXQIxDilqROorDi
wczXCDhi+qeCGxocysjJq3pIuY1zfVUlP8ecQpc9uNYycPWv/iGpjlVeUDdSPiy6T88x0AUVRNhV
g0E0qDgYuyCVeQ3sigNmRKrAynuL+lPWBHrSKvPwLJL1TVVefadGA5Q/yxI0PCT1b87YcNjhLWEy
ht1uweAIL3OECqCxyDi8wrkvKIIM3Ep07pcUjXFHgINXk0So/e09LnFeGRJ86fbUIhfDL0QQHX4X
8u/LT1uOAMALbkOJmuB6tSrA1VC3pqBS9ZERzjGVuJNqXo9r98NrLpQGssdXH45K24txGs/hNIi3
ait/i7EAPY656g1M2KWLeIgw4dUOTyF0XANETaNCwWFC4pUCuWzPUgAM7gJo4XXrZM5EmX9c+RaN
sW1ZVyohyUB8qpufkLgAYrEGoh95cs/woCW5Liry+2wWekCVOUHb/4TDcYgQhuzMjrnPn4Xjeb0/
UPZUzhDo0WZV04wfmDTvoor840C/OoaLSckfKNRasUweuoh8+dbL5dONH1LHKu595cuvOG0Ld6OZ
H/BCdy3xv7H9+FfwumkmZj6vexX2ZpnU0zFOcMcLpkcXsGRw2gu/Kg6nu9BlfOaGj8LYUwkZ1lxB
wc4L75yUTE/tYxzyTUIXEDZwWm5IbQs7HeVUq7adRzWYD4sUa65BJGzInvygtj0OjRmyUhCJ7MIp
Dx9oW2MWF9lfcA0S4WIdxW/M1wrHnm2/gsqB0MUq82ygT4jkVr8KE6pKbPnL32e2rvhuV6iUGVEg
VS3Qgw5HybKGS8hOqpbLIVsj4Fx2nomnUJGueIgAejr38/e9sG0eTfnUyxYpXRHUoEpAV4Tl1ABg
YfnEH2EVnr39jK3/BBJu1+PjQ+/cXeMHVF8bwod0hwDMoPOFzz2Rzyv+8d7b969u4zlKMK4DXKTl
J2HkeBBuxSgHisgshVIvyRrMX5J3Am52w1GFkzzoqA==
`pragma protect end_protected
