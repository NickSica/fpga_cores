`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
iQbEix3JHZTwa1vhipHlmwS1/G9xw/soq5c1aH9r1Ikmd5PFC6vG8hcczrO5Gm238/UZKbDRHhQl
8vxxX1eWXA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NYO2r/VW0Uk9iILO9avt3Skw+TFdXKrXeDrkjkY6MrmMZXqmt1ljuTdXla3Px6GiDC5iNRfSB1LJ
jlz9x6ZyMo5VxrDlXmNLima4xlcLjwQ5Ldngl558uz/vr1FbORoJ+gk4f03PWwyf42EKOYFnCVfd
LJfFRdBml66XWTkIRRs=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hXM/negBdYIePK99VNL4dA9qZWSDCbIcZGIF+wzwJF2GeTdZiC6Sv8N9/cF1YoJ4PmeE+1cpGoYE
hr+rxDAb1wjgZvfDyEG1QWzKRSG5E+oNC6Bj2Xk8erPPxuHL0sXJnNFmZt3mRdMMjzJ/oBGkUF0h
iYE6DHIS9BMznThGr4tm6wOQ24nLfv2CkGw5FtsfpBEceglyVNwc5KmDZpqUutO1UmcXWgUVf6aG
3t7duiHDJKzCaRYGI47UkrEGgYTLtr4N4clyKbc4ZaAFsMfafXuq7UodHyHPGa7sQYA60+7yMSq7
lZ6oowJsQLQdpXSegbc7gK8ezWVXMGToMCUX4g==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
IZkumnZp/JsuGCxK7A5f04eL3wOhVC/HIkiq9ThWDUN6/jAV9gkhdECfPCdAYxhe0IfGI1mwNrRJ
CATeVriO+TbtGJF8trisSNtrtJxyu7w+ARrQ3i7xJ5OugSeDn5jrGtPVCeIVbs8Otz0RthJD/ia+
zMRiRhN8wPr8+wtwChbS7LbmoKzd361OLqaC8TX6Ab1GBUHFOMfYyAPJdl/jXbS9u43VHuRY6Yc6
WqrfDJE3842973TEArl3DaaLzZwM28WBp6JNk4Z1zR+7/fPjneoZl3Dvksdx4ThM0a5s9BNPAH9V
WF7gF4b9Me6TfP8DfbNOy0URIYx+xbfpe++9uQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eaRvVH2iXg+bRFhfU/Zdu0OhZxAtLuP0NVIWmdEUooi3G/jC4AtcmpPrp7p/DrHH2FZwIvu+AbK3
sY3ybtP3ICKGUwlnIt7XryFabcZX+wxEJ33rwyvMH3qSJUvv0NnXC8IHlKKyRjDylY/oANDzbz6D
+mWDv16FdHx/0RgRk2HTfCPx8qBZ+fT4hbE6exCfOH2KzbFjubsbEmNkNU+HUDcusYXP2EoAnNGO
lFufKr3GhljOMYxxaVeKpXEcKWjQB5Uu1M3JdONHHSUP3iVPekneDcajTRMfHD9FJggiLA6mAgel
cdhHqUxScYsWsL7cenQphjXngVDIxqnSMZgGGg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
heQDXwsWtguDyBBqy+N/Xr88McxL4tQSR2XBCb/lxs8IKaambMExKMCiF+uYl01VHmTIU2W66UkM
7t9z8H1Gdw289KkEy+LLNQNFvy4xiQp3che0cCrsbm5/JjwMeuGavzmF6wwMkz5sW4oMgRBAsxzn
RRGXDS1r2TiNXhNi68I=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WZqwWujfHGXV7wBEePMjGLVWUeV/ygCmf158CXpAhJC77z2vuuagSDsOpGgtqyakG2cswti5bhBy
iGqPgNkEY7Q4T3NMe5WssA5nf18Sw3LU1MCehsK5WrHeKiMOyz9QpdgScXEE86/e3qniqvFlM2/c
HpI+I2e/HN1QOgChXb7HzAEEqCCdY9VD1a+p15IoOmU/8Gs718QdaPMJOt3XdTu5pAmq/PWuICaZ
VFSPDj57xVELte/pDBIXo8hgI5sad9ci34UyXovDzhRyUKzLY0u+gqRalObdZFD1Ph6hGQiLfmwO
JTvUCIjoFwTzhh0dCXYGcwc8O9kaaOIiiwpgyg==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
B4GVIi6TGeAAKF2mV42cg9jGmUkeJ9TkEGN3HtEus1MF1Zmt7Nh1Y005XEEzr57ufgLlM872beae
bxX2U/dQHyW4OCP8KBTn49Kmkdu8j6t5b8W5HRsXXHYSGPOo9IxUSHBdhwxHpNWauRDmTFNl2lia
Ton0toY2wVDxIcyINRYIpxD8YGHOnHSHPMsgAGtuP7kRvUnSvNzqqhzVcNm3oeIMTawuhFgBXD+f
0S45sDt4HAERXJfO2RXmlDCCLpg7FQxibRHwoppbdhT48SpFRar2SU9FLaP1Rhu4f8UN/BXG8JDH
IE70hcE1uVmlqXL3h64Aaql7Kf0Mt19/bANOBQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2480)
`pragma protect data_block
8fgGNC4HfskTXIPOSZDcR6dwMGdMbTtu/lw4gVjAq5h3bL7NAq3IdqfiWFu7+ci13CNpcvSGoQrn
TyoLiue4wNrmKn2N1jZCUEOft6hN6l3PWjD9Pjv3vWsDH7iINrF8kxrX0AdayWDdqJCRI1Tf6w6y
xMGaMyEntvUZdwwJ1sIc3+TXp/eld1rmEEA+/zmrnA5L7ycxXf2+RE8ewGkQLDAxo283HUKK7py1
o4wWHJiFx0VLdfeetIMKq9tNAz2ZDBz4GQSkD5VlAQrDKPym4IXSYasR2IN2S5RPpq1E8WlEDKxT
QT+8aVRKFK/HaJI7CTNGjECHtX+dThZpSjOQA78xsNk1jYmwdiyQSwFfq7ReGj11A/+d1Y8ZQp8b
uL74VlSatjktAoHnRfJm+46CEkK1FwBsL7bEVI3eIe6wemEDr+bEal4v4py2vgXYP+6wavIz42dV
kjqdnpNNH+Nk+Y6flIgNmFoXDR+iBHBq2Kwd4WrZFykxxilMih8lUKresceEU3f1iK4gdLbtMFpF
ZeneN6wDYn2BRZWJK6DKScrUQQg6zwVuQD3pqwkZupIAJKlMHkUbQpR/l2XZSBWeBafW2li8Z/N1
VvKjQOlMHVPyCiT1pG54ohDJXajSjrXL/v82JqpmgTZmiqjTIEimoPsSAifIrovfVKDeeQM6KHBx
1IMcJzxesfYyLvYOkHBmGVtGohob1+KZ/qhncRuDHUt8RvOZFlgvbyCeGVvBxK9ALnR1N0yFtxTw
+RHHA0Vy5+I5yvI19VCXiO+TjiypRhHYvyiVTO60YIbtb0D2M4YQGzRnmR6WM7PJYr3dfyvs3yvT
7Vj1OYTNHxBYtn7CNSH2sDGNCEIAH+D95qEuNYJ4QcelOv/MY+nUnVP1dp+fU+WNI7Gy6LwO7d6T
/OL7rLDBx+3VP2VqUR7P2yGxjF3xpu0o9D9Ssi9BAbFoz44uLhVlIUR5ClMLSNUjVKhIx7nFZAIB
7E7z+YYYXoX0TGF2Z5jTLbA94TgnSpy6ETYpYDrGQ69W2xSex/4FSVcEUhLJYP/xgFbL5771SXS7
0GZCFrJBKRSlajYLpoEYlq3FrFKAOu5gI7lXZya84mavTm8ItU60YcnhUN+ElvGRhEk7ROB2eIrb
8cQLOZw1hlj73SqHjFLQmP9QrL4TV6Dr6UX2sXq63meKqxACaAXdq01QrB8nrml5xvoxlf/2rrfV
gPgLhZErd2lnjz7+Wj3N4Y5EffWKK7hvCMNBVoSiQcXBT3xf4nCdT4NbEgih+XOkhZUdBC/3DbGm
nnZjOzHUswpm75t5XGv+0fxtxPRSWR+jyYCpANvl5JXDooUnhasXamdUK08uRAN0HUQx53f2taNA
f1V9moOYdPu3kmoyBBgo925LGGZ2r6wxpKgwjLoC6hzfaNcbveMLy74Fdq3NnCs7ZMeT4qdwP+fs
Ud02q0B4ss5ToIXAR5VPlTICF5s3QYE/Kqz79ydUeBnraK7MRoI4avzQDp4OsMeKbVlHtZ/vf6RO
w+xYsDRDAgmZKGvErz3O68hWxygAv+Nft8XPLSuWwP1lcLUlnm7TqeGN2+RjZuPJelgE41OzEYrm
jXxoNozDRrVtb8W+0YUbkFJ9ZE9J19oeNfBLyiG7LTc9nmHpM4cAph6nB8t+1yJ5MnjG7CeR3Y6O
+EyVdCGP5gm4nx/etPkF9hD2FaAcq2ylYpzhHcG3S9/AcOg9ezErNVYjzvFuySrDoMOCp/MuvPUN
d5IYtu8rmq5vAQKlTua1SR9/RMzd8SSrS8ocy7T/bg06tVxzsbbV/7wBcS9j80lFIXWCDsSxp8wk
LfC6KKQdKm2g0dOueKIKiux1hKdwwqsKQEGurwnhwt7bfIZMZ/g8e5IH3r8yVYjt+V80w05UG5xm
HA+bwYGJHsYvKOaCyVF72lHQzT5Sz7eBLmjqqvk+TacCoNr0wcEjjHeQagIjOPN2nPC17qPYqt+R
2fGUqoRLVkt4njn6eil69GwAYs7sf7+13IIwgCI41255SDOaICaY3yvddFUHjbqfYQnYwUZYR7Bo
p9/PK15obcl4SIBUhWpMVyVUou7Uj3mjSBZElPHmwz1b26h6GYidDcoB+MWV3VY2GUy3dlAsDXW+
rq3Fy3reGEHsgtg4s1BLVbjlKibPrULPdXJ95SAWS4Ux11JuQcQKivlUBAj0HrC1f37KIptjAALv
czOlTZmJH0ogpR2LAHH5VQqyQPx5LZRda6aNxk6eOvdo8pKjB5teffbte7x30NLaUC3EMxJLm+T2
fBpJwll459BbH8ONxYIeuR+eIQ23K0Y7TDFBBri+j/3sVjadvLnGTOLLuwrZIt1/hwZhtE1jTUY5
1sYT5eMzL8wE53FFXKqGE9EVtCXCFvJTGN50LKDNWzQTZsN7bFjQbwEEiUx1+Mal6a1gAIP1Ejvl
3e6nHAtmcu0DA/FJ0HcgPwu43/mlGQ+Aat+AFqNTWMa3hcm3ZG8Mzx6GiWu5wMuTCkY8tJtHJWGw
oEVQqhuySrxYQJwW2QzbypB76vfhazac+8wOuMf6UEcnwakkmk30eBvaWS57kuOcD7cI5iJGZdO6
Dc4IbnpanP6s0RKsU5wzEIhid/lIlY9iadRo/fD0zBkUCzJsaiMRTgaDK2JGCKTMry2rhA3V+kg1
pKf/tyGydCvRsIrDOZ9Uf0zDYFQ1xeTgIuIQRmXcR4GoCqki9fVJYVUh55dok4xPwo9vk8NUD9Cm
KJCutOMiAtnLjVYiLX7sfnUx+q85mfmQiFwjXnylqwAmw/1/NWJcUM70IsZgIcjbkkwPHiV8LjSA
CWUEDBlbKdoH4nNR7AtinLhBRorins57CiYIW0eGOY7u4KH+LQYWqVriitblBAS3+GvXEHTjkQ/u
bsh0zbC0lkBHYwwC91dBBSdp2nUY9ZyKP15CX0Cz05KYRw8vSNsTMx4hwczeZq3nK/SCFcEDJKxu
1DgI1ZIbfMO5NbOvMtvK/xl0kBQ7M3hGxJhlJU+jOnHzJEl/3NZboboZmhuMNvVol0QjdizqOVdY
8iluENuLjESw1TZmYVnnjfOZFfyRn1it5R3F+/rlh3FMfwKxaU9tpgw1J1zMYiR7miV0rhW7/Aro
E1YcUFcCbcMxT2oCqqB0lefANAJu96nWZaMlXfAeet7EtGjL7hTd+oYbC4zctmsLFuSMaZ9K/cQR
0c0R1eIqaKVoBaWRkh2fKpDtdLAHN4T74rpcqvQTY9tEo7gPbXsLx6gxoX4+nCeAHv2frRn/8v//
bTM8hW0XsgCOgsHenmcaLvGqAl21cGAsHXMsV2c=
`pragma protect end_protected
