    .INIT_00(256'h022bfc2052220778022bfc204fe2200a022bfc204d8205a0022bfc00cf020572),
    .INIT_01(256'h022bfc01c002b04f022bfc2050a2b80f022bfc205002b40f022bfc205342b20f),
    .INIT_02(256'h022bfc204d82d010022bfc11c01010e0022bfc14c002b10f022bfc0d5042b08f),
    .INIT_03(256'h022bfc205422f032022bfc2054401001022bfc250002d010022bfc204fe0101c),
    .INIT_04(256'h022bfc09c0c20500022bfc2b03c20504022bfc2b80c20524022bfc205002058e),
    .INIT_05(256'h022bfc204d8204fe022bfc09c0c20532022bfc2b02c2053a022bfc204d82200a),
    .INIT_06(256'h022bfc2b00c2051e022bfc204d820522022bfc09c0c2052e022bfc2b01c25000),
    .INIT_07(256'h022bfc250002052e022bfc204fe25000022bfc204d820500022bfc09c0c2053c),
    .INIT_08(256'h022bfc2054c20500022bfc2054c20544022bfc2054c2052e022bfc2054c20538),
    .INIT_09(256'h022bfc2054c20520022bfc2054c20524022bfc2054c20540022bfc2054c25000),
    .INIT_0A(256'h022bfc3663020528022bfc1d00025000022bfc0b03220500022bfc2500020532),
    .INIT_0B(256'h022bfc204fe0300f022bfc2054009001022bfc2053a20500022bfc2052220542),
    .INIT_0C(256'h022bfc2051e2051e022bfc2053425000022bfc20522204fe022bfc25000204d7),
    .INIT_0D(256'h022bfc1d00003008022bfc0b03209002022bfc2500020500022bfc204fe20528),
    .INIT_0E(256'h022bfc20524204d7022bfc205381400e022bfc205261400e022bfc3663d1400e),
    .INIT_0F(256'h022bfc2052201100022bfc20526010c0022bfc2500025000022bfc204fe204fe),
    .INIT_10(256'h022bfc2053c01d00022bfc2060e01e02022bfc204fe01f00022bfc20522207d0),
    .INIT_11(256'h022bfc1410601000022bfc0b11325000022bfc20500207fe022bfc2051e01c00),
    .INIT_12(256'h022bfc0b00f01e00022bfc1410601f00022bfc14106207d0022bfc1410601103),
    .INIT_13(256'h022bfc204d725000022bfc0b00e207fe022bfc204d701c00022bfc0401001d00),
    .INIT_14(256'h022bfc204d701f00022bfc0b00c207d0022bfc204d701100022bfc0b00d010c0),
    .INIT_15(256'h022bfc20500207fe022bfc2051e01c00022bfc2053401d01022bfc204fe01e00),
    .INIT_16(256'h022bfc14106207d0022bfc0b11301100022bfc204d7010a0022bfc0100025000),
    .INIT_17(256'h022bfc204d701c00022bfc0401001d00022bfc0b01201e00022bfc1410601f00),
    .INIT_18(256'h022bfc204d703f81022bfc0b010207ee022bfc204d725000022bfc0b011207fe),
    .INIT_19(256'h022bfc1dcff05f00022bfc0bc1703c3f022bfc2500003d7c022bfc204fe03e3c),
    .INIT_1A(256'h022bfc346aa207fe022bfc1dcff05c00022bfc0bc1605d02022bfc346a405e40),
    .INIT_1B(256'h022bfc0bc1803e7f022bfc346a403fff022bfc1dcff207ee022bfc0bc1925000),
    .INIT_1C(256'h022bfc1dcff05e80022bfc0bc1b05f00022bfc346aa03cff022bfc1dcff03dfd),
    .INIT_1D(256'h022bfc346aa25000022bfc1dcff207fe022bfc0bc1a05c00022bfc346a405d00),
    .INIT_1E(256'h022bfc0bc1c25000022bfc346a4207d0022bfc1dcff01101022bfc0bc1d010c0),
    .INIT_1F(256'h022bfc0bd2003dfe022bfc2500003eff022bfc346aa03fff022bfc1dcff207ee),
    .INIT_20(256'h022bfc206a4206bc022bfc0bc1725000022bfc32688207fe022bfc1dd0003cff),
    .INIT_21(256'h022bfc206b62027c022bfc0bc2001100022bfc206b001010022bfc0bc1620278),
    .INIT_22(256'h022bfc0bc1925000022bfc32691207e7022bfc1dd0001010022bfc0bd2101100),
    .INIT_23(256'h022bfc0bc2101100022bfc206b001014022bfc0bc1820278022bfc206a4207b2),
    .INIT_24(256'h022bfc3269a207e7022bfc1dd0001014022bfc0bd2201100022bfc206b62027c),
    .INIT_25(256'h022bfc206b001018022bfc0bc1a20278022bfc206a4207b8022bfc0bc1b25000),
    .INIT_26(256'h022bfc1dd0001018022bfc0bd2301100022bfc206b62027c022bfc0bc2201100),
    .INIT_27(256'h022bfc0bc1c20278022bfc206a4207c2022bfc0bc1d25000022bfc326a3207e7),
    .INIT_28(256'h022bfc250000101c022bfc206b62027c022bfc0bc2301100022bfc206b00101c),
    .INIT_29(256'h022bfc204d8207ee022bfc2050025000022bfc20524207e7022bfc2054a01100),
    .INIT_2A(256'h022bfc2054403cff022bfc2052003dfe022bfc2500003eff022bfc2050003fff),
    .INIT_2B(256'h022bfc2500005c00022bfc204fe05d01022bfc204d805e00022bfc2050005f00),
    .INIT_2C(256'h022bfc204d820278022bfc20500206bc022bfc2054425000022bfc20520207fe),
    .INIT_2D(256'h022bfc2054801100022bfc20534202a7022bfc2500001100022bfc2050001010),
    .INIT_2E(256'h022bfc25000207b2022bfc204fe25000022bfc204d8207e7022bfc2050001010),
    .INIT_2F(256'h022bfc2b08e202a7022bfc2b1bb01100022bfc2b21a01014022bfc2bec920278),
    .INIT_30(256'h022bfc01c0025000022bfc25000207e7022bfc2007301014022bfc2084101100),
    .INIT_31(256'h022bfc206d501100022bfc01c1001018022bfc2500020278022bfc206d5207b8),
    .INIT_32(256'h022bfc25000207e7022bfc206d501018022bfc01c0701100022bfc25000202a7),
    .INIT_33(256'h022bfc01c010101c022bfc2500020278022bfc206d5207c2022bfc01c0d25000),
    .INIT_34(256'h022bfc206d501100022bfc01c040101c022bfc25000202a7022bfc206d501100),
    .INIT_35(256'h022bfc01f001d001022bfc01e000b01e022bfc01d0025000022bfc25000207e7),
    .INIT_36(256'h022bfc207d00b517022bfc011000b416022bfc0108001200022bfc207d93633f),
    .INIT_37(256'h022bfc2b00a04210022bfc2b3892f917022bfc250002f816022bfc206e420855),
    .INIT_38(256'h022bfc250002f818022bfc2084120855022bfc2b08e0b519022bfc2b63b0b418),
    .INIT_39(256'h022bfc2b08e0b51b022bfc2b37b0b41a022bfc2b00a04210022bfc2b2092f919),
    .INIT_3A(256'h022bfc2b64904210022bfc206d22f91b022bfc250002f81a022bfc2084120855),
    .INIT_3B(256'h022bfc208412f81c022bfc2b08e20855022bfc2b5bb0b51d022bfc2b62a0b41c),
    .INIT_3C(256'h022bfc206bc32301022bfc207720d202022bfc206bc04210022bfc250002f91d),
    .INIT_3D(256'h022bfc2b5bb20629022bfc2b62a2063e022bfc2b6492f21e022bfc206d201202),
    .INIT_3E(256'h022bfc206bc32384022bfc250001d001022bfc208410b032022bfc2b08e20636),
    .INIT_3F(256'h022bfc206bc05020022bfc207722055d022bfc206bc323aa022bfc207721d002),
    .INIT_40(256'h022bfc2b5bb208b7022bfc2b62a2f21e022bfc2b64901204022bfc206d222380),
    .INIT_41(256'h022bfc206bc2f115022bfc250002f014022bfc208410b117022bfc2b08e0b016),
    .INIT_42(256'h022bfc206bc0b018022bfc20772344a2022bfc206bc1f1ff022bfc207721d0ff),
    .INIT_43(256'h022bfc2b6491d0ff022bfc206d22f115022bfc206bc2f014022bfc207720b119),
    .INIT_44(256'h022bfc208410b11b022bfc2b08e0b01a022bfc2b5bb344a2022bfc2b62a1f1ff),
    .INIT_45(256'h022bfc2b10a1f1ff022bfc2b6491d0ff022bfc206cf2f115022bfc250002f014),
    .INIT_46(256'h022bfc2b6c92f014022bfc208410b11d022bfc2b08e0b01c022bfc2bdfb344a2),
    .INIT_47(256'h022bfc20841344a2022bfc2b08e1f1ff022bfc2bebb1d0ff022bfc2b10a2f115),
    .INIT_48(256'h022bfc207f50b013022bfc01ccc36333022bfc206bc1d000022bfc250000b032),
    .INIT_49(256'h022bfc2b6493232e022bfc206cf1d001022bfc206bc3232c022bfc207661d000),
    .INIT_4A(256'h022bfc2084132332022bfc2b08e1d003022bfc2bdfb32330022bfc2b10a1d002),
    .INIT_4B(256'h022bfc2b08e22333022bfc2bebb20820022bfc2b10a22333022bfc2b6c920816),
    .INIT_4C(256'h022bfc01cd82063e022bfc206bc20836022bfc2500022333022bfc208412082b),
    .INIT_4D(256'h022bfc01ccc0b032022bfc206bc20636022bfc2076620666022bfc207f520629),
    .INIT_4E(256'h022bfc206cf323aa022bfc206bc1d002022bfc2076632384022bfc207f51d001),
    .INIT_4F(256'h022bfc2b08e1d008022bfc2bdfb22380022bfc2b10a030df022bfc2b6492055d),
    .INIT_50(256'h022bfc2bebb20522022bfc2b10a20540022bfc2b6c920522022bfc208413634c),
    .INIT_51(256'h022bfc206bc1d001022bfc250000b032022bfc208412060e022bfc2b08e204fe),
    .INIT_52(256'h022bfc206bc22380022bfc2076605020022bfc207f52055d022bfc01ce432384),
    .INIT_53(256'h022bfc206bc20546022bfc207662051e022bfc207f536359022bfc01cd81d010),
    .INIT_54(256'h022bfc206bc0b032022bfc207662060e022bfc207f5204fe022bfc01ccc2054c),
    .INIT_55(256'h022bfc2bdfb05020022bfc2b10a2055d022bfc2b64932384022bfc206cf1d001),
    .INIT_56(256'h022bfc2b10a2051e022bfc2b6c936366022bfc208411d020022bfc2b08e22380),
    .INIT_57(256'h022bfc250002060e022bfc20841204fe022bfc2b08e2054c022bfc2bebb20546),
    .INIT_58(256'h022bfc2b08e2055d022bfc2b47b32384022bfc2b22a1d001022bfc2b1c90b032),
    .INIT_59(256'h022bfc2b22a36373022bfc2b4891d040022bfc2500022380022bfc20841030df),
    .INIT_5A(256'h022bfc25000204fe022bfc208412054c022bfc2b08e20546022bfc2b57b2051e),
    .INIT_5B(256'h022bfc2b08e32384022bfc2b6bb1d001022bfc2b66a0b032022bfc2b5c92060e),
    .INIT_5C(256'h022bfc2b66a1d080022bfc2b6c922380022bfc25000030df022bfc208412055d),
    .INIT_5D(256'h022bfc2500020536022bfc208412053a022bfc2b08e20540022bfc2b7bb3602a),
    .INIT_5E(256'h022bfc010801d001022bfc206bc0b032022bfc207722060e022bfc206bc204fe),
    .INIT_5F(256'h022bfc2500022380022bfc206de030df022bfc207d02055d022bfc0110132384),
    .INIT_60(256'h022bfc207662200a022bfc207f520572022bfc01c0e01008022bfc206bc20566),
    .INIT_61(256'h022bfc206bc1d002022bfc250000b002022bfc206c32028c022bfc206bc20283),
    .INIT_62(256'h022bfc206bc1d003022bfc207660b002022bfc207f520295022bfc01c1e3238e),
    .INIT_63(256'h022bfc2076601060022bfc207f520778022bfc01c0e2029e022bfc206c33238e),
    .INIT_64(256'h022bfc206bc2d003022bfc250002f032022bfc206c301000022bfc206bc20566),
    .INIT_65(256'h022bfc206bc2b04f022bfc207662b08f022bfc207f52b20f022bfc01c2e2b40f),
    .INIT_66(256'h022bfc207662d010022bfc207f501020022bfc01c1e2d010022bfc206c301040),
    .INIT_67(256'h022bfc207f52d010022bfc01c0e01004022bfc206c32d010022bfc206bc01008),
    .INIT_68(256'h022bfc250002d010022bfc206c301080022bfc206bc2b10f022bfc207662b80f),
    .INIT_69(256'h022bfc1d00320572022bfc327ab01000022bfc1d0022d010022bfc0b00201010),
    .INIT_6A(256'h022bfc207802d003022bfc327af01002022bfc1d0042200a022bfc327ad205a0),
    .INIT_6B(256'h022bfc207933641e022bfc227b01d004022bfc207870b01e022bfc227b02200a),
    .INIT_6C(256'h022bfc01c0e2046b022bfc206bc32402022bfc250000d004022bfc0b00209002),
    .INIT_6D(256'h022bfc25000011b3022bfc206bc01e40022bfc2076601f0a022bfc207f520491),
    .INIT_6E(256'h022bfc207662df0a022bfc207f509d07022bfc01c1a2044b022bfc206bc0120b),
    .INIT_6F(256'h022bfc20766363c3022bfc207f51ce10022bfc01c0e2dd08022bfc206bc2de09),
    .INIT_70(256'h022bfc01c2611e01022bfc206bc223c6022bfc25000363c3022bfc206bc1cf20),
    .INIT_71(256'h022bfc01c1a0b117022bfc206bc0b016022bfc20766223b9022bfc207f513f00),
    .INIT_72(256'h022bfc01c0e1f1ff022bfc206bc1d0ff022bfc207662f115022bfc207f52f014),
    .INIT_73(256'h022bfc250000d0ff022bfc206bc01200022bfc2076620453022bfc207f5323d2),
    .INIT_74(256'h022bfc2d1080b119022bfc2d0080b018022bfc2b4192f220022bfc2b00a14200),
    .INIT_75(256'h022bfc2d1081f1ff022bfc2d0081d0ff022bfc2b2592f115022bfc2b00a2f014),
    .INIT_76(256'h022bfc2dc080d0ff022bfc2b28901200022bfc2b00a20453022bfc25000323de),
    .INIT_77(256'h022bfc250000b11b022bfc2df080b01a022bfc2de082f221022bfc2dd0814200),
    .INIT_78(256'h022bfc09d081f1ff022bfc09c081d0ff022bfc2b2892f115022bfc2b00a2f014),
    .INIT_79(256'h022bfc2d10a0d0ff022bfc2500001200022bfc09f0820453022bfc09e08323ea),
    .INIT_7A(256'h022bfc2de080b11d022bfc2dd080b01c022bfc2dc082f222022bfc2d00914200),
    .INIT_7B(256'h022bfc2d0091d0ff022bfc2d10a2f115022bfc250002f014022bfc2df0801200),
    .INIT_7C(256'h022bfc09f0801200022bfc09e0820453022bfc09d08323f7022bfc09c081f1ff),
    .INIT_7D(256'h022bfc2d10a20631022bfc011022f223022bfc0105014200022bfc250000d0ff),
    .INIT_7E(256'h022bfc206de0b121022bfc250000b020022bfc2dc0820636022bfc2d0092067f),
    .INIT_7F(256'h022bfc206e40b12302d003207d9040100010ff250000b12202bff0207e004010),
    .INITP_00(256'h764f53d75f5cdbc8ded34c4055d5f8f84ec9e0444bc547f964766e72f5d85556),
    .INITP_01(256'h7ee87c46f0ff7b54c672f8467969797bd8c0f77ad1d1657eda5c5bd450ddde54),
    .INITP_02(256'hca79ede67cc9d279fe6dfa5cc9fed9e4d7ebca79e8e67cf0fbc7fe6de4ff51f4),
    .INITP_03(256'h477f44d3e7d4dd794a5ae9d45bf047d5745ed3e140d9e0dcda71f6cdd5e6d775),
    .INITP_04(256'he05afd4b7c4b5672dd67d07a4dfd5156f35cfc52e1517bd056e9dae65bfb45fc),
    .INITP_05(256'he1c5e7f3fc4fd07ec6e7727ed07d49e1f548507e44687ffa54f4f05d7756685b),
    .INITP_06(256'h53e66163435ad65aea56597be66df2e66b7b60e17b65e9f2e6697bea7a7b5f61),
    .INITP_07(256'hccef55fadb6bece867cff5fd52e2536df07fe2cdf267e07f60ed5363657fe5cf),
    .INITP_08(256'he7e6d875dbec62e17be7f775ef6166c6e7f2d8ee5a63587c56756ee076cafbef),
    .INITP_09(256'hfcf36b74f4c063c37b566c5dfa466f737c52e1cfe9fd6ae3fe67dafd5e6945ff),
    .INITP_0A(256'hff6661c3fbc471f574f67a6752eaddf65d6046674b74d070c6ffec66c47d5971),
    .INITP_0B(256'he66dc94acc5268d8f86ae0d5f648e56b657e6dd67561e3e4f048e6f66bc47df3),
    .INITP_0C(256'h48e56dd5f55d62f9cff0cfe5c2fcf2d7eb51697943e9dc76c0fcf453fedd64d7),
    .INITP_0D(256'h7c4b6150e35161ddfbc9f5db69d878f378c9e74ce1685af759f1d6eae07ec9ed),
    .INITP_0E(256'hfc416df6495bdc76615c4cd8ed4069ccfddc645fe946eedde35e74cf64436940),
    .INITP_0F(256'hf7ef177ff5f34fd974455bfd4764ea4446f47542efe6cfccf27147e6675ad1d8),
