`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3760)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5K27DQVGG6kX+kzvXCm1RYB9q4zmQJjdA8e9uyn+Lkd99r0fgweNYdsq
9stXj5LSD/ovmmupf0stG+75rBKjyhtmXFt9pvAJh+LJ7Zz8OtuNE8roI+hSi0ohAfCHY8fHPb3J
4x2G89uxjjwn6dK65pHuJf3oiNA5SvNNm7yBmHzvCbpenl5I0Uq1jFgKxKdG33Wd5C/PipyEFAuF
0ZuytMIQRnQ/iZ5ysh+RyTnM0gN5Wk0yvswklHDkK5PCQwKGKwSJas/+r4sLJq0xt3Plv+TUazIL
+0yZ3iJ8iuH0M+oM9ROOqWmDjvgjrC6N43ChHX/6PHYmM6i9Qggk62V69R1Nh+MJXHqz9ncqyFtc
Z+IDOvuBwWVFlcyYnje+vb4tOaVtdWztAvsk3NSuBv+eY9PqK4CVghHjfNBdac3DWd+Tx3zKSB6i
706e6FOrDL+zpQdExXsHXuEpkyXwtzcy+ZtUPpK23EqIjwBHIYmDjyqJxi4RvSX+sT2VQuXNbdrK
9qg7j4c7Y5dLd2FJX7dx82mORKvqvtDvKhO76GCszTrkQLPRtcKh60zZjEvbK8jSXZStmc1m5mff
HTss9tuM/UptwrGYbktIrcudjeNvLqrJCFSzs11RK91mvcHR2sfCvJ5pnTFUU2LFC+0EXvYJfejL
0KWO6/e1XLcQmevXWLrBQCSYvs5+XT6VoeG/k4Kh7kbEEWvwCAaFzV12hKjqsNFAGeYyVXsQp2QH
1wv3akPi270xoWoXpAKe7yIzntW67BgAWAjGrDOZGTIk6/md/VBQ5kfkzrY8jUADlsXGqx92yhzg
o+bXGSXdXZM55dDSs7gbwSfbMLxKajDh8XGcsHnvEOLb/gqKH3cqjGXYUUNukBr6RWqXxGe/ONUH
rjQ94RZkVUZY3pghXTQXp/7Tf3rJ7MggSvi7zOmOTHtezcTRQbt3vvwbfJLA9cLib38CuHW74Jr8
dds9uHi6giNFu6Xnfj95Yk1yBrCX9Reu7rgR+meYnvOQjs/wgbBKbsJKU9nOqnH9eFrNA2DzyKFU
9AHm+9y+JIoFE/BrEqbwijMlGzhZYlN2YUa/vfXV2SwFk6w9Doo1yizcY0Ym2HN2WOm0vPQD0t4c
Vr8f8NSLMa6tI+HUoMqumczwl4uXpXLVUBMBt8UXxECMISJrpf+XPKEzrYJoyS/TbSHgX1SwegkI
/6IPPF3gN8oJt9SA4tMQReEz7y4czdrXYoNcP6vvJlhB4DRlrLZCkGBi2FUetqso5KQlipgp/3+c
XMaheS2m1ofwNofh/c1T52+9SeGLzdFqN+48dl2hvqyrKZOiNE5FtG5JjszjKmZsohxxSRsf5iPz
55xZxhA8Hl6P41WkMO7kLfzp7XU/1LedXzDI1898uWSQzlHCxlzujFRHk7BaveXglp3UwO8uEE1v
q4ypeAYwGc27HxyHRdHOSzhb41X1m9YgN0Y8/PsiW7F5EBdI8fI+CCskrRw+ztRMJevKpQdHCeCe
KEcyWoDbiZFF747RK0CgaN0iPY5LIkp0AYFEgbLz9mDZyqsh8NUgv6PgA9ZOMPrfkNLuyG75Bjji
XfMKe0eq2Mc1PStlFfAiFaHA4GCKz2L5D8/X36N2Ikv95MwlVhuY0imwNDW9qUnaVWNnpBebMP/d
FiC1G/BzWilVyXbZDPcKQOQovs600FriR3gvNgLKp+bbL5vijrcEM9bnSYBGcgyh6aK+5x6oVnUK
W4qqIoA99YHlDE+W3gMOXO+7odBrwZZQsOeVNZH+Ym+3Ps4AzM4urdKXR5WhCetlwnMOJR1zZHyX
LYc9+bErXXJQw+lx7D8tQyS8eDQiKoIaiqRd0equMc3El+qnBCwbhknQk5pgqPw79m2yAKaYCIJm
DGqRALxDCPBNlBFRYvqC0cyGa+f0S5kZ8ZteNLT/ogXjt928Agg/k+NWvCT7qrSFPoNaOFX0LRBl
U3jG2AwRJLspih5B8B9JDsgSPFGxIVNNFcY0s12GQ4RkYJcl+Ds/ONV8EJJfQ+v+yrcY4ZKYHTUH
7FBl6nrD9VnL/www7sqKZWSSA+4v7RjCGr9II8FHOPcYE/4tEqVsi2P1l+WWaRp4OKhHg2t/JPbV
UpTR8mv2T0CBo20B2xyzp1lt+Du36Z4yZwXpZyaXHXPahXU9peTbf7nvKZXHNN6aHn6HMXZiHMd0
y3ksONTfnn0LrbfulCC3yBeASc6gd5WHxfY6kcfyln/6ff5cE4PfMlDIAivkRubKumAnFRPsb4AD
44RDZDAH6bA0wXzWBx2cofbuHZMWZvv0M0v6W69LKVWDzq11oaxKcXjpJwjW9jY2B7cgzstSKTvf
c5HAykmFLxW+5RTfUwtbc2dMS1Hp0GYn5bS0hwBXJqx0jtfnY1dC/ijw6Fj/C2exrOw/z+W4rObD
DrZ2rS09CHhqDlM8jdiDKsChPaLqwNlzvnDHzbqnLTlwHl6vLnIffDqUWSg7PdZTVmstDtGL3V4q
TXmLdBhKrtsoohmisvw9NtVTSeKmmxeLFIxEMPtw/D3+oxQCklRTe9YIUATtX0XJsovv8GIYjL+e
FlkhdZ+G+ZdXykjfC4cxgVXn3unBTobVtfDI5r/X1WFkA7x6UPTOB55J7xdmRO1cGTU0wEFOqqmR
btLhXT6Phv66L9WKQOJ/AAzCZoyRVkHM808fgcyivyLyd1RGd65i0yYvuuCQHuecrdHPMhnNLOXr
NtsxWcmNWi16Jxy8texw5SVz+WHk1IYkHxaN8t9s+OK4nI3GjpvRpXefpf+eFjDvW9jrmT7mTcyg
GhJLnLDZrN1/qXmG+1BssGuWbexA9VzyocOyBT+qT8EwF9kwYeCqWCcFwwMBS9/gDRT8sogU87WV
Iz+Edu7vMI31i3Q6MGJ8yHOse/RVJ6IM8RXVthMCq2VVZUyzKj/NxbOOvZMvgw7jBV1tmqARxky8
iBuKPV72wSS+NAG71G6BnWVFn5vvWXMpqAbNSXEN3ZDyFgP36DRRhwuuWKAHAlaj+Zy6rqPW3/D0
VkBdOzH+WETxAOp01bhKzn0t8ympJ5Ddp+o8TVmDeduLr7I8c4xbgclnnc00HNbmWzCEnD5T/Zoh
H3TeztUgUOfXsDUclb1SKW94a1Nhc0uSzGvBTsuwSVxg9a2BAzl9zh5pj12/FuaUMj2zweZmpl3q
K7InpppqKv/rFz+IA176YWonLmQCiwONIkZsZCSkW7aFym+CGkgc3RZtYiP1hFsGJlUr86IwjAp5
iRNqcF8toL1ndVKsXc1yEBi4xqxOQEHLyc5sBkI4ePiHaX4LQFo6pRCRTtuaVm85WaB+ia9u5Emu
X9HsKbdJ6ml+St6wFK/Na2Yxtegl0zBo4JlaxefwQLkRJXUobOQmAz9NoWzS5lL3FXP6L6m11cR2
6NkRsJUHccysQ/SWVH4NrZwmWcDDDxyX3tPBIISQSntic8CtMRBBfAk9yPQnIbucn/fn1aM/bWtv
H3adnDhKoqyz678N1c/PKLlxrNTMkGq3ErppPtT1hQA8e7pcVAPuvLS6pb2QF94LJJ7MKvdecAqF
GEQqEb9IEphaaWq6br0ekl++GDqAR5xlU1HlWsApl1F3g5Fun1HbnvWre8r0bToDFiw8InwEERB4
jhBS7PgOB9Dh7AbNqiL0/nr6lrIcM51qBQDk3GDW/ZS9BxNtVkb6ZhU+7YrUV3L1IV0XTTK6rYcO
1hZHaGZGmaGDDmuuCW0V7A0NSODGsqBWuVooL5p5qUDaLedErnPhIXTgXwrqX7g2cRgxn4ubHEPR
wvy+Y2Gp9zhLfCbRT/lBFVJQzcctH/l/XuVMPp5CgM0f9yXXU1DEnGQ5J2Z5Y8oYmnuqjLVbus+8
9PAHoYBNmnyt02qUeAPDb+Vs/isJeKI7QlnSG9qd/qIQwdUzy9UVL7P821TJMNZdZWOOB4MNxYBM
CfEvqr+jIVg07zKGw5nCzwj5srLEIzPkypCKOrAUUkuWG/o5KkRdYXKeM/xsN+HNK6bnWuUHLlwH
qvlRf+AP8GMye/DGw6PWs87/AFeCnyjE4VYzpfw2C1coBA868pCSQ0GWFM72+J+Apvc2ygIAvHlu
MLS6XFh5lLY0BaIOsazZ9YFVPrlEiq0HYAjtHQijudBe2F70FeTXpKwRV+VToaSwb00KkIxgPHrz
8rDG8JQ7cuqvXNrbgiap5Ck9yJx0qHMrBx1DlxQw3arBx+eS2Bl7HDUJN1PW4nQOx80sTl0bUvVt
hVHITR+cNeZxxV5MBW36EQtTKxD+AuG9OMQE4knCdkPeSVq21Iy1UYKAx7WCV+uSnLBGyV7GAr7B
DMtIudTirGyiDHYlwDFpRz10Sb8iCy7/K5I7Q8ZtHP0sg7n7AhyaxOXHzcWAvd8MzefYYDT0wDKh
6DmqhE042cxZ+EEbzM1AZJ8rsZyzzkI/DKl84bM4BwmqjwaD5UKeMt1/oJ1YX40NDgYlLkLRCu1B
zaDcK2DULF06PGlii7zjEBirXHATzzEz299FV6h4wiOjIZHMrHlBTm5hBz+YG/f+zuCZc1tScvVy
Qkjx65NuWPMYKmP+ghVmsHqfbCfo2iXIZ/U4nzTOQTjSncr3v6SCLwag0U/KqQpF7vBU9i0XpsMb
tCZMT7qIriN4ClHo2h/IoFXeNdU9gdRa71Jk99v5cO8RkiWm3RamudSpRVb/v7d7BUn8QQtsRwwy
ph7njDl4xizxmCjeHZ8b+p62Seyu9ezKlxI490UDkkx8aft9OgYrhb2CXtjT0f8AvIm/CeEeiHd+
zm51huHLhppL9LpwW5ncDw+zg/vsB6VTriQo2HcC20LQpcUH1KVrOoqwFl2iXkHLP/lli1kfOaiP
4f/g7v9I0CxU7+KwlmQt7WfLw0Ydl8a7EnXUQN8tNRXpucZiA7A2PvFcnPYuSgmj2pt02puRdeYh
Oo1aC0W9DsWhGPqnHcYuNGVA3atu7UlbVOpHUKNTkkYjqZRRgo+cJBE0ICyo17Qx9U0vL1RkvQ==
`pragma protect end_protected
