`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 36880)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5IQJj49NipZ8M+awYasSToxRopi5Djl3gm8/L0sS747S5+TDdrrPUCKt
i9mrMvtWGVGnN1VKZJiuVj/J/SkW8KW/vs2v1OrDSMGbrKgXftdvTXzPhRLfBBgRYQs8NMW0+H74
JApjy89HsDELmwmSTSkEAZGEcaEkfi1aRzT3bJV02bJAsJmsNPGJ/Z4ZNAGqhjZmoShaUdRBX7IU
IEgWILa7VX3kPCRxVYa4cwaN54az+X+kWfm7qUMcSSlRaWW2gUFsKo5J/mzjFRTO5GNfdkXywUSC
qNLVPQBnG9ZqXDrANlMQMaSSfReVdjTqt5hM1gdtChTCWmzVgee0HUtsIPuoEQ8Zo+aHxArMxqgG
daWb5IZvEYTYBi9+MQhXsRZqasLYZ/A5GKglGwZqZbYxUCsnjE8y/h1+rTP99sKdgHRn2q1wqe3l
fpf7GC0+bZnOt15hDUqeFjT8E1DRr7G+XlrNObJSsvD5FQ0PQFL8xu9Vk/JWQBWlbkhsYLIzY2pN
3q6ePuQYRyfyCnPM7ToiEMYnyV2kRoI5UyQqxieSPPLf9InHsj5UUUWOksp48Pu1befYKLO+htEu
3I1Klw2CPFUMMvt8yb3STwQZE8xHSDutBFN8QnNE/5gpr6tJGlsr0BOuFgUrk6PxLOZ4WaUEUXJ+
0zL8aaEGDC4roKoSQcRVK26v07SokdR7T8vnU6NaOnU8mn4ZKzmx6V40ybNWVxaTkcFfkHp36Kmw
vqSNfRXkImupxhjF8IRJ/ebJ6ujC9XskUmsf/UUPABzM+oCkjYAHkn/ZLfI77Kgosv/wNCKXNZgC
ThqK7jRgLW8Y4plv3Y0KBSVYPWfJ/50X63F8iPsd4xRH6o7QBHzRbEPiE4dJTzr7sdSTyqU5/Iu3
2irl6+ZC4E6EeqElVQ0scY9ia9a8vKEMYjcLoF03z/swbochmWzWKO06DMl9LBAsQf9RyKxEsscq
/RtakaNFNk8zkXocT+W4R4R8bCMne9Rg61qd/FGWqbNus+W7Bla07VLwiWV/38XeqPZ3WymmihPI
IMlmlV9/R94nW84CwFrd3zwVxRnQ6ThNIHqbaF9W/7vsJE7FTX6N0SROAgi6IIbAoqoftKNLcOy6
TKaWcdPVrcQKheo98baHEkx/jMsTQj/htfkKT5c/1zgdTuVUcwQY8qRrAzA/HKoRDgmASnnhBQZu
Sp7/gDcvm582DXi5N2zLY1TkKpP/hcOubKcHbjeZg+Ydsfa/0bcRHbKyuuh8BdvdciiE9a4NoxEf
oIO8wqKN+oD2otaQT+Kh5IJZOy280CRwQCPzSVRKFZCYH+g0mPZMnKcmI1w9yp8cG11QM5OdjBGn
ze6AKRuhNWyDpOFjRmnu4vC8M5WokmpR99Uauv5/gdPZa+df5s5AULm28+a2WZDNSbTqd54oGx8+
tsDE55K+cjccKFNBhBxvNtRfs02rw8joTNZFcus46wMecofyiMngyXaqy6/KQZwHB95Lx3zQ+fwC
QJccp51LdFQXe74Nt2KZdkXixC3WvHbZi4+fH734bYpI8QXviabpEegCoqmME1TF9SMOsyH4pjtk
UVDVlcQrpcZ1G2bxgCxYyZGjDrEjaJmEDUBgFHq02H/k1R4pOlzJetDSX3aQjPvcl1+b5EeIV78B
yxP49hpf9FU7CE62PWXOun77JVLk0BWXqPlI5yqJIHXyDGgBeFgYR9jYC6eSW9IE0U+QlFbSP9o5
IunBIUpergvmWXFlKGG+tldopjdy/5ICEiNlhjgBZ6ovtjgHJetaUkAqZZ+2SJo2Z3p395WZkT+M
7sUhawVcqyiNq1F6LEZQ+s75DtdVyM4EkB4asvqZy2BlBZXHN2r5MjI2ZdN/j+cy4+fZrtC0vK7/
MvtQy1iE+GJdaLuecBHXkmZPdJlUM0CRfsbnOZrQA3csCwaWHTOKnC7bOrs1C0IVvqOCa/CC2pc0
9RRzbfRhh9JI+inM4dqJld1UEAgz54rzctSf4w0eim5Gt11u4jeN6McFo1h3sDvjrfk8Ao9mW+IS
kwh/Y4e6b96uSXCDGCBWwGBpfIXifKz0QoNaMsVyFXCxE97DdBeI3U8bFhEvhwG0gpQ12pYExZFR
V6IsbMLzP8G9wzzacligIrEM8TRo9hIa3YV+BtjuRYyf8oxZt32bqs+p5Py5ZQNwuWbjvTUUPXu1
+gnEgClXVJX8VKfYnFPnIAYBqsGzqNnJ60cOfLT237n2VxSpIe5pfxRN4EwOt/is1IlLdAom7JlU
RuLaL+RC863H0OP37T7/j21tYAJzAczhVSpe2qHM049Armv2955hRVIrZPBI00lmRo+RLzFksVTv
N2/FLkiXnUBkyOkJKsRYxth0jIO93RY2OqoeoeBawezcMTOnn0KSGWYoukwVCOOY80bLSYCXd8bR
WUhJFB0s1DY6pD8uiBsfF+SaUFyQuqpnPWrfzZsvvx0dd0A3KyWsLpBsFztZPi412P+VGbtWB/j/
svv8D6y54WSpZmt5e41hY2W6RZ7VPcfm9vs4P/u9nyFgt61oHBvMUEPqjD3WLRmoAD+OwXc/SIa3
7gPnfPEwNoH/tZDJFNJTdY4xtLq4+2LfYUL1lQUsyrwzymEQLLlXEPD3JFUJsthWG/ScKbT/bYL7
DDOPsz0I1YNAJp+5zCF59eNO273RnTrAV2pK754lPR6dOiRLuCWhP8PG+EJbhtNIkVHCut87eaEg
j3D4TxjPnrOHrF58lxv2h34+MeJctMLYruuOYA+v9UgnABde6bxA6ugyfq/wKxeOxltqqRc2k7yG
iM02buIpgeu5ZJX/6KIVhNgXbxQJSYFPc9UlMc+/qhVw52uqk9+7vr3uLcYGv5etnSJiarR8/YUk
PYP5EhuczuPMoyF0L+NUkcWs5/IEyis8xorcdcFE9pA9m+PS206FZRTstLbijHyanQFNlIIIHQ1B
RiHwFIYTQi2dLgzA7BS8dC6Tr0azmAJqnygUsUElWF8ime58KovYYclfpkm4TtEO8CyqGEOwL9be
6AYA0pGw6gwq7B2R/LytjNezE1/WprU7H0itxsHeaqORQ0QYgLwQoB8SEkDvZovALXO2xZuYL3C8
8jHEaOwWkPOo/Vc4RyYPwR/FXIG9W9063VMXHWM2WengVUCae3wqk9XRT0MrF3bYT3couPITNKcC
4eyXmOOY5OthZoqJXmAhtCE9D+WUZJlTxNFLCreNflQe34kAVBDxvB+eVY0V5QdaHfMKGlO5Sjhe
Icdl9E/GvOaCh6w2aQ7Su6eGiE39b4AFY2asCa+lT/yn5plnBdVvh8wv17MnKqY92yy7EMLHMJOf
fjF1z06+mkGDA/Mfvt+Bq4klbUE1NyYjffy5DWGOhIXfKWbxoG8uYA6M8VqXCBEeO5BzY+dHCccP
2m6dXpuQeC8PoF8PWqKRzmw6MYOGpbjMweBs8Jmok8+05cYp7jNfe4c//ODrO62YgLgf3IPst1bF
w62VuPemZVBXXjJ2a1N+japgVUu+0E8Jcs6frmgky32zR6cQJ+TesiLM8WaeAPe/GPpakUav5MfV
OkXBvo1F3oYLxgrvFk850pHIuuWC/ZqQ94fRAcz0wDMz67ulBi0K+r13YpX9yJShX7SSFApF8ytJ
keClU8E500dOe2ycytaDMxNVtuxncBbFyNzqxQmTgcuS4qsinCFh4j2tcnd5Zo1SbLd9sL2/PgWH
AKrSa5FROQdOSMFznc11vd7tOPaJRWKHf51UhyDYErXkfH3llEDXjlfzhpqK/rkDsQDiqGUf8at1
lsk1Pv/7tbd4PVeFs54Tvg5E4qoIsjBiOKDQGMbbQw00Fvs6gfeoJspee2dVhj8ci0mSJ0FVzpP3
A1CmXYOO1ZRGDcAllT6kcmHRFH3xTFfX6gyM6Nmw+QKQ+jg1kVFWzlww5I/LaOyZYOfOI9sr8Zjp
BsXo40i59stNvTvb5R19h1VX1VRD8LR5SPT7EWP3Z+TRJaOZQ9xV3j871FDcudycwcMRfM3D/0KN
3C4RM2CN0uIDqXa8oZWuGz8uhfolY5cO5GTpSICI8rlNuqgHn3Tnp2R9IDnmc4PrWHAodhh3LLdH
TYs2pNErP2IoTsliNEx3eepC1zRaG2N+a36z/NF2MOhfrXy9fqEGdMDG3seQuJ/ifr3qlt5IRy2t
X7UcSYmHuXNFdBcC5N0mssOvMZ5VfMAJBYPpscnx2EXsFKBt2ktYqz/fVwaFHZQEvuo/wgpX4DJa
/QdgdjkkYR8aQFuhuimWh5PmRF2JhuU38X+wAId/6J0IG9pn+YFbfnZZmtoGc4MSXJKNdNp/V0/p
NfwQfpoTRRd0XOSa7+7aY8wterOLopZRP2hrX/7OeoqgnpssjrnW9JekrxRrsaKrOHF5HAFuxrWV
DL9gqArnzK2+l1et4g66A62VIFZF1r56+KcFsi3Jghs//CER7ehDDFm4ISHgevirnjh9nayETnAx
ZlASiwNeNFT33oD+ZslI0LlyNsH5quMI1RwEKfZddJDq9ROJuaEfPDhbCRmKj1LZ+3vff1KcO4uv
cjZEMDl7zvtkUQPkqr0hTZolMR+CoLN0B3lddYejuhSb905nyISiQkkX8kDgn+CXTc2wr3fQ++zi
6rglq+xs5VZYufce9GQNAr5OfTyefS5it0UxMDv/AcO1hItJxLrojaHEy0SnfLjar79djCdbLR3v
KmJIGT0Qzah0nKi4Bv7lD9igcwXC+S4YkPMXI1mZ1En7MJaOzOGjaC3oGJW6GfoTUhi/pHcpD1YM
eW+DawFxkx/i1qhoYvCItkn/4VgVPsZfqpzSBrxrl3++dyoaqR/0zIT2k1o+dHq0L3MqjJmFne2G
z2B1aS+XDjEBjweTqx/5oDR3KyS5Cu9ukQv73WiGX1drcT6Qv+3sJrgxkLXnZJOxWIliT9oJSZh2
55EEWSc34xCLWpT4O1Fi7JcwrqldNrxdyR1Pi81UFus/RZsdJBBij7d5Yaf5T9FegaFIA3RHgHKv
jpgOwiX78Vm4Fi7y+zQki2rLC/Mdz0Ksf3jTG1JXSDVpkfXMnn+JXJCrFGmjo1xmH7Jybzaq1U5J
sWzkw36qtNQV9zT+4dxsnspiKyIjCOb5qxLf9E2GCKE6vOQ9qYX4V602xkVumw6fgen2heecDHkZ
kNwrcZHVYQ62djVAJ1MqXUPbF3mK0DAnHcjj+0S/KUrCEHhoEShangbVUXTKpN3HfqBOeXpx7oEv
ZvTEatqkfig3xHNHzxI2PmePtsMIXErPQ+CAOqCyS3wnyt6tTrTuKiObgwRDAuylTtDzzqlqm8Fx
DScNX35ooIoUwKH272KUKwkTzwk6ZX5Lg9cgZDZK3jvq/f43YGJkT3OjNZ3CKp3Ls+14ZUhWPh+x
5wvNraqfeU4doozd+9+w0wfVD/WgiAfCN6vid/i1OnIM3xa1KJs2AlpHbHpAV0pynVasajb1b3cI
I6b4aocPOvKQHfVWcATuW2gImaQULunXg/7j1HlhILTFK0TEFJwPJWMRKzc3VOGegwGtXvRmHjYl
oIGcSnfRksbWOr5VjppupzdM8U+IyWmtSGMs1fRyyDsMwU1PmBOPM860Qu3l0ebVosoQRfDUJkU3
G51jRm1eGarRQjFrpCX//G7OdDYKB7XCMbqc1osAAopQxkVsbFwr2BeLg8kSJwnxIDqI6XRAYkiN
aju3toChTS7tPichq1f6h/BqcNlqsiuWQhgKRY3by117HiVEz8jQqenfJyUAwJvI4v/SG4/bOav8
h68UbjdYlvDG9bPh/qa2Zel2DLHwduiHD4DY7fD554I9AGCEym02U3GA+1BRRD4UAv1CHzpZ2wUq
BSBFf6hgwXC+MI9d0P6HKfSD/+mKDCsqz1wzBEfob/tDZ/t9qmQ19zg0r8hsgkVQ9yB/zZeI0P+p
aiztUbFZKBzPCkfnIwvJOGlpDoMCzxF00Cxu3R69ruHzi5PF31mg++73IclZazOfcyE8xVjTRNcD
P1sF4H+y/+/r2zjybcaPkKy9rItzkw8NvyEIWbEyiOqCCdMiw+I5wTCKTTRQ/sXxo34z16iQVzEU
x0/mTMseAxLJ2WW3XnqJZw/4D6UN2rg7HJN1UPbzkPEAn3wjXlMCaD/5HSwyQt96EJseU+AqS/VC
laET1VsmYTro9xtG5GOicppMt139BbIX+zc/N3j17M+biS/kRdqZjC2VMYMuCCjSJmtCREZ3sTrF
yAjm4RW3bzxg1XjvUXxq46J6LERU5OjO5WDqMwX2+vIZqCWd+JmAD9DawyOmAW99moTK30eSrzOY
3S3ywsLdxRgJovmoThPxbYnRwAM7E6aqzwPqC4R/xRe7ojYqNkUPBZR7IO/hNnyNe1zVWaHreVuj
R3jxdETgd+cZasLteDdwohFf3mpUUbPjwYzwBYEaXEOEPPG7inzVV/SE4X3379lkpUqRP6rAi3DF
0vNdvBl1IazhlscZ+ENUX0+NewKI/wP45nd8iVo+WNes0XcmA+gyHJe1Ru1xMjvftPVUug8GLYF9
oJi5pd200nrU0lNjoj+zxvD31cw1vdYhTIoTn8TCYzDyixEZOXMLqfwPVuQCI1gyU1BKB0GBy21U
2d3WbKxWuCcTX9XPjZMB7WqTY/LXE1icygNQVO6FSx8EYPUGSt4pDHXEjxYhbYBQAtem/DgRRMOI
iPYH+QBNxoymsyZidl7fSPcb58TouGoi+h5IhcsSFEsmslqEC3x406qyTGFtExTSrwWvaG7lbg4i
wjP1Aej+efOPa/Nzd3lGR5460K57Eg5WUuN9N2peff9c3BO8qOuqJTTOyiYZdQMX8MeIYJ+Ui3Gg
40471nHJWgtME6xaUTIc+pQdGIMtMs7adPYVyxEvULNisyNvPhatPjZG1MzLX2jlNVnokfHNDA1e
8Tw/XUeh7SYCuzUL70+XIBXBLh2IqK1qlDC3w/MpL7dkZMfxTmTeANZrXg8DHGyzTEJeV6/7gEUd
qPKUomokKCmo4rr/reOwCjQsOejSOHJkWI5QRrMXaejvo4ryk9IQWUeFJbJUnHbCvb2Mq1JX8Igr
H2DiEopOPf2sQ+kBpAVmqoZFVdEnAz59BaTJMCbN5aAE1JH9H7+GW6G9In5jb39vizobsGpbWxtp
HoLXU4gNgjXH0GQBcN9VM5tIPYgVzLyos5PEJbCUa5bbEA+72RRbed3LjqDRsmVzOVVlUxQMK5gD
IKCgVQVeeXKnKIioyfBOrSaqvEfzpZqrTRDkGxl5Z8r0Z5nuk+QbMx2aamGOSSyIQANJQfYH2TNh
5y9OHbOW18w64W2RK5IaCV1DQLZBsuxdTYyASOp+wEgPHe/OhZEH+kywn1KZ2UPBcKtJL9X3zMB8
lcBzAQlt678U56uH3SWJh2OrXIIYN4G8jIIDzpEpVbU1BScG1SkrkKoFx70oVxoOUK29wF6w+zdU
+dnipD7d1fjylg9Rk6o/CowM9oBHMxMPqh6LlAi7f6gxH8tEU3kTv5QfF7OtEDFsdoawBnq5sb+s
DL6CSABkt0Xip3xIisA9/mfgBKHnPXQDuIjGBYwOagp3oO+zwI39/tjDp7F+OwHHD6jYPvplH14e
sLxuKNkAKkXAx8xwXkilYYGGunc4baJKwIPyyU0gV9JqAm4S36HcC5Mojng8zSI8hDNxbngKN6no
2nVXL11HD4KBvfULWfwRnhHqH+9Q/VflozYOJfaVePhsmVqFfYbae1+a5nVnZLGFIfRczYh0Hjqn
geh2kR2/90p+eeoxbrkrCQ269Jx6pjvJgRz213WDnsNeUpuIbzOEXDre51VsXJ1Cd9vyq02Fd31g
YmttJxq0byuzCGdYYoWYRzBUyrs4nVTVErqv3K6F5PUTkJxYPzI5BsGaD9roNyQzuWQtjVbdLknt
HJRCeSy4nhGI3ym6Q22qe5P3nuwdVWw785D1WCNP5jvQz8/pXzw+jjTU4HHIP7V0+DGTMdUjwev+
FJbzbjbR4IOKX2A/72p7PG6IqNkC4TEMAURuUBmXJ3bNTenTG7cxrjYgeVQWK4AraCHM3qpqkYsp
eogeVvzOhiVjIr0o7oypfT8I3/7ihk+9buHFHs66IGhe6QpM26fZBRKFtomapb7eJrqRX4y4bMqs
+5lm1EpMw7ktW8KUgnMHPQlPLl1jKvdkai50aRWt2CL1dXFBo0joZbyBpljPVmD/OZAm/rm28DJS
swz/ZxAm2/Tvt9gea1//QyRBFM1UVjb5NwHw/LljBRrBnmzwxCsYrQYz8pcuNBZxMM5lL4tMqNf6
dQmo/b2tUPM1zjGPXmo++MOpwJX2OVjhyS4+eJvHC7NMKB2GNSzvhsyC/Bb/jgxCr4MJrk1zVgi7
rxXxBZvaqeQALYRBHIsjGhowT8Co/mhqsMDr3aRB4ZF4idcU3tDX4ilnpCFpKxBeu4YjQ/3i9jOK
4I+CehKHQy6f//GgIsBFXAtrthnw1lug/WHtjd11L6oLiR3UiblhmAkWT0HMhQhb6+Cx6bL6pgfB
XGIT7h6U3h5msPyGMdkwwYDsuh/cMyzbD7JDSqvaz6t8bEox6zmJfu0jxejCP4hZcdm2SP/ZMMCP
3C2pJ3rUk/ykSWKxCiU0n1toHctlhWkZNwwYCkVoGw0xVdCDo7AD1TiciuP/MGo0qO0l96Trf9TR
3E/EE/u2iw5Ck8JM+coqLE/oQRakWLKS+T/L5N6njvJehK9fUeN4nd6VftA7hJ8aMLYseVCF1lGq
4vnjHWKZkcUoHxL3JfJXfXDa9fJkCqpHGwB6XHsa6xOHwceh8ILSoWCMhEbGFYb/vXrMXXIXvkNr
jxL/az4TAdA3/TPJYzz3A9ghH6KoKt3bN2WK535PzCX29lvGvdAgpwBzFazsj4eFO8+m0g1N/8qo
nev6a+eEEpsNzF2rUGWs31k9oliHW4bne8gGGlVnNoTdPcdm/51KZMSK7+EPsp4gsny3HaMwEoAo
yavurP9EZQHKNmc9mHmIHdV6C7MurlAlTtJYlejqvkS9ntVJV6HD7R8YKkyMt0Cj/KHIFzOXvz6p
uFkmjdwTfEoYJ0u/ni/kCFCHW4vOhfvg8ilY+1sR9TC4EXDtCI7QHbk/CktRqr5NTJWZRGnfeTKB
L9EK62CaIibk6Upb+oneAep1uoz4HolNPFwZEncbJAiYq8LrF6yrQmFdBT9TNgRjsqxrPZ++Kesl
CvTyP2ckywUX9dU4HgVov3Lb0WLfGzzGdnRvaWvBLu/zxVreRkgUywg94sZMHzB7/H+lAoEQWykj
zqXAr1thIW2bWubvsPyfUAXoBAGd08QYfd6AuL15z+3KHiMM+Pc516fPNK8E6XLTbwxfGQzh2cLi
4569y9oakk5692NBcxceCqst6o8U/e5Ex57e2Bu44Ri5av296+TUbcb6yCR9EelwKWCDsnyNM3e4
IK8z2CLRUGz7zz4x5RnDq999CuJ3Mwxau36tETGIAE5L/1et42i/qerkB6WU4PksVxxbn/eGYGCj
dEbJg5E8sxO97Cv1CqYKWHrMXIfyc7gzi1+TSKWgd82pcG+QOqs/a0lDCLTHlRtaEkU7iAAswHmZ
o8pW7YBI8vRzhHgQxvCIFt/MAABFBKMrXHoujZWgG/1rY4kVBwWQKoctKGKxZneeXWnNKDVNz1gI
fqWb3gakh2VGvBr51uO7TQIl2DX10BlQt5xeK4i9J+LpkE+oaWNtgoniB4nyZ9A2J795QzOPFK2i
k6oYem7PtNNYcC7EdLwpTc9vbxpPZpmrcCcWCupzWEb4vxFjON1ErxLzK8juF2NXPxCeKkKhjwyy
gft1Jhoe7xlXCXpWfTT+ksrvOLukGeBpTpnGxRhPm5hOgyhZecE2+01T5o2Txq7shb9Lw4593m+N
8Dnpaqeq+WyyahrjBHBwAIxFauWCp099Bj4r7ATl8IAz7EAAUBHe05d79PhWl04HcEQs9D6bTijT
BY+QnhoSrzhXwokG5t1369+CJou7ZT+WMp0VwAXgS3nQReGEN0Vd7dPojVis+KoOKLdBoAayLrmC
klbmFN1SSOOajElkYfRRh7GEOtVyTboYBMebE8IOGf2DnCLRdFhUlSVWIz9cgl9xb/wLwnYYhdOT
YzYjnlPofhVBJiZX/Lkc3C06jyqSUgyh3CKIyCQYKH9eOzXHd3i1v2q7qaqGuocwvC4Y/y8ILcPS
xYehxyVy03v6pwW+B7+cPCWVOAyA1NaetOrb81A7wCT64XVqe0Q8uEEOrsdjBGEZ6lfVwCiQYcTu
GrjpEfCxRRIxyYf30gMc/myBbtfREY+pu3iODX53zpKkXvJy3RiBYnEbJg0EAuLXPNQVGu0Kt1Y0
3CugpShC5X2deoiZh/HRhH/NX0b//iDxdBpY3/J4P42q8NdjpR7e6nWc0RKeKkFoz7xgOfH0T0uE
8ZNSOj0c6cefK+7HQqkh8mSccYzO0VjLn9D9KPrxLyrE0Fj7JCMkZUN2/aGJpjiQ1F+U20IwRXsh
YxN9xNA4XNELSYqS5ZKOKMXj60GPpcl/nGS3lgpxd2LwO0Ctpoxi3uriPtkythQMJKZjJoyJZJMa
gEYsfJFI1pAJdP0yEmNJ7MJga+aEJdAP3BZIxyLGzjYaZxtidfU0AsgTTZ8iBg75BXyLNxvkHxAG
vPemFCSpl3WJe2X07moo6leWTeA/1fee7lrAzbC5Tfb77xclvCbBQS4+/BXpArNkZgJqWETU2su8
EJzHc1fJPiSRjHzMPhLut87Pxk4T3mygNN1a3FZ442Q0yU6EMemg3ZhP5C4gAjxZoPB5UMXEFw0P
0nbAQUaLQcfaSQwKadPj/5dNElMS0MblTiywlU1NhWHkGitYew0F5cX4BOMj4AMBdJmmUPGzHoq+
RnlZ1Y+9Di4zaf+j1eidAOtJn8apO8wPHoyI/7wsEcBnCSutNfImZvtPf285g2GLh0frkXTrGXZU
ZvC9wttbgG0Z7EuXe11tEUOm4zg8r0lqoatwc/8pcOxR39JjnWbJXGPKxWd/VWINQqENVFPycQ5g
c7OfMWCDJKH5P0ZZpO1Oe1qtuGr5OU6czo/fc07IKYsp15x+gzMqnF0VuVPOiLl2BXbEnFj5wWD0
gqgv7oT44DeJ+sBhPetdlu3FXDJyFuImgYtfo99q2PC2ZXYsfpog2Vd/LE0cL713Tzfx6zD3Hhr+
BzG4/LPmyY3Ma/EeAi4KzfBCvagGUAccyr3ebn8f8saNYJOFuFJqxSXWK3LRL5+89Fw//W3gzCzp
RI1Ybo/BO8RqSL3DVX19/mml8LRANsiNYvXV4UE/4k/888CBnLqTdmew6yzhxn8nZsNgRAsebFE4
yWIRZFymtC/D/6yADhHn2xnh4vvXfcKNYvV5LY1Xvy4N5WuS4iwYbLN/DObMWyR3jvWkQO4scyqU
5BMydO51aAxQiNK9NQYOXtETnTSYC400ksXzuCUoDoNgW09diwln8+FTBtXTu80jOjrc5uQzBLUD
M2Fm76cw/uFmY2gBGwlVZDsNkGqx6as2zfaobnm3jVzzJcBN2NiZQkXnczbHr0h7yeGMpYWjfC90
8IXEOAvgG9mMAwgWK1MSsYogyemFBrmqX+NQPNov1DrswkFkFJdsucOsvz2WdEU1VedXsqPEj7Ce
OtCh/XnSp6nRYF88e2OHtifyaElQOHLBhrx9q9/slFr8TcCgbatU1tUim0fwiYcYeStupRhZG3fp
SsWMPNjt3/wzU/6VYCZOitOQjzRYzFhQEa5UJ09Iem1oUJf0oaPZnxdIJ1Wpf8i/YDz6wWmnwiaE
3F9wMZbrWaSZTt2x2i2BrI68nv/CQaXGt8qU7xTXYOCRCklxrGMg02be/v/c+srZO40VQlKxPfPR
C2WXJ15YoavtJOU8Hfqpu7lUWpmlErKmKxKjvdVx6u7vbh8d2txe/lK57gQv1jdjFf7sbWa2SuTa
yPM77m7ItYBJzoKpZRfOlicWaDR+jyJAvDuCx11j6P9SQqvG34ePGquFyOmK0a8odoy+W7PskEka
MLWL8R+p/D0ZZZrPESmdp0GBQxXTFxxKxqmkdN0yDM+jhzml+w9CiyQ/UounaXi4fPMI5+9XBlGB
uRQ2xcKAp8ZWDG0ogEp6Ayv+PVMGXjIBfSR2NeJOBzJ6eigGhBtkMmllU3fgAptnNZRokl/wOsOI
7hvo20q5r7WVOXH9bieODnGPGQxYWwKuLxFlfpgZFVLM35BEMyLgJ48dLMVafz6gAF979uQUlnVy
CwWVTHZxk3ckved7NcCeQoMEeLdmrPTFLY1jVSjoy+4mfyassl1QBESlJqHUJLekFyX9VK1w8Ebf
Br0/SeFeocqOoWwRoghAFF52mVVSv4OsM7Z2Hu9xcJQQKJ4Ot0262kNLiG91rcGv2y5jqc3cTK30
cyZ8UHxpEqFezq+PREQ7okxQPFLKWcTqHOYZZuG06SiAJIe2S8BD5fa4n/rpySxW77ub2TiGW2x9
o504I+SyQWp4ZghbHE9MshpklHJlBeruacNeZmCLqabosC9LpaC3VPzyStWDuqyyZ/U6O+QMVnA/
4lHy4rylA8HHHsXj+sm+kTjhdf9VGDZZn8TtOAdcYNpSzzudw510OIbrRoK06YsA1+9j3H0wahGK
VQAboV0J/ofuGNk2DiR304Xi+Wa9a5mbdv8O9oKTG3j28N5Daha8s/MFUlzABsMScXRkkLkA3eOg
dlrPiIz6drDb8BQulQ9OKtECFWHUqp9kbA6KySrXxBwHnOVyAdg3jhTRADTM0STMTXG/6vjDffuk
lxr5eRnsGbrIL9Tbe90I0SKXQQqta62y+A5CvEeR2Ylw4BGRAe8zZ1J4HWvh/2j5BixN3M6bLHtn
1MJ/yDTVgGO8kK6gN8Y+jeVtkBxnb/FMZhkTKwybAHFGlmH7mWPV7U59zYv9JWWESQgZSygh1CA9
VUlm/3wg3j4tbwZfyaSsbIJc0ZGJUG9w4F7ghZj0rNz60hQxxeBt0ryK0RXF4vof32y24Bytb3UE
6vwuIGm3DD9+9r4oKoAgiGy2ArzmqJgX/GjH93hWiGxKTJW1mY0pN8VlclpW+Fd8KI3j7+nk/CZQ
mmQSWB0CUYgU6GcX30s0WHhyPrT9x8+tK1gmYYQgzPtRT45jJY+PqrjV7K0NDqkJAvoMDO9ZhKrZ
dXA2QnqujNrSVWFJhwSaspujr5lV429CRK9TczSvGMlMeDer1FUv5bBJF4bYkTW/pd0kcN6Z2l7u
ozTZZ62uFLj7wV/z8RqWw3TXCma3s1cASB4+cRy/kycLj7OKf3cwSFDUA72ZxXvU9tBhQAa0mLm9
HmuDWH8iX0V+vT/hwBXbKEJV5aVnvWmnptrRXJJb/Ap/P5ROpOMHyyvUn4DssBCq2n2oTAvWPmlz
TQxTD8CeFn6/97hV2l74PQDiTyOxV9g3KIvnXz/OQPzOVSDmLUcs3yB9j8oFTFCYbuSgA0WH0Icq
roavafN9qCiAv9d1OdoAKols224JahTwZGd9K8l1qV0fnLD+dCu2ZVU1/3GZcPjapUtdhNEWLOUp
eHudSfGzxBMizX1tWuuj0qEu49MZNOKnECMmvZ/gLUoz7ABL3NUFuMfzgJb9oB79O69tUlPqoLw6
llzxFb0e4ohdup5WjgX6vduKrLVgBVOzrn1GlN/viIa7BmbK+RKZlKrazdWEo3vPI6oIaTWYJqH3
1MGYIw+f4sszdpvg51gAO4IaC0ImD4sLxaO9l9TI2SExwLSpl0PUGrVwVMe1XZNJYqsQYkIUIOR+
UgpikttF7XIioZg8Zd4WZvL5GVbj34ktipBanbBUXP2M8R0Tqh0B3vihYJuKD9X8zW+jHHfs6+a1
pjkzCKBNQ2R4DKNCpyj7zMJE+X5CMclb3h5mGxrOf7e5Gyrj+vYWM3mJYaYJnjZe20mtYW+5ttzZ
HTp0n40mN1jvB00Q0zhhdF8+4wzkQSpKvRp5SVIJZOZ0nNS9PM+QXDs5IncoIRQHSbhnSC1irSBJ
eO8kIoSLI96f+XS2v3WluRpUX7fz6/Jn6EqhRpRKixMa37Mhlwn//GUguptTXNtyaHsgF4IhuqvU
NBBEqiak8064dBqFqJw3vxJi2QTzy4MNj7c0UOUBbl5DFEvGzEcH1X7394LZsXpjf/a4LKc4P7IQ
odjdDqurl9dDRll0AhObv8IN2vD1+9vhy3xYz8hgqePFomD1Wezitn0VHrGfU5feAxXc3nFRYavB
Wdk0j6umQvxR6OznEoJLokVSgTd2x5DZe5mDAvNfh+2PASf6ZwIeJh4jYCdrQ5QaFjFmm6sVzwzr
Dfx/cgmgTzOEUxD6z3oyygEJG28XWA6Uw7LHeo3pkgPscOIBpl0gJHJLCleeUTEt64ujwEnAJNND
wijZjIQrVgAKVJg/fgXs9IgBLPymWxEXKxjs9P4lYV6LK6Eq9jgyW1etLPmb/7iUkdEkj3gQb7so
S6C0piNp198bDgZ+Gq/VHMS0Ow7eOZ59bZYwyZfdZgUykeiRJ/VRwhG5ueP1tBEDLNttyKKDXIGe
x11KBgBE5Uxka8jTZEoLA8x+u1SHndmNReeVuI3vac6Jj6T1WE/236Z1px1onabeB+iGxJDXPt6j
zq9Aco5eg2Ph4lhT5rPfbkc11zo8fY4PyHCo9xbXxnXWkAtRiS7cIRkbdhZsgJTi6/XHGRSdWJNO
f6rj8D/AfKk15x7+F+4ziL466ywwkm3vAYtJwrh5M6DOFwBqJkz5b6QC/zdBOEaHHz9mG9OUmeMa
iqqV5iOGQ2uWvT4QaewXPDOGNI1GdkGQy/rMeaPSHo5c57REfZb8ZNt++28yWGR+PWwnMNQmfUv7
GC0mc5KlqGMM0KfxsaMu/CP0RUdJapKrYZyoftC33otJYhGxRhE3fg40Eg0gzUnQ8rKLW0o8FH5m
Szer1XLpADck22gxW5d/iOUruzJ2Un+7nxpRvyTK7xan8D8VcPZme9whOtd8fQHtIWPb8kYqxbsy
kicXpE2ruWpHeJNGB0GUbUFf0kFoLN/eG2tHETulkju23SbJDrt+oxDQL07CBOXF7TVhbYmZBYB8
9Vq12wlOhqV8htKYTVWIKiRBBMmow9DjotbwIE6UI7zuEVI0fb8MlNOHX1yTvrgau7SfJtQty+ho
LG2vpGDVMU6zPAN6qnZt/8dRzrLM5oB8iaFWpS5iJ3S/k9JEwLhw2EC0Ve4TRephiOEOsOADEoVt
7K8Zix43cZsEMu0o8JFoMk24c3WlMR6axQXXO3gB8guTgfEsSdauVvIo+4zsrjatXYfKGpcQVVCO
ZCli7/+4W0WWl/UhwDit0VW1RnPFn0AIh/2W1J/TEAsFmCOT2YyLjKlNXQlsj6NKgb2Pu8BL0JPd
FbKNxNL7yFw+eF0htOGpbgbH6U5g23pV9CE8saiNneYwa+h2wO+P3t1zfODIfCkdjwr+1kFjFOeW
MUj+WZgYjLu1DagOx0FcmgK1oIspVJ0v3UYmctt0kK+UQz9XJ8/N9YEoreXbAtgx7xrWFxEiywNH
ok8yKWR0tZgwLLDkiHgIyqez+2F7dGJftxUQ75i7Uc0j4SswItfpAIX2JsdkfIiTnlrv8puoCPti
ECOSGhG+Pt5wxodn25q+SHAboTmXmrpL7Hk6W7xdbYbxuLNmfbK7XU1eHjLhE2mFWrrApbopwIzs
YcxOM9Ue/iBntVo+UzJCF5yO0GWxVzi6H44e9ttnbgPj28HJmlKl27Bq0qOHRClefBiXJjzYKQiJ
opfJHLQRc9ajHNnrWWkVJFJl/UB18RUIvccDWy9CfQ8/dpMLy1vGQzafInpy2S2liZpwZ874JVVU
B/RfMj8XPCrzxd6AjKjgW172AafUF0ddKLt4jSxivOu0kVFxiaCg4+KwHgISPpIf38Tj7WqYzayC
rw4QPIhWo5Rn8/fPrZopklNBUWipPBS/55HbxLiPHpD8F+ZtBnbMcsVF7Zrc7ILneUtJ1WH0VNMe
Bwkj17IJUuD8POblEIxwuZtNPoshYspSgtCXnICDvhXbbaZWuogbegdyovmjhGCLbWYsbjgMmiya
ihTIDwJZBcHfFVZm9/nz4CuGa8wherWoiP+G8tX6eEBUaNSKA1gWSv7v6/sCeiBVTes1ZTbKQZSp
U22hmEvRiKu0By9xOrRYv+wfx0rj2U7xq5xvK4eTgHr/9EaVHktVO0MAmEhLrwVWsEpFoKqxk5Dt
Hc/sSH7UeBAjlos6QoixgyPv+PaRwHknT4Pe+t9254PhcnMRR2ZCroO208QpvlgbXnQdQZ12/N04
xmbzLIdcbZvjvK+2OjcEudc+OjG8saLkQPYnYs2vDMXjnO8OsrjpAs8LW+y92zHpXicsLQOoGMJM
nUInNKSVFFBnAO5cjzaLiUR5WFuWa8Pd2oxhBE3K5mw2/5YHvZhA7Msuw+3SSJ+I7vkckV9SDPCM
vH3/OR1AgAvbr3piz3ym6H4kaz95tNDUQuz+HtJEv5hprEEaimYfsYdrn+d1kj95nsbop2bwdPJ6
BPYVjvVFTr2zRJyxLcuK1g5LjG8QWNNt8Qkc7NnMXTtkbw0K9sToZgQQaN3JZbvz+JiZC7KDbw8f
GMu2UCskBJtEjRj3hO2esv6+VcBLTXxTdG0C6q8VwDiImthNE6sxlbyqzDcJKHIfJAM20NojGUEE
g0sx+BKh9UUcrLZ6re5ELTmFuYUW6JzeqPIx1eizc0c0YUbdzau7D8FBzt+FP6E2XSqatNyi6uin
ztodhv0RomGYIg1PS7L5bTu9iKLXh3pwe6mabUJzUTGPmLLD+wpRRpz5LriLqbPd6gfCCcZCE4JW
cKKEvxbcWABGZQirWoIwm/nM1fzcyvG2Z2AVvJLkDjClcw0r1zJFzKPGhYYPlrU2c8jKJw5Kr4iB
Ss9MYQEtNjW5xni/4HC0QtjF9fxvOsIWtWZT57Oi6+qn5tXnzM5vuHX8zUiEsIgF4pIzzPFJMDLb
ANyAvBhPh/mm9CtKO2vWMbVNO2aAGvRBYyED37BJYRqaPl/1yuiadMRlQLWW/GBkprXEfOiti4/e
S4p2Oq38msw4h2x/cNTB4WC3aS/XB/1oMmt5M2YuDLBPtVrIYnj2MnqkW2/H43u0ZVFOMEuP2yOa
60qD2kitwu1yw2wrD1oLlrkCAmmYQ2FuL5h/WI8UgfwqfVTBsK2mUnQ/UffnPUQsGCZw4WdMYBNl
/wUibg4ur34T/vyui7JT/103UyndiWlFW0P5kNgjrCAUqXEvjhu3GTK4hKBZRhhiRf1pOE4EEQWj
1uecLd/3w1trLnwfl1W82qYcpLhgmT6iKvZTqBTsXCER/MbeGPLeJLCbHFhQPrHj/yj36w+xWqpR
ZDfzdUj5dGkZanI8DUJTDK2WlyRI1Qor1jB4Ql/y6VmfcAhy86ILsn9TgI21RKGplY7xvZk4s6uf
7xZi4YrjKhwckYAfCdhKsmu1QaQzWAFFSIJyJDrGHm/SHrUGuCOHt5JrkLk3kZ1M777nF0GTd17T
sgr27oynJ/Pc6E6BvZ+zCwJ5jRWgOj5oRJua14ZLhys2w67FoXk+39xucw1yPXL85T6BDRgsVIZo
8G9YVQWeeGxmikm6tbewwS+gSDXMbOa3yjntnuuUmmO6QYr6S4VDs0thrQhmg1Y31L4Idbhpgnx5
G2c+IDjtHpv6kvKEM5kUbxcufCbYv8CTEpAOZsjxqVLsTk8xWWvxoUwGRLxxOP98hkreefNyppmq
VveRapbBrJgCF49D2X5gdKAFa3Mu/2avWI74ppwUMyG6MRZ5iTt5aG/ghZeDmyubgdo+zN5akwML
izv7nhMOQAflvO8tVBsmerxxXASz+v3YAcdE0O4MD2+XSGjCu/UeSYuZDDVTOaEYIyU42Rb/bW/L
M/m5zB62in5GOLXorMuN8rW9nD4+ryLzsNwjldZyWcE/8RR3RQHATlsA9VVkSM6cCZrAP+ALMzRP
qoZXQsEq7SLmaWVMjHlkeRAZX2q69f+JwRYZsFLaoHGtSd7W8r1gChHwYuV9CGzWSJEPko5m//73
BeGf3a4cK8bzvt/9OtWgUvL9xMGBjRHG+C0+MmMWv4X+De7NpVD9jchEft9FRAOe3c38n8tYbv7Q
RE8VsI/GptLXQQv05xGq5Xo4W0aR4Ec+p1KGorYxU5XjJEPL4jwerXzEBYQfgQ4Bll/tBE+3Xus8
LTpEDeREDBnhtv1v3Z9JFSg7kVJpxwX8DqARvc4SgJt5qZJRA5c7lD9xB44kUELyOoxj1As+gVvW
cMizHi0Ed8IXrhe6eVQmTFA9j6fyKrW8vQBkTYEBkD42ZBeq2R35wqJDuPlMO6h7St/mepDFfB3D
rwNOpOQ80dhwXOGowBxoKsSuewoVmxPKk8YG1FmNLdbcTqTNb3edb3wFD34X4tp6hiNu8Yq6HzV6
ZvT1swOYdiIt1mdKOFMtnn+jKvu2cwhLMEZx2sFWff4nwfEZABxSoYaxXwDu6lVPygnmSJIm1vSi
oIUxO0JkJnMJtsEdFMl7Dw0C5LVDA5p/fdDUDKngeB+58Mq0QqWZSSGP4AOQ+sca8WZEbHevlGHN
sKuAPbJwJ4g3XxyclP6neZW0SgPZck6EQJTYT6maVEQ2u0NpWU2jgn5bkFa4kTNIem1MCJNKm6Bu
JtylIcutbnVDfuLu+mNDh/j/ZoqLQyzAMcc7PSWvJPXpe1NoAAEPkzgVvu2rJjzK4NfW1NR5/Rkw
XRPrE9Y1SITkfePqL1AVv1IcxxtzFYY5+75RFZsj/WS0iD6MZATwFygLzS4py/4rU4s2inuFxjWE
Tmt/2laAEeRurhU0sA8wO/M3YkdkB6GmXVAI8ds4ed9xxHaTcdiSOQq605+0LlJqzEYak+kx4GBa
KcZbxw6abl3i7LUNLCa75lN1Hx00i1dcZL53f+zWciPEq1ojJ9jQ+OUivKhr+/+5hQscxLenzEOQ
koPou2SBusfyLd2iql1EuufpbhmUVEvZjyuNG4xrxFy/am3U0VlRVLqKPhTEDxXC3q4q6/VDZmDY
fHozppEEXpR6864SDfQI3cQfALYE1u8eet47h7duEOoXzHDKUoMzLgAs4p3ye7bvYGIkfiJvAzwu
vZKJaB0039gFvparZmbt9Qr9dKgjhun///fZc3HlQDmGQ7nlwLW2BOmNhtEKv2Fk+H1HsgVYHY/B
Rdv4OXO4bCn2fwogaJtaJ/vz0EHZif/Gy5au0nK35no8+/XTA+bO+bXsQbCuReYRkmdV1n1oDK0Q
abS2+pKeVqGpNSe73FLCXxIK8XvF3LVai6N6w0NF9cpQ95DzP/IQGnrzod/nJNC1tuzJaQj1nVAS
s6+wM36GgSFgsXBdra0gfXqOU6/SmjrAsenUmAeY+4+HqWpF/mu3MJjJ32hdHRlKMB/corMKk8qd
y2rml7jHQ7z+NuI9OHuNo/NhrhYXiqqz9gaomf2BwpIBy1vfeHXXsuJ1KnXflhc2mPYFhawksCns
H4ZHQfUjYdaopyc0NTFIOjSGLZJVGmJZNYdHkaYGRAQ+QQkTeeC2jN7pBCJ8gXW75uYbF9JN6DNj
govFG75PZOFP4Kovs9JyaR08h/xnYm0B9MKHF9QqAFZOtGYudLM/wcKf/H1H4TXv2ukyJaW1unVE
NxXN0XjLVDOc546+yzP0PC+F21W8Fk+8bHHHoymnCwheOXENLSXzQ8O/GbzfTelhTfzNRj7NwHdo
+QtYLPYyEB/04ZSxF1JE36uRtuOyZ/sy4NFfi1ypImC8lLuBWhs7A3JPTSeyS9VxITbLtcCd0vt/
hd4dC2m4uDbCsn7J7/uJkGkBRcsLiRH5ExK8c53Bq5vp0raFzZflVYlxmWDnVtco391pPxflXWQ9
s8JSOQakVBSdEugUT9zfn3xM8d+T+lYqonHyaAJM45U13JxJGJWKgRC/4Dr/4eW9Tsv//ZNbdRku
tUcCTnmOxMtVHfXpcVPYGe+5oZ0zbIhRQfZ8LwgRjRzi7ywtIzpfDMr0+Fvehblh+B8loXVjANz5
LEwAXJT9G7LwWcatc+3F8vrezL/lJ/8mg5CpzsI0gR04JXljDbCThN0Oy16ygGfQQJAUS6nX+4fG
1xf5Tpudch1wFS1fF07o0RzLao2p9uw21fAZmOrpWfBKrUZGj4OSRSjSjb+Dj9TfRlOPjlfQ4tot
FfE3hkjl5/gfQY7shPa0MAjPP73eqZUwL47Gw89fcsatzLbHYs+M9nCzQNzK8wlRUqH5bYK8HTKf
ewRh9V9/B7kMyVzMlJwubIsZjotum5w1uu0HprRH/2g4piGPtWe1C8zPUIUQnylI6ihpApwei7dG
DwFHLVXfvwKeSdXMi20ZxPc4Dx5NmFt+/Lg7u0OPevpq8/01hT0kSgYr4nQpBuVgXMA9A+DL/5VD
X63iKIJXg7bGQUhZtsZLEhsccDtYyO7kCh7N5jyulJc+SWTjlBTA0ham0B7s7w+PvgHe/MjhOGo6
8PGV5Pe5oeaV+brEsjk9C/Azbe+b525dxFOMY4teHhrkuFpQU6RrHhTOBXsJpO7+wA8A8ygpx5hl
EMa0Fl1LidXgxNKtiSVF7csEBLJD/ZoVXJzlQCuk+fMw8SyNV2OKfarwrC1jHSQKmUMENXY/hEh9
x4A3iu1V0Na4wxvVld3RforbQDk0ubkvhaLpH5BGoP2JjpcuAMCtJIsdz7MgoSGAYc9Uqxvm2cZ/
51buOsFh+fZaRVocZrEXdfl0zOF2dC8iHpK4QchL+21G/lbbX3XnuYRT8ZY9RA1NaCWxDGETdGZV
4NVAoqz2YvdgkJb3HYoRAGx0L6AGySDLgmF0TzO/n4cBqOq9NmI7hKhYdasCAe4CaysxfqP5zSgT
gu+Ftk/RD3tTxBpr4ItVAUP0IF2gIhCtS5/2sV9s/taJ6x5HU733oKOBnGYe+4+7hmeLLyztwkV6
DlLbuGQVi2WHhvDk8iuU6cK6KJTc8QeK2o1tmPiqH46+tHUwvHG+Bp21KB+l+janeTsDoTH3zSTT
zJUj/GJAp4yuZ5beFchGbJcngLQ9FZr4VBKBTmSfR3r2WEksrLVT8mTXx9xkXo78F1EjLZlyfG5G
0GrR+8VcvmYhV+ke+F1DhyI4m7H/BfVdf78Z0vcXTx/emR/JLEjuI9RlYfEsW9tJ87TTJ4/O3Ixu
DoUWbn0F1/5569QBxpaS1k+wDLQkwRGLbgewGUSOVijjt9RlZ8yYft9Vp1kyQ5ZX/oYx7C4FlKbU
4n6LjQUsa5hxtr9VpR6GNrh+xwzXX9xKeGEjL1We3u/NLDtCuyrIQvu0wYEz1xMWC1+s/9ASRGaO
ehYO3K4lT5vqS8LQBm0YrZttxTPunx6JDmHVEH/91zQDrgyZHObuAK4FE5va2WFyRb7jw/Fi2R0Z
ZZHTBU26IzYwqHIyVrmidF+wa3rOXYCbrSa5bFvujLlX0KaEdbw9w1iNqxj+ojbO+B/C0AOlqiWa
D8yqQWxaMUuuSbo94cQCpTtZq1AQeBew3BFbUUdHuLZo9sJrGAh6fJpbttFXk4syJi6Geq7Lpcs9
VVGn/ycR06VKfdPVCjbEg6mQp5/8o+/puR1qNd7sWnopjNc3q9kfV4YBgVhYouJN/rF4nCMCrGU2
wPkWoagTHybdBqqVDeUaABaHy0Mler/sIJjVJ9LUstCMMhlfvjgdA+w1xhiYH5LMDEnn+8/HvGsn
tgbrcWhMKaUZgiyrLynD8eWjEXsaEYXieNN70MDdsOcG8c7vfypsGWiER4Cx11/RJw3/uN4H1f7c
TXfJhv7YLVCYpD7WkkaSyka6wMgycA7TQvjgPqG1WZavTs3WygrhRkOlHE57SFjcg0h1cmbS1e1p
s6epGTNeRozdt7OnrLmFVj2ACxEtwG39/c+5KtFd3vXA8M2EsPRM7t9IA/7W/uEJme7T3NpcDUpq
Akm8d1ERkKGvEO5/B9xCYMEOWxzsBowdrDDadlN8CgNr6ze2hYrPvjgSkN8BHu57C4L6YUqrBzqf
aJU6sn3fL9QsNmv+uNbLHvgy55Ut074hcSRGDgJ37ED4bCAZMlkNFh0JogTyk2P4D6J9f8l/fb0D
HmftcOMvCJIH7RqHjsrEKrYUtqMqTkc2WCGi5iyX0ueyxFurFB9RPiyXrdPhb4Iqccq6a3XbHnHm
rMyuhKcex90pf00r1X+rr6HSBRuI17BxmwHCCuH1h3M6BIrHy0K3EP8qGD/A2+XkwGxu9jwxppLF
hoWZvps+On0/gjoFU23bZQlSZgdkkBmrdtRrxbs5u69oQvbQ3hG7PkqTJvJGMnOur6GCtoJ+wE0b
HkeV1L5NSrl862JZbvTaoSivnJfm6frXQGQ26dmQ1Qpuc594xYzsi0dlt+UNa3CPg7iwfseYel1W
iI6KDcFDr6iQTDvDRlD2TldyhjSAUddwT3ki50LDEcTm6k+jH5+qgX6EwXLkz8xvh+JbKS0pZ5v9
DUyuvmmzZe89scv27LAKCl3GSvLbVU9U0uwpkDUIyZKsvnG3H/F8e0LRtwSb3Pg2B1n/leXucqbE
qeOypALa1t8EF+l2z6h699kamYWnxz+Z8xIZBWwgqC64hvk9LIwxaAqlSNd+nlP+ze0B4MZNn1/w
/eggZSY4tRq4ump0PDryTeNxIKoVsp/F8rR7aYUOovDjjI66uP/ccRx6Rsu70T/JakOk5ilp4mt8
brpyXOW8FgjpZkvgpTi3rKXODWEtr+t4L2Pk5EwreNqVwquk5qj0apCOcXLRCi0PVdr/0FRez0EZ
yV2j/tGhzavpSGyp3nj1fBUbfLql9qDSx5Kj3EAWQHQaFH6PQY9W/DwWyYqngLST67OGkVxpoyAw
qkkWxGiKJLq15n493Cu9zBqF4fv9LLm7qZlu3TNo9dqMxajqUJZ30qBvoOkYXzbbERVxuTyxZ6K8
vo5AdKjGqbgX3s6NXp/2t4/pSNI7Ka54HRueVJCn1Q6pjINg7ysaIc+DpGX+5UI96D0uCFieVSzN
uFmLGgW+nHc8TGuJ1LTG1OTXOHbGXcW38xuebryVRYpQsepcLuRFx7qfZXJZNMJ3dz2bZrATjxMP
81WPmt2xwClz0Zj61dG4O8OA12B+V5GnV0rekEu+D2Y8qNU4I2E227q13RtI0OGKLfGHkBt8CRMy
x8wtcx2yle+lIfIZ6wviN+ORvp+q32Yoq5v5V6tsQk80yTZvpCEAatFtmHqD1YYuNwWxR0496raV
fu7q/yfCflH+dustTxgKdqB+GR3KsHbxKpU1KemA20IL8TcTUAzb58JXZC4dx4mxPydBM+Zct5aM
FReedm+XzqNAO29ZsyrrkEiZ1zq70IWP/25BxhUhmfP2U3lIF6zKt9g1Qf+zfjAuLCi5AFXB3uvm
eHemV6vqaavhwYORhphAUaaoWj+nnm0ajPLekIYijAACTcCKppGXAnKG0w38auadJ5+grx3Bd7ui
ziIJsVrpFMmLVE+f+fbIpX82Ayn3yAG5KRGnk0eNR3StEiKQ4l3dZik7BPdm7sPxS38GQ2kLUqVL
XvqnRAuoClbs1Odn8b9lIiEq7ADbXSXoNCWc5+TMy9ZsNsRpZJytXTrq24p128WXaWAuExZ/RcMy
OFSam+iEiTSX/yTwHaqElGdlcedbANx151J1ASKhrhfLd2qTb1jkK0uoH9xpaTK+RyfgtVXjbCNr
XEMnBMBHSrIVVuTkp17C57IEkUHJljNN6+C+IZPz0zE/yomJU4cYO3xZ4zYNG0P58zcqAeH0BN1u
JGXtb0ZuaYibIafzPTWyFG2GsLQakAuQxnab+f4xCqKBbiJQ5OaE9cI0mcreB3XWILPyFo6YUBcu
KeFdH5MBfl5DuIdhJG5upBnogtovNPH2qvD7Zar3jA6nZIcLVhFts6ujoP9t4RLWGY2rviAcKoD7
GQsR0lPB6A2LsySLlyNTRgBwt+iXB0wZT92MxzX7pTaYgPX/vbghUdm+j8iasyQxN8ZBPYZ5/ze6
PGzf/7NQQ2vTOXarq9g7PDZn+mBdQkHKeVXtllafE9JffTqx4O9gzTpdMjmGOy22pKJ/AT/OptCI
rN02o7uqTstlqQKVhelYSd02hg+xx8dDd8b1oh5zj6S9uHj9rSyHeOHxFXAbEx1sYKCIH1MkU3xL
5YIQvRdwThHB0cXCp4V5nfKOt+zC+Ds3uHIPl+c4hzqz1EOALzasFz/p57W2Pnox8QVo/LDIX6+a
FnKeDTsaGMn+SF3N99n/N1m4cx3hmNbxPqhjh9Py4b+Tdnl+SEYi/NxP42ib9geu3UsU8P37jjb+
ni/lAS4MeAtHPIBT473hHg4MVFDMv2DfSg/NlcLQh3cTjbYjQ5vM7iVXRQwZ9oKZTT8o9vz2WEjV
LdeFNaBQ+xEMi3D4bfmJP0GLqQ3t1hKuZJIGLnN3yFp97S5FiKxbdMZVwXfsRTSNz1xab/rtDvG6
box5HC7hENqXqm07/WEzF1eCSYlGBVGYWEvs1EjDRr58jenFnKXDI/yZmyiisD4+JTMLr3zoY8RW
HcspPTkEAEWu2xG9DYgONDGQk9bDc+y4ZVhoaU1e0WAl0tTEPMFwKXVadNX/lddnkSaa93vDMFw9
gEVn1JlPa1aTa0BRiqdzzOTKXa3MyR2E0Cxlc7oDIytc+ofgLGy8QNEt0tKrKZNeLIUKPcHesyov
/Bx9n3/2LgssEAqW4Zs12u2nSjt5v+3btRLi8pmCk/2GnbpoybamNSdpjQUEsaM8XwLYhI2SvES+
bfWBq6YHs54eCKJrsETKrxkl/pdyMDialxvhXDUKdz2GH0nx/tNwwljo5ohOIPxW6+Cc4n0mfLhQ
UXOiGfOCXq8zu5ISb6GXo0WYlmx+MlrCYCtBbsZCLebmDM3VD+u0IC80gAXxBx+CZ6kap8pIa56g
AF372biIEAp6rpWVB3nPnwPXEj7tizAN8cYA8n87GwlydPazI6h4AdS7eBYtLLxhs054HaskvmQC
KmkZQrQREAvkxhUa6plpHBN52y8guO06q2wFjXraDAgbSCTCaQSqgq0Rb2sjU/b3B6k4cUB2qPYD
kKryf45a16koo9WxABY4zGmeDAsaW2j/qrehAAbf1ui11HWbfQyiuMdFnPZ4aEVodktomUgmDh7M
iVxDnHLvOwOrBVQ8FK/HryVXmZ3sayYZdVOFJWDrcRer0JO9rdcNzxb3Ob51XdC5CivDweXovCuE
4w+KCx14zmWEi1PyKsygcE7qewfsX2gLt2CH/qzX6PgNqMWnWrgzOXzgDGsaVN4jyAzfjzswdYe+
4vrSSXnyFvLyskp6gk/vV4Op2ApUwRo3xK4jvTznsqyIexF79v5WGfiZ5BNP/T2H6wix0Oo8WtDh
QApx8X6OwHCKNcIae9pLxGKL89SUAI4UGjjclO8HaFWpCGczxBNOWSZnaznihMCkMdP3tHDKh3Sa
NeAycdCZ/XqlU9pfKeuJfwhkEoM6a3I1Y0jvcqE8c7bPAjVumAhhKtojC9X5Yz3VPg6dZzKszTVk
Rrd9DFmmlFSFo381Z2y5ODjV2+LEZkXJKTSzbGd/Jt/xDFedLwtCQ71rPWYT7f05CbBY4dachVNU
3KbtIeZB2FVgfWdqpiFzRi1BfAQw/5FjmKLljKYwQAMbhD0/vAZC56+nckoxzdIEt7z8OToGkMFE
6cKnLqvdh//VhIMgxbZxU8EiiKd5+v0cesFMzzlc+qmd5Tk90hfsAcXImrlF0Iqu2h+37slzDhIC
64y8pWpB2zHi9V96DuRY5e6/1BT4dBK+6uA1745Ngpe+vn8ruPyxB/kuRkONqm50PFwfqaKvIlnb
AiQybn9tKkJjTsZ3fg1eprB6Ge46YXmEPgf9yKZwaEALjyvxksyGZzDwkub99zDcLZjWeZaL7gB4
7UyF4I6ANztMMDDzJK17hwX8xoJTeAyKXGLdnTOqJOgbrozx3A7Ib+gkZKZ5yg+e2kIbkGEVnrqy
SoYK7qdGl5xBoCTLBzbAHOcjVaDWHalPwZTyTNCHfsFvOTh5GWE2dlZCkc8w/V+FmPr3UFdTWC/r
ExSYDtcyzgDFAxgXfH48UbMjCDFIM4rfSbXONzNXiaLOBZY+WdkstQ0KzxsEcbaHeWNLzqugjhEK
NwjUF6ciwwiAMZvn61wSy9QZyDTe9eNWL7s9g2OCHfMWEPPD9cZWKPCVUxgWlOxPzRPX8q7RsSKq
8qHThg0eQYymxdjQQs+nbGvI27RkSWqxRKDOFC3/5/jwZLVaEJa+T6UEDdz5BvxBvs9BQ0jVoXH1
6Zwky4vkqpTtSRJd69m5/WzNucmXUh9ScWrLn4ulqVoZWtrW4XsEtoPWlwY3HRHx9XMPrMpBgEKq
t8dcgcSnxlOlCVl9J5ZCb7N9nwNWzn9lPrGzsL8ra8Wi4bKVtYXPNP8zEUYoJqfb/wPqkO2wMExG
+ffklIFZofCYb0ZsusgSfr+6S39NnT9hmMgTxo83HNIs28FZSyibq/+a8Uags7gg92yjv5ieZ7Sj
IwzzMC5ieoL5nuoz23MugokqQJxfNNYwRX6DnLtGzXD6+yiEGYmI+Aa1jgiaPgSgAViWCdk7h43z
lT2+iSoP2ZmNzqYKIWDx2+MpxRBIm2+y/mH6wWJK+PZ/BdDyXFTE/c9NzDNFMjNU+DQEY23TJR9j
Yws4KsknxIo8DTfKaxoAaZar5TfF1GYe6+A99kQ4Mu/SU68//YEEf+cuUvYmCmBgqPu3CtliTUvE
NIUFwuu4cn/PPfFN79GBKQfkyHzcacDYsYawEfbE2AV8uEKZcb/Sp4m8s2qL9IcesKZnVJyLKYKX
zAHyrsuOMI7KxRGAu3s/ev0qxWW2tyRkrOo6SskDxTEJTDlgtfc0QJ8E8g5rg1Zxe6BY2sCQIDLP
IDPiHhxdeD4W3tqAShlbZUl0kgfxAJk/TU889YiRzO+0UqsNlUjK34A+ssK2qsy2xPu02xX7RF3m
7/zCjAoap4jljyUyEBlIjG+ZXqD6mKvo6OcCgCaGKMjxjxIYPx7Ep1fkTfq6tz+zRoP/sKPfln0z
YVYUl6+k272NadeFbHCNDkHUncn4G0fHJWzM+45zlCvu8cSz2zzo3TJfJQgoKkp3fZRFruY7WkOj
mPSGtcRQVQRdj2HvtZn2ERmGTYdKOWnbpwBwmh0cPx1bLKnd9gfmLCdPtog9sSZu9txX8x4VqT32
iA3PGFtDzBxlMvynLz1VSRilyrO/sRLLZbLv4PkE8GOhxL16afoyvSiDFdxRerrYM+VQ5dupyyKb
jrmgwfMoaMl6HR0jo+V9Y33DvGG1OBan9cD59USuKwldsnUXDzkSrrNHunDmL8QAGByWXqKS4HeX
cS2fxAnUH1c40ZbTBFIYKkRWziJ/7tzhjSR8Mg5e7BmW0QC7EBrIQGiulmUDdDfPpidGPxvBHsfy
HUfHIneeX4QGyQgfViHCc3zbbr0h2xQ5LhqM0Z7UJVrtuwfbJXyWILPiC0N8vmDDsJUObJqNF3MM
vCc0F3xYwxtEkK/ACpfP4hzXZ+01AHPXFtyNVDho/gpgZIL1l3wU7cNUkT571cJ2U5oerNS93os2
uziGIFVbvkXdGgN2k0gBeguAWkJEbe6uurSYwAcUTNLkyMNd8uV5cw+euZNZzcqHMcpmrN+5kLWw
wzWewu056l9rPYPHOe/naaoFsfAArxRQvGoNy/uyuviSsTTg0SfgvPK73oW9WAxQ7Jy8acgM3K8N
/Iko+9ktOwSVg8gCbjEIjl68NFb5EJAbLfv3ixS1DtliUDtvRhDoUNhTRy59lvLRQuTnjK8GGbca
u/Qi9Asdi19DKJW+7TJmSSmYbGN9U4jPI7teyyq0T1HLmGvQNZ0PSreijfxomAAq7TabkRbU5l2i
1kqQ+hcunHWGFtEMy2jXHtmM72hRpu8KEC3X9dzvDANfW5ycRODfi+IwCxraMzYSACMjo32rSWTE
bk/U4ZKvLx4rvviJYsQBCT9lJXkSCKIN0tIy0mv4vOARK26b1x1QPJs5gM0GZAz3MStNlGWNtppx
xK/MJ+XFDkThC1tMyvt4T5/4jRtlNfYvMmYuEEVH1jx2tAZC3PYREfoSXYMuvbGBzjaj4OUuJwOb
HFTtoCkb6hMTc0JiOhbZsi9wWwpYizz8vvGmc3eIxb6EhV/ccW8sDHNiZafK9SwvUOluQOYrDAzM
waZ7j+fmgoXAPeB7c7FCLNFwNi2iZfPPOiwI3nW7f92F2w+0j9caM9auB+eLd6DGZtbiUyeCqdkL
WLOoBBrbDIvMiJFOsftFAL1k/pN0pX/Y9Zb8lX4JUYov2e0P5g1zDhLqfgofrrTh7oCY+6pRGjdU
ndcpHdddvlz1YsC/tPsGCRULDrh1E5ZaNRRIeCz+XrUMLpc+SkNmO8tELOVUbLJl0PMjclJznPim
VdK9OBP0WMpXGlL+5tvV0cuGouzN9AzcP8U6lyKVLcvcMIDvzQZZZVdMjoj0rwndPNevSoy/5bK2
ydqEOk+1JtA3sfwW+WrRkJVwPkNneNkV6T25KiZKlDlwRzHLbO2RCTlADlYjk1T3XdrkAXz7HsXO
AC85PmXep+t1SaZ3lH+6lm7roPrxP4oyx21nZIPPkPmQOToFD8XKfVAEwqdE1mBb9d1CtesTCg5R
IVo0+ReRj378uR8YgJjYufO1qQco1jnhDXT5ImOlAs7QAhgoXpvJ5/IWTfWNqkHqLGc6vhJB2duD
7voXozABvcLuw/eoS1RnH1Kwmj+0+H0Jf91/fSZraH/mRHjLWvT9S6sGGq+5JjM5Bz4l23kqX2Kv
NpDsRaQ63h4hkz/57IQJDy8Ez85OuOI1Xc0ztbMFh16aVmL7ymFDWaG49LH1ASIV1be/VRBCdljU
/Mu9hJhipMG2RXEg98rTtHwx7Lp2SBBYtoj7/GmrVeeX4Bsn47cKB2iLnys+cJnp5B6pzBa/3Ty5
KPjS+vVZ+yDbAT141P5MZoPkXW3UZWlxDbbpytvqqSECZLnuzSkH/2fwYxFMO1jzZmIAp0/xvx6+
FKiwgAZ1rtGwo962KqlWZNnYO/O+dTCWvKAr6K6B8u+9jGbZ42SNRsghtNdvD3UIQSLZXtiENfOu
mPnpc9JGdbMziP88ZCa+AtHc1m99goIP0n7FZOFIGx46ba4O69xYE9VOBPqQemmNfQy4Qr5yHYDx
WPeZIYDbIXFp7Pm113NlLEu4+yD6cxIRhicFBC/syQjqJX7Ta1A9wwqCmhxOEG8RiDG0pjPI1g9g
iOdGRTXlGOnwbtDme/iVmyfT6skHhVP28UVUz8NHmXkm/IVROH+iCYe56jlU590i/RK3snzz4O4s
XUm95yBcXRSgLdw20A/vQ+abNS323pSO2Hc4s0EeCiBHsxaqmuFo2+SK7CzXlZrvpn+gS2qEGgWX
0raOR9c5TuCoCHpVfnG9qi5kuSIhaqiF+oblJXoBEeG1BOWvN0p1nFdmCZd1yxgNeZ8CRVHivht6
iPCpx1ddL/bABXZcIfZJO8/cMX3q5/qyhGnPeGeeCjvVTJ4eIFljCGtk1OLb4UxiZNfwQfT+0czY
MoJ3Z9QofCZsvVy1JW858797UL1S9BhkJiJKITdGgPhokwhK2tixIOul4m1Hor+BNM4oEsT5T1fX
VyNzcv1q+vKtcyK/9/sWWvAS/PTm/SPioTJm+R6PiEkSFkFikISWa+FD3fm81sbIDN/lCHxbXCmU
k71xaE3ngwnlC5uFidVu02BsrNFodR23fpGh1kWiHaEtAbqPqVEqnoRqlYcQyPUdvyf3gMm4RqMW
eXQw24vuZDoAHUa36VTswdSS9DgJ64xUv6LFmHDlnHf4p+SIMg4LnbeQf1AQsAv18Ui6pX057oqz
u8+3mu6uX2W82jSCl14bezKgGzkkKkdxZXF0FjHYWLib7/7aQNYuzfqbg9AQHpcsHUy5i+P7aKUD
Pj1M+oQesGQ+HiK/db/JlCH1XWc7Ub9Wb0S3/R2J6mF8mifyt9ryoDqKhnqtFchEytBHTNxPDTgs
++SmkvXhOC3juZFXX0v6ybqsxmdueIfjiUlDngF6AeMhpNz1M2DnBIi5yr+OSvsDOf5Z2ZeZT2fl
YdZKIScc+CFtBRAN//y1RImqsE6CI7+7Ozj2bAe+KMdHu0+byQTV2ndNwAtEypcoxkx1H8czUbyK
Ujhwwf3AsIR7tAcBrA7fPSKLmWJ5kzc/NTaYFb49G755+q7PBoCvPb9Mkiub5wn0u0IFfy3e/Qyl
yq+akQlFKpwCgmdBExObXFuyymST+dwN5uJrLpalj02Eu2bQ37eJm+m7JoP748gxapKvJ6EdZd3K
yUbtVJQw4IqBb+oXdjy78WA71q5t9YMZB3L2XIXmwrMrVp0uHOFC6J2AwlDthEEnAzMC26XZOSBh
CKQKhJACyw4Ajqrw4fKIdbGjaIP/FE+gW7qjMkjFlYWG9gB31bENSuGFL+EZV8YspYxANsR9nNBA
hkJ3lSqLxs84nAV4yziMn6IyPxPGliF/DTPwDXr7rt2u9ZBoRZdzaaZ+wJig8N+c248gj6HDUq0L
Pe4hteSsAG3CuC2gMNb3aDWhNS2TAWum03hxTM8OFCC8uuMMpbhzMuVZXiqwmPHCidGd/UpdftTf
LxkvBKJRBFEiRWbDg8KrrGASIOeZJWBVusWNT9vSJbTgF2+NILPtCZhcqR4FR03uA27nNMx4BT4S
rLF3Rp7USb59Skn9WPl18Blz9+fzXvBMRZ5RztWWpyJizOiRkYdOAuoXKB7jrS9UHGKIl5pQXV42
B36sdmxOrpJia9e8xIeduX+2dK+CL36qO8hLUJbW558BKyJEItV2fmICQldS3mh1bvPG2zMel/iA
Plzn5DXQhYWNF/Lwkha+A9Re9s0twsSVSS4vHarHLpJ8n1tI8+lD3ovtMbBhx8a5++UMT4P7dWRf
wv9Nn8xeUc96lW4w0krVOJbd3oK8NwWHPAX2oJTbPxgohPKONQ2SS5mQC0MBdGNrOwbGK3tapBkG
aX+Zf2A9pp5O58AFfIscnvjLV7PCtvcidso54EFdNuovwbmr78DjQgsx6xpqbwO5jfwRaggnqL/k
TolrA6sNJka1GMXPqdCu6p5SVNGFTvxXlZKXKso520HhGNkGvOhD/p2vVhdn2/Lb56bfkacWpwdO
UdMz+Y8qJPBj7RUiHkCdpQkkmq/UMIhppDz6GfLIp9P7lWOdaBJUrIepodq5n1ue96ll/BgvVp6D
uBhioxFoJ+N3x2EVmrITz2bI7/Ow73YxosBEpPsjgcC7f/TpubVk5nNtLnZJqCt0MMebzqV7w9HZ
FxmMZm2wGjO4f+K3W+p1tljXrqESFZ9PSwo8PBE0ukOpAHoenmS+cZ7qrjCLJ0ZckWDj1YOCtWXY
K4mNaktmHx/lBxS105M26S/3K6A5szXEKMuIw/SlILTUZR42SLuhpUiTgOmpSnd8oJkru9qsaqcs
d5zkxiXbM+OOhBkVX6bgUKuYDEl8dQq3uJ9fMGSg1voUOVvBv/rxSpS3SQDM9b8OpfnR+lPJAk3G
6ujEwjPCANNSPCqVBVOTqrOOPvM0oXnUOvd6IPk5UvGmUez3sPsySF1RTRbMKtxuMSxoLWEJJzaA
c9/7M43yKn/a1qTo5tsF8GzImITnj9kn5CFht9NnbUh24JxT1hVRctaLvVB/r/omQaCs+PID83YQ
2He2DC9qpV7VRczzC71/oS9C29Qnop3+mJip7856U2MrAz0ksTAl1dqe+Fa8bNqx/olrcMSJ3sQ+
4oSjqXAUnvqhCRBkOjrdW77l7OyGYzqqXxwG2j5LxiIYiioUQZnwcYx2jLHXazUU1HXvggvLo7J6
8H9wDZrmoWxRmVSBvEEndvAuJwAgZGwhElpbi5QTCHn17yeimEJ79CaaNnEa2aSrbMTXNLrQFsTh
SMfepHCwrYAqrW79JA666IZA7dypv3797YWZKpaWM425PD4QFcDf/apx+MMROcynTHMoKIcVgCq4
f1J+4ilOyq5slYqzxvmcC3D+MSZPLbmD8IMPtrFgL6lLCFRGf7ycMwSqKtoN910dheTKhE+gsUhC
CTrQ2pCbXmchVPZonOw0j0rZa2tkjphvjYwdVfp9kVJZ3krmj2exFYYExMctR9Yhb6w0MRHwbsER
MItSQYf2NvkcbHRPfzEC/Zfm9rBxNCVJ10hAMBtLH+ars7qCTP9kiEWmHdYs+WizpioypfEDxquK
PUajIe9zaaXc8lGoRDVCbUqi/Fr47d2R67bv2FUQGRHy3mXN1AFMVXDOU2l/Pe7oTJyefFBPtrUS
RGbOYecH0aeu3wV8m1ptPl0YOME98Rn7HQ6kxDMAfoDFmhxGhuix381XWDgWFeegmWr6NtYrmsB+
Mo26e1PLX0tfWHCWvkLCkh6sRLSdIwy8iWBXS+jNo6IDi8dYAooUZdVwDlF/SAySpRNpG2Iv1kQE
qrms27sh0IlbdjNpXEEFtFDdZESx+F7BKisf8/+3imnZrA3Z4aLmEbZdyalgHZSEYoagdhZhB5jD
T7adFImyI2XEwLQ5x6vgR6z5fbD7RstNPjg1M8Q3zwkGNq2/d1vKOHhN4Qbmf7BbhYWvX5jtkayP
o3Ot6ve+WdVs244Jkg8I0CIW1Evl3wGb7T+O6y5UvIBpKGsxceeRsd7U8N2A0dIYIQAb2zEfH6A/
axJk88Uyuw0UM91DDUTDeTpPTJ9obIJBAtsZtv7W8woozasV7zRxClq895Z38u5kLS1MLsN+YOr1
sZK+DiaH6qxSfRlY+0B4cD2BS5c/seaX1K8/dIe1Z1ce9QL6xlKoM6sVdOx9pb4i+iufCV9W31P/
BeyWUjliUixPgMDok9nmB7EcF8BU5OeC9vUlZvsWoYO3XESmhDWZhwk5mcNr0yE9bUW2/k5llrxJ
Y00c8gDznK90GDFdKkcMyhdK8UXmzF8P07stiElgDcYteyTUaqeYuv9t0mMXXeOw0Kjsy3ofmh1h
D4SBnpPXebUsTsutdSZUQ+uvOycbSDt2LH9mpsF/l8YZCcSmC60A2YGSZK3vGiGv8Gcme8QoRMTU
yf/QT/k1BgS9D0XS4XRURCPTOtwv0L26FtzvlIny2xUlUK2dLySwbzigp1elmfZJMZ0y2uNfAlmH
aLa4/tzyjAuy6ZSjyZpIkxidDJ8AezovjGpaFn6HOFrOYSK+I9y74Wc9aDrnVYKCg9FOkCCU2lEO
py/DIxUxoxtNkvp2QecD7Km4j9YPYfkp6jg0+7BsfEzFZfpkGLsppd9dkiM2nEHdX4oVwEmdmOqu
y7lkuL0BWL+RcXbQptNRAoIWvpOi/ignL/Io7ZySEjMSncGsfQKB5NNxvMkZE+u3Gu/WWMlzxvuR
gI+Qpba+LwnSBf0YsfZZ5SJSAJ51KVYvNPh160cQmZU7V/dbW6I7VxZHIbTL4/TW6L+AJGBfA/8u
F0UulfVZ7KDTJgMKU70Ed06joXZ+UIyalrCnEz7g4dSGsDPD7Pjc8eaNSyZcxbTO47qa8UMWPXL3
UY9KbY4Y/CiODgDdBZljJZEAMk3ZtBb8dEpseT46jn3ruIhm++ZK2CyPkRbatabZWwmWgmYKhfnc
bzqw+p8jmfRF0vZY6+8KUqmR4bY3EbYmj7qUmjoAxtpiSE6DoJLIrpUa8ATy6oCtbUpVMaLiEwUB
DaplSROk32xJYYzMTFDZv66mvsCaYQrww/mK3+le1xyG3eu2Xhd8mXWuSEkJTHgBWjkMYyU9KT9m
7OXSoVearVh+Cu4H1FStWItNQQUzH+zxsH7z+QJpNuw2KTW7IY/m+usP3j8S3VCZ3/ws8GQra9Rm
se/7ygENdwoQSUqS8lwDVccYkjm2C3sjqcM2NiWbFj17m/dWgqzgViY7ZEcVP7ziBvS8ZPzwhXv9
MoAo2UnJPmYlG2iFYoGxxDWVDb6R3mbJaY2b8sK7a5O8I7rkVmijzi2XKP717ZLxI64gNi3cMdIC
Iu9oJtaXbBt7ZqYw1vHDQ4spIcP6k/GKRr/bbUCRfG1U7YzWx4cPTxPuo+xj/Z8mBqoHoPZt6+f0
V7AlD/3nGnKAeB5/hdNOuYFjgpQKBZ8AhNtEt0dIKFXjciSkrRZ1+kjCVYbr8GQ6Q0tixu2nAgNG
OOyo6eQDlDJ6B9wOKPhaXaTjFs+tBFEwAZunTSpSx6t5aXp79zCL2o4qe/2mGEPKJhV07WKp1fVl
p4By+6z7/mprQNu+24lOMDE6AfE/XwbLcboGk7KzYeJIAu+UnYXdsnTVhhplNiyFvBmq4sGvI3EM
zGevePja8TSuY1th/KQDL/giaSEpYJ4a5Gkm9SYpVHC9+Qqa7Sy3t15Y1nXZOJHCBOZPVhxcV0Ah
5j8Y/RcRybJN2JpPv7/o2FPeBPg/qDywo7taEspV95rgtJWYBXxD2i5TqwMtIfD1i8wkzQMq1EvQ
AK6TYxNDqjISA29v0xeM1kUW00B0OgRt1akrJzQGPdhqweAlI4hQIiTAvdvPHhsGZnWYeJJ80Ah4
aDR9OzdGz6h2EVPoRdIhKQahlSFJGT0cn1DFW+G2iiOR5m+TwYfYJO9hJ+uruVa00dlWYsq/ZBYm
wGPjjoIetAFuMnhL4f4dlag5Ws0EWwL3G/2riKpRX28cKr+VviO4qghWxf2k5xOtva4AEfq6egW2
V0eain70zA0AF55OOk1sMKl+EfnMrLnGs0cSIrSZ/qvtQ6JPUQlHpEzZmFRkmdi1VQJZc/njsk9b
3q24HP99wP8nIXk4dU5darhF4dv3qseOQlIV6lw9Qf1ZixCx6DZtV1DcXsQBthvIHucurMZYpEGT
lvcred5ZlBnXi/j33m2/CC6FYKcgLHB1LS2WToc43fgunSUk3yWCwkvxlCfUk8sO1P7UAcCAp0Ah
X/XxP5nVolWEIGDZso9ysYLqtsL5/QYtO0KIUxpVhYn4QeK0rgCDwkdUoXKxEo1hgbB7cQ1snYqV
5rLcltXMu8wXwDQD/CQ972k3k23xs5zAvWT5AC/VRFekhX1U5sr5cxx1clLfnYmwYW/4klaBZe5u
AfA7fXsmCFk/dNk+zVJA9k13UpNlgNiurfYXb0RqaN1BiDTB6xgV+qi5BXo0+9sVzh7aZDNngQZf
1LmnsIdkrzQxnfOEUetpYSJG2aerjaKbCj4k6DfJQD8s6ghb4jTvY63X+entIFPMYlQHxuDBH5Pc
7pYxlaQaTUhoMAz8TIfSGX6gJIa7i8ODyJTCqNp6exuL/RpNwA+eHWEHIYNjl7AkfQHXqJFVXvom
BVogQaDv7ai++5XJp7mjnAR+H8gLHWbymvHB+HkvMWi3iOg5RtYudbck/CjX33QOEERQpOcfKSKc
o3Ulqs67qsEXtousQbCddzPWvZvo7RIWme+Yl1hXG32lh3/jRbeJYjuT0jxIkZM5Apza7rAbKURO
Kfw+hQ5FZA56xpJhrbmHZ5fzDtchNTsdGzzxh3avr+SKDM2Dbz+XD0srZszPckmNwG1nTcjPYqEt
Ah1tywFK/Iv8XZ+uEdgZlQKCiPtCYgKCgF0JCoIFVKC8M4juY83v9UrE9Z4b4CAE0BWt/yL3+ttL
0AYLLd2nFSi8E9Twc55FoJAkY4ZwSaAztMt1oXwFEBDggkKWFF+qc2XIxMsYb6b6kGYODoLATw3a
zDKwRdls5Tf18AqBWJnVthl68T2qCmEfe/EdIwdEOzidCo354+yLCcuSVtuorrSWJH9ObC/ydQ7+
UJm2mjseDO8TjPRIUnDOcBiIN5DR3PEij7n5h8CE5SVWPGVZWvzdxM00ko4Hh8ZV0qsF5rAv9Y59
GRf+/7LMIH5eFl4ZWETAvqWwIadmhRI+cMXWJzX/aiGSw6ttyDzRQr+CEETVb4EUVGfvYst1huvz
RTxnRuNqeXngYc6neICdAmjYXWYR9NbP6zTU6d4Fhn0emipGAddeukj/tgRTGuNKNCO2ruJaXLzJ
Avc8gBuSApCOpPcrX/hVhEuUuyIpilqDpKdr6rSjS22M0+l+46p2XZQzkJXJFRoScsLlE1x/sV6M
krFwrRDCtKTRK4Dg/vA8giiLuDpIKbCu9vwanqq8TVTYNATlP2hLLA89vhgIVXq+Nj2oiQEt4kKE
Uo/25XEM8Mcy2rySV+Z68DdW8va2urycc9kpzZ7gHP8FDL/rI9Vsfp9IqP50YUWSdihvioJYipuY
cINRPWleGnGgq3d7VyNLyuHXkC1mBkBsOImTjNn2GIorEZTA8YOItdzVoRsPkHuPeBSUEW5UMb9F
Wcx5csiq1LnRYiMngcIbrL2nKpdjpWocSEhbt46bdfxPMyaqufaxXhFFYQv2YC7mQf1oFqQmKqTx
lUF5Jt9CgtrORqIOT8fegHO/LPOqQpdq/q4QBhrWkMCt4Ot2vbxo6lkAd3zD6x8BKeSc+BOp1NUB
3XsQ3eQJe45y9TgwNmRv+WSQNQROL9Oap9UtxqTBm0YVoaX5+Rh5RqEF+/F7BeJH0TDLOpbrf2jB
yqF9JMMjvt0K/ttvT63sjb9wtu4D6XqC7iU6ZhXOYkfLEuZFjJa1/m1CgwBR48FhB6YmBp340DuN
48b+eqAvRvGsaVV5PRjp+oEh77fIHk8KAQ6nORsJeYhDpanIPwg+i/NwpEWNUnwCPGKhiJnVbsUM
0Zz+BWBX0sWdO1q9d+i+AlbEHy1BTnM86mNG/fdbqF6kIICA5Ld8iJLT6uubD9O02f4xreoZLDV2
mdNa2Kv5mo8UQYfsXZ7wqooPUZWGVJWDaJFuQRMf+ACiGWvXGvVgJisMiV42MRWiVF23uvqFeYP2
rdz3Fi6eIWBhMEvp+mf9Psh6kNnGAvtEnZ9yUYH/bOvar9SeS7YPFPuKvlTFpa8jPKHEKhel4ZrW
BuXNgiRdTODYpF/4waCg2NceQZ78Nhz/hXKNMudy7etYT5YFyWNJjldLMOlwbl2YXnl7378HnU+z
7ezuvjvXUEPYDbRWoFzAM9TlvScLNzEE0gNztc+hFpJdOdNxwPM/ifuBxfYqadsiwU/B/sgotTL9
3wOdsBsG72CRDx9b7xnOCPpPENfNsB0NdvBoWRkdty87tYK3yYj9wA+u/a8IQIB7NviAKWpwZTcN
IPHI5J4urnnUhcmYkMPziAYnQ/qzLOapFVU2Wxe2lb8/C7PLeY+3Mpo1fv2NhU9lywOh9yL9FzhZ
xt9Ck2oiac13ID3fyIlhkh6GG9FfAI83C6OT11m3RFxSJ7fNU4jquFQ6FCvpUpkHFJTr7Jq6EUPA
ILPI3FCHUkzqO3ZQCnBdLNsZUTV5WEzsMOKgYOWZboToOu6R/pZb3h9N5F/rBujK2lLx3CUi1jwW
Gmnt7VoagbPsf/xkktM+Sofard5EYXCgu3GMGdd0mSqZv7ZEfYIDU29dgr7sV4zlL3lZoIYSxLRo
zdPuXfuzYiXuzodtc+HKaUwM0QV36hpfMZzuvxaR2TbYljGr1qNQuEq2vRdfaWLJXNhpNFCcpcWn
yKMBMY2M8B8r3L+DxfYYzMFLF65DfeTEEvaQXenhHJ+k5ivqBWA4nBkOFAow655flU0jKPePVfzC
emWeJSWBe4gol8OnATAdcAOSIh6TtgaHYRDCga3RlZmzHcisuqd6JbBkPVql+o5jzFtnMG6YK8rU
dvL2sQKnuWoA4qOI5tsFNwslKHCeRvQ1/M2u8RDII7zRK6JJW8V8f8TUuzhx/pv9J1xLPsQXyOnR
KRn7Q+QG34+dH+gdA5LnvGh1YfyZk6hxd6iVuM56vt5WNUcq18xZcNU9dY5bCJtIpTpPKVDCARYR
HKUkBLI8udgc0NuzMJwO1v0AZhY1liI3uyJ7U9QSJRamGTKrWBcoMywO7RmpibbnL+wd3La4c+4l
+bh+YplcTfrVW6tDPELK2c2IZ/5ZwgMzheDwmXeamtKLUl5C4KEYfKmFMG8Z+lodEVHcxPTjwMTP
/C1qZGSE6+kwMrtWmDEnyHbTjQJ3ZP1BcDayun/KBzswdf9fZl0pIH8IniIGQTTXOqIDO/dTG0kr
PwxLg0zR8p3KeDY3Kjf8KGIjJVUCH8zKPu7ORfSoj0J3Rv+wE8/+AoL87OWIkLaFMRV3IO3aaQEG
Jq+CLngu0WB8sr7cU8uauZDxGHER569eeEx/z8q8Z1O14/NB3G8yLETIFJu5tyDYzVypoJnHJEYP
y0CLm7y56AV+qR6rKhZwfEAv8XfaEzTA3xEvFSIGPYL7rZBhd10Nbtzj7mrCCyRDGo34vJP6Omhz
p8thfVCEgoVvLAr2ndYDPRhKxmqQ4L1GYxFz6925+au4L3IfXRVs5I/ZO4HMDViXVVQDHp1Jc1XJ
bHJHrmXunk1lovajbDTN5F+BijNS+Xsys5TYZAAFlszpr5O3hj9JdWttb/gVaavn0cNrw/GVvV8h
q2Tj6Lt8S6I2mWtNIc+jRoO1xTc2QufxPAFqFCtQ0aYOy0i6uRVBfkeb3wJRg08ub1sSdkuyt2dn
QiAOn6sB50wbFn1Nt97+eUhMIBzvOtpM9136ovjROrDalq7fZkrrnxP3DhN3v2+IoZElPXXD2ezZ
NcdTQQKR7MyM01lHK9PaSmSmvDRwvNtJdVtyyTyu5nrb6tKEbkNC97h51NDLAR5VBYVcyZ9Xc3gL
xfwD2z/9F3pYAeuCg6UP1I6fXG+qUqC8tCdJLcRUw1NTApw7iZDbilZpBvfVYpVPAyqGakkeUYem
aOBmTv40oltPTZMfElhoqwl3wP1AxUXyqnRXjEyeFIFUPSdEoZBm3DXc+hd/nnbl5jIejWUyJ2yk
lWZRglyIiHTTCuDiI4cS/WgwQQVXhoSZTeSt241cc97QbY99HOMQawCCk42wK6uT2stq6IBw4rdj
6HKROql4LjFv/Wx5qIv8Vo5+BGL6wY/+RyHa40ASCLetP1xwOX0sLkDOw+uClC9hLtSpjMk5B9vh
YdYbRhy14OmJwuCp38Wg+3ebzPSdn3tx8cnW1sMCX3CL7L8p5nREUvmAg63rM7cJ5sb/PszyukD9
NMZzFmXCX/PXXpdzPAC11C1wK4l4iu3XW/cEqs2PFgvg1ZqQUY9f5zq4yX3tPDdPoNhVZAHl/hqb
aCXH/lDapD6WJBx84Kqr979Vs3IMh2ZGJfQIoKrLdRH2AiKsk+bNgxlNLxcmY2ZRJ6XoMGHXvk6W
Q/xcWg7cj1usUpu8B2EtupC5qijXuvzQsSJeP7DroG4RFUB6Pha/37M4q4O25aSVtbdfVRPuNkMJ
PC3WOCH7iWtv5xgO5ymXL1w4Lcb/2IpCldguMURsBD+dsMjnUwM/6pYsH57jjsehDT+u5t0PWhZY
3h+AN4GjW+z0qyZXOmyM6zmORb5y038Ow+f3+EyZTUELAl1ISsnsgMJMdvw0DNAHwoMX2OievIQU
GZUPPOlrRfJtVdIcB05YG/o7heaV74Vtw+/P+OYA7889ThmyDpsCmsSIfYXnVxqGifA2rhb3hHEL
HlK8291RThbRRbjCugw95z904Od+CNydM53muawI2KSGDy8pW4cEv6cU9c+OgFS17DhzvcZr3S10
W88F3uxsYgCNlNl5b5xldeLlZlHSq0uflLsgKb0KOCUn4fZKcaImzNlTtrvex3KCf6p3aMgU4NpI
XRxJFswcrlPQfLSc+JjcbB1GabaTsxHSmz35WhsAaIOTV6x5v3W9qQ9CTyik7307x0UQuh0mrGRm
9zWZ28Req7moN91lUp/89CqwFMztCOnJn3w0qIrH/fxkt7xmDspKY1zQZdRohKUAaoVbDKr0DB50
i6oTHg8RiepRkuW/Auf61v1k2kl0JzCmKE9Ypzfop81EV4utfC82Ui/7Mo2K2/dh+EqMgd6/J0nf
gS+fzYEygL8lueAGxdywKwPB2RuuS220tH70+CISXHmCB+W56vNOTchAVwhRGimgQANS8RZlk5NA
SuZ4BTfwHmpdeo9XT2FCwjQMkybBLhRYG0X7q4/KIhZAXfqzl0gJbi5cfYCzAYyWsdkb9mhAANPA
Mjtdlzqf8Chtp8y/aHqgWQ3g19IH3NCm2omAXRFl2nJ79Z0RSRY2H9IspDx9O1mw9LECPDUkF5A1
u4xBrMxNtqXPy4lHZnoRK/osjyjcnqglZaMyzOdkis3RY7DCL7O6jtzOf6HsHQpVblvjLesvxiUV
ToNwQhbOtd512jZHN068nM/jMsMss4isdlEt3fLO/ZV4x/AG7aETBMPLw0ccvHsx6xmgfM9vZfJH
CGvT2v6fZslpSdlHhDLLcpGCewjOXqDrbJs8fxM0vbwtWkp7DWntAPCvKVMve+XM0eFYyde+cYBJ
WpVyCF8whs2zurhmXQD4Ser4JMTZH01CAsaEre4XM7Ah9ag52RHHHhlnwgo2Z4y+f4zBvYSVig8m
gG9KnD8wM7zQ0ZFhh5HKcxbbadNCRKUC+cpK3U7dSx1bgvDVrfU3WPTeK4Lyz4c4dHPS6EnA3UdN
TV3XHQgxD+LOfV7UKDvtAh9L2DPlxSn5hP+fw9WRb0LDe8dZXio33EYi86aNHVJ58sxG8d6skItQ
jNfybtfT80aBfUPBpZL7qBqdGHYSsCvE0zO7dC5W8r9s1KbqN6WHmRQa30a2ub5kCQx0yOBEqMZY
+fyfJ3ZOdnTqdJeImTyPYXx00xR31Fr7yjDhrqyzxqIKz/RCNhvhLb9w1J1TQWqL1xsgHyg40Yu7
qnBHGtaISK/KO+4B+3c7zy2wmd++klz7yGN65nV52aljB5jt3s91XAxZTrOGxmYOp/7lNIz+9B+s
8bQNbvhF4ztJ/OhJCm22EIWUcgfvnt8VkuSVmpKPiGSjP+CbF0sYGNwvRooHlgRZgWbp2LsV6CV4
T3MzV4HIGkgsM473DaLDtSHiGFZSEQLbmaIwNQt/bA0Hm19XjYvgeVsGXdJXd8BoB1+7O8Km0vEs
QPSX08SZvu8gxLV+cKVRq0seZpYswCwPvONXsC2CG0A0QK9evOf5xzU6c7Dfqi1Z+nQyb9VdXuPb
dq+tUB2Z6JPkPZG2T4H7Bgccl3t4g9Ppp2h8iYahN7P2rtpU/fPSVeVOTtU2NKe4rrydG/rhpwuu
B38hogO6lB2mVwhTsUslVfnL3ulZIM7GknTefPo79UiOTihPqXe6K+kCu1D98I212Jhd4llCpVcL
Y8OBdcOobieVyTixskE0GN4y+MI5NIajxZt3dOi1pdFhWnVUSHCwKE7ReHIL4mCoX6eqQ8T0PT9Y
91eeXeL+bN46+b6cwG1K4PURcMLeaY7cxSP0nNlXvyeZrb9fRzfTH5MErnx1wNiBPg6SgW+dMr2m
DGC+ZKxJFVrXxhXd+g0YHzCgscyK1Zck8b/LALDd2lB7M7lh1zz6sKxWXg+xtYElRMY4adFpnXiZ
ttX20tKV1gpBob/FLhdVZUnvs7YrXZIY196lQI56SeA+Rs75J2/M/hzSnrRz1+YHfJe/9V5dLqGs
n/M6LH7J/dzAJYUioJd6+6rD0KJXA4Pc76ilkumVgav1HUP04aTu5qlAMqDrCUgnKYstwm7Msiik
c24IjR0lgtBXcG4JDxOJxmdvHs5BXDZcujh0P0PMFM/XDxPnpZKddnRQuiqYAUyEpTzUp4202YWk
KxmJjL2n2RHPb3FwwNkrm7L3x7TeeVFmSn+zrXDrrEDMZCF7GYG3G7AF3YhPaAThIGmywdvmuq6j
bZ533cWZucIJypgivcpP5WaY2F4lbLw12v1w5WCkgiNP3octmk4O9g9FJS558Mio8GIHkprrVzcb
aXMC1pFWZwn9gLoMq+6zqNiQ0t+3Gj2FhiY4BYrZqEbhWzY/VVRZYmnOtaQaeTFxU1XHBGRx46cB
t9yOru1KFYKdvsqHCy92MdrbmIEOFgO2RsERKSenwbd9irt8Uc2ASAd+Q0eGeP+tvVI8ZOY5yIAp
mhgyMIc5suOs7j0iLdGaOA8cJu7jyAfTsp6MZgpq8WSTHtNm6CJGnesXBenYVmynVFycYLfvD5o8
bImgI01F3EStl3gBbfDnADzvz99/oDMQG8gJUiSwPFEjCyR/+ZWY9IIdICG3u4idGaxVILz+BTNk
0cDMUu1YffUWXjz9LO4ZVfQI2mbhnekK8K7UWqxosz5QsqDlQmIP4HqI/kYsdS6YXVOgaKO4wv2V
ALfkV1bLW4MZRAlEOf+oE7dDMxFbGTUPeBX4i6BnzsugJuE6UA18MpMu9xCcICkul5i5hfE8NSe3
ihrm+0YznVJr+MqpfsCNuaa6u8Tf0WSa5Ug7eD21BowvzL6a3BJWduijNN0wOZcQHznkgoNhfTgx
zsC9lTHCMmtmXkPt7vzv0SATBKKbZYyWUE5RH2YFJRygZqmmQ6f2zpR/31uM6VsWW3ehIMi6j2DU
o9vEd294s6qFk3tRXaW1VZKbB5d3zSTK0EwTOwcyqRfP+lfW5dagVTFIeUr65GjO/X46gF2GZ+VX
5szLUKJ8JEZdiLL8L6paJwYV9umluk/zZmUzSgBcE8bXOJo9lACWbyb3WQ3hOWwl62C8S7c1cKj/
bqLWYYD2ABPze04BzTZM5ry4ZWVDJq0oPvz4f1CSDme+qdGxFrCpr6abOjYmGYI89w97EJAESX00
Qit1DN9/fwTuCSsNTP4IBAi4qS9aSws3jLdonDYOC9//NFAiKp5uvMzxq4jOldeqc/kaUItUkuPH
Y9qIMfJ8i5Ucn/pA95/rTJkpR+MhWzJfUNp7fGNhqCshFzKMFL3fx4B/jRsmYp7JRcSQQEw+06zm
n4M3lixvt/aDzUHE7nYMpXRnVDxURz8Y4ealoO7I+hsUgD/8/w5cO7IamVRWgAWq2IFHF+acjrWQ
tOdy1tapLiam2C97S5xAVVpVQCR5uaXN55vNzyATGgFvht3ID7qmTkEd2zLvJIv/Qf/M3xDTJnLL
Vuv+LDabZvHQy3GzWxAjwFsWED96ErGn4sMMzXVbM/uQRPFQt/qKZGi7Cd6k+XlZCzq/iE/KU1eU
i9SIlL93rdljQfXNWpGsSZgwYaajGWxhYVgW5syn0pRtJed1gbJV3TlJtsWtHZgtvNDAk+JloJS8
entlvrBw5GX5rW1dnWVCLWOKbzPykCZc5Arcuohtx8dm0/Vqbt6aycesdrWGn2Zgw55qUYOkyFFn
DfwqrcfQJN9miRgLp0wRUp9bM0VWR/DSJdrEX4sSRc/tRxSzZ/oQUeKaWchZNXMPwMK90FJggQyV
aN2yG2InTgJU8QPJ864dv/DXdvIE7T/uLLumhAeWOIHKQ2r24HtoqtS/2n1Kpi8s78QhbLsn2hCl
Vy3bemYPrM3Fw8RwkWnZOw0p3/e3bWjo81bUNcMEa/UvlbjSIiwbAh8g9gxHj6Fxk0RnuRTcN1Dw
4uVEHlwoddjh83nRXeVZetXz95mDUtwGuwyj9/3QtbSJg2LofXrKLUYGYki3vy2z0eqUup8mHWF0
f13AyACuJekpDDwuXqmtjXXwKb3rUTeW07gH3YpSVWYVf8OBWZPROPkTbgKp9LZyVme1lV/f70dJ
JuDF2kBNCnW7ExjOd1/rnzofpXBAnvHxSLtyurOJW0Em6brmmfLvd8eRRKkZSPjXFqkZG4U4Xllm
XiUJFnQBH/CN5ovsjvcVFodaNM7GH5lVPaf3edHVr9DRSFAAa1IZSS2N++IhXbLPVN7sqZVE4WQ9
CATA3M8omjPC2GItRyGixw41Ce8+Q85MMh18uVRnP11L12xoeppeOieXo6ge/jrNupZA2zsjsFre
PajKDnL/A6qLQ3VrA7R5FIpZiKuc17f2QW2r0d+cNNAEO61kSfMCHnzWY/1gJkE0fenOdwAFqncO
RtS43dir3RGR0CDCbS0F5Q5ZkKYmPICW0Z/NjrkONN/P0fymj5Slp8qbUMUW0mT0i7LB2NlnxwfY
iD9BIoZ78oUc8JvPiZFJq+gJ6nvSgxMeZVlk/EodsEOAP2Jm2c1v9zP+HszhzzoEMhcP7tWnFl74
OOln3LeHZmL74S48yPuGIm4DqcRmeZvtSlL46PcEjDTOK2bf0OWFxyOypDYa/H+gZvq71HSgxcnH
+sWewpWou1hBFTF8hnwpr4RWYOoRVYiO5Gc1aENJxudmoQV4phLqJgSma9akaF28nR5gNHeBxq5B
jLRSWVgcf73XmKNKuibdYov2C2osgiEa0Xwd+WxZiswAZYfDqH7aZRBnS0B6t3prNPKcLKhQej2n
b+coWHGmnkWdxw8WacblKX6GnKoJBpAsUYs+2Vkn8CctrAyV10alM8VYYcY3LDCJEIOva6i1qitU
A7Zji+jUHmH2kaJOYIhy6nvOc/kbIREbsc8OA3D4vT/LWN2xdrm9NOyt6R3OHJKRv0Q4kRlr1MmO
UrStWzFJ9EBCZ1eK0ezC13TrPHHRKgsRFSmolgKzvyec8OE20AepomdZHF3AY2FGpO6Q/6qGkDr6
0ppE/GO2murfCk267yv1de3ECsrTRDDfQOfvvUOcRdkj9LCpQvq+GSicm+1nagzVkLPOJhIIrBwi
xNs7bLekzFHRmCYm4ErOfBNL1aflkeOzxdARoM31RdIDJ/v4iFMQlc6NHQyL7pXzRu9WayyWtnu+
LSgTS5VO8vMVtPIDSSv7pSIy8CjfVsSDKa1LIMvUUebmAvjQR2i5UOLy/xNTmPBCB8NGejhZD5tz
YXJIW4OUBM/Wx4hv7bVhazueONmTCgmshpkBsehzvK7dLI8nPfjn3hjT29wyuSS309RrDr7dOKO2
Q/EBb4zctABgYREqqtAPqFZ3Nw5N6ww6eca2Ad8yKVALBfPDknn+GwtwUoKimemsAFun6cJzw79A
Te4WiEx5wz8HgxpAO0k2mIIxB3Biwwmf7c3JIDpVkgnT/IcWH8XgjA+2YchQb+z4WD7zDJekhpXR
xTNfvnS503oDr3XyCeaITF+MfSd0i6XFxl4XdRMkJekxOVAtW6fmDRPUsqMVTVskIh89umk4/mb4
niYnLwOwVu1tlguNzDxVl2jIj9RwtPCUPNz8T6atokHrGwwdHCAMIH8v4sa8eU/AM1aKXl9TvO9r
HzfMgo9nEdEcB+S/Iikkg84GM+MjdrpU/a47hTCGoExAXWmOtj2PQLOcN06kYvnMQu4+nrn3L+yX
2J1tfHctVE4HId2ta2X7CZJ6Obrm7gdz+n4bNwz7eIFX02Bti/x6bZb4BV/Eo0LgZe8gzN9ncdiy
PwBufedcvJw3cQOEivwhOpEgIFTYzveBM4VqYpkOxWOdB7P50bBz/cuHrn7QaJe7+JObLRjceyXO
X54Nn2Ccf+RvLBGwWKxovRyXAhLFtaiy5p0Iyc9GtY0ZuV383Gi44f0uvacS6YQ0kL0lkCQ/5S+7
fRxaTlNMst4G1egx2fWtK1rsMLiOPl7HpoYDsHlC2bi3f0ZsVz0EMp/EjO2A7hcu0ECWUE49DtZE
eV3SDFqLAh+eo0YEDQojzfL6rlNM+4rS9mUxfl6avU6fdpahA4Pjrf1/4fEmvR6xRXwoy0FEiUne
YltdAijIJENCRlK6US3vOCz974pymDih1zKMPkhnHdWhQFr6Azyt8BrRNwBqvZSVOQeLmNxBJzkO
UfEceoOOOJOAh8EIjSmKzxEX9oAa/d8PpUSf3SE4tZwOb70pKUjZUWxxIeYkxguU4wwFwuuUrK0/
6cLR8c2gfDQx86d7vFdkh848Kvx+SeOiwWGOB5zasGDTV3Hs7D48a4oHBx5q/l+4/yH/YgApbg1w
3X7q2BXspLbEFTeDlsiUBOtMqbp9pp4NWkLAh9zlbSFGgaL1HnBErrC1kZi+mH62MEt6DKOZROLC
P8b7tRTejiUzUFJ3xMOYBvHn/gGha7vkdX7eDvZaLgN2ko6gP08IUqUeN2Oox6VHhpNN4anJApF2
Z262F+RGmPGp5aASmKEd2iAKw8KiyJwXas6r5Qq0BjRCbDeOzkRhMy3LLjOOj0sLHk9s7RUlnjSr
iyWOyFrzL852jQni6uWPLwPSW0kMd/mf+8hhgp6NYIhjzBqyFSTvDx1HsGgMHPYSdsJQa/tZ7DVT
m/fVMHLBP0GONi+SDy4JeYAd5/Fpuu/l0zM1Nt470aPgamGjA8d7VatXxgFpghy4eUAce3Gy5pzo
BA/ji6CqU3caFzRbXuBilql7bqX+EOMZyNU9hiA/tKyRgh+cnUqggWYL2p0TQIcFLrGqFDquy8tt
SIiZuw5CEvLpPwwyXpGS8HRq1Xhl1PNHdkQkbI1y4p9ARy+RQrpYA9pU/LB8ipytdhYTHyDM+stx
SJoTFB4fkn8Z/1qQtgDz514LybwOH6qjPwr2kTjmZXD+GEOEX0yspDOzK/xV/FWtd7TDi2GJmmF3
gse6wLYw9Jba9tSRbBGJhSuxUXGio7lPOtkcs6n08ZRe2itxfMZVYf4Rp6yekTpNiUe3kS5tTlEF
wjQ2iItr82uZI7xE3EPx18K/Oz73s5D7Kzqkaqx5nRZS8OB3K8Xg16xaVc18EZc9ys9g2HEVu14B
g6gZLeSvfdUWJ2cVQImOg6KLtS1hbVy3QeY9tu7+V/Txg7VqPVIC1cHIPPMuRmclMH1hH0gY3kzA
jux2r/OsvSbxDK4gieYZhfQo1bDEze0Wxy3pjE+OhTgrD89zWv1fd0YpxCtXpUsQvm8UP2jy2s5/
9aMH2yLGcTiVxlihgZE196lbExU8xABBI2ttYQIUlPQ+yMHaK+q/T3UW1vHq0MvPN5+QXy2GJTOy
hatL5AT4RstUPDPbKidiKlByzCMZbTk8ydHi8qEiHGZR2GZueuhNgLxZgJrx5WIStojye6x6yDL8
65RTqtux269N7JRPVRmuqBmTUpA7V5/SrdzCPsq1z1BVxlYJRXeoiq8AmD6mGhCsqLAcaKeK48d/
iUnIvSbSf5xlJS2Y9KbucBnkIDhEs7EeK+UKYzj8s4n5lvjCwNRUyRKDForO2oHtHnT4/qknvY5b
r2R7Ak6P49mjsu723f89Q7iyxqGYoUSnYfuzi4xiE+BHq3i9/BaX8mWChe3OkLogDvInmOoiDbFB
Hixm/aR91NTTyj1tVYha6ri4Vl6EVeCCIYll1PwkP4kn3cCF4FsrIIh/WUxGMaS7eCok78bpFIhg
gktuOoVctTc9PjG8wOr8maFEAvQiCaJa7HqBrJiyj4fUoD7ve/thoJzXpNImytaL+txIrZ/2eoyP
469GSuN9MhR9Me7NiB39yTT0sY4ewHHwQyApUfJbvTjecYg5uMEi7TqB+QOzzK0DRGW3v3UQ75Nb
xf2UX+qzmJYaeZOFxdCcwoBKlE9NUCNFY/sclVlzDb3n45HFFeTSl9aD8KsXIxhznXpKuLoUUnUL
4raD4iWRc7nf8nKpaVQWsF+jPPM2xb9zGY44fW6dbsSjIFWwwzenSpAA9WiUt+hY4eGjmW9WPUEW
3npf/acrRj6EKhK9pCLVKgH0wrNjV8fnXbXg7JVHyTSj9uK5DHBxAnKfXwLkSD0Nc0AWC7L0uO/9
F/uuk/fxIj2ZEBa4py8tHGZkwt9yWut5+/kJ+hqQV8Poic8ABREuGdhY66HnvPm+vSCGFVggt1Qz
oTvru2iZ48waqdoZtSlMvaeDjDmKTPMLH7UyDWKEFvXKBixmASVmSoQpVqedglE5EZ9q5GeloXCx
qUwLn/kaMzIQ+ZC62D14MQqIsJJAM0pfzrFg2oZDA8BaCpQjp5W0TgJWqaOB7r0NUvIzuhHbBmQH
8ziQzYSaY+imrQ8iEzv5VsFRCFGuN0f4809cvz0UxEfhDFIC5SAjeAmWrDSh2IVHSj83wqfWgIzr
8rCKQK9ieNREbbpsE6HbaA3cdq+U/VY58wQGrIvBE8YdygnptFvnwq2meFiim+yTTSRU+lA88KjX
+ZMGZfyXgHJcjYXXX5waSdKjpq6uOgxCcpNgbL6+LISt76bOI2PI7PeNm6dkQ9VWXInWP7uBF8qx
T5aZydbzjCM3Oiu0g0V1FEFvPRfgkj/QE6+K5AYtZz+MqSvQ8DC1jSeHv1HiO5/VyTqIucw3pqCH
RIGh9iTl2USDW0Nm8adwBbe1YR6ak0VHttkZJEJLSjooX2SZOneLDTypVH67R3NrOBedM0W3SwSN
FTTLl/llKTdOVfNdT2geR/ykQyu2gHIKIV5WKAJbJdbkZIJohNlUSfbfo7t+US1ZQp0kBR9mObes
DhaN1XinOS9vU/dWIe03zUunvKx2RGy4pqyVn8xhlxYR86UbT2XwAIjv/nfLnBrVo0HT5e9Z9Cuw
eewlgLFd4mkqV0d7XGdioTn5R3ECHAhJ2yFodQq08PZ0zBUoggYC8w6V4U4KLxmPiNydcdfbc455
AZzrNdwtv9AjLH6XWSX10JSgJ96BZAWeSxZQ/bYjblUhgt/SQ1wvyRdHoLu9GXfli2hryjGE/ycD
iK55zIXYWRLMAoi5JnFTdwYYPdDcerj+fXOhVvzeCz2tcJ6bBlDHmGt3llDEpW8yAl3OLJsWRyfj
aWpd1wafmlMBo9E/FVbcl+PCAonAoDUDPjs8rj+Nm1RrsPs91vGOqLiFO6dOqMMMt1N6WJElLuMr
GWjghnJVTQODd+m9dh/zeVjHKlxnEmm6POR5S8t3sM+7W0rFWqOwnNFFqkDl7Z1H+eOlH6/yQ37T
8lPh/jVUUqB88b+JUVArTugBSoJOOq1YL1VaXaj7y2OrO3zLIPrQYEmG+bWoaysGOMTlo+JQ5dlV
rwXtIXNBYaO1MbPIx1sS3KOvNGcn8ipO2p3nBPa7AJ03UmOia/FJPbxaIQL6WDpe8I5h9550nTrp
Xdb80xsssfQrkdZUh7hrIR3Or91oKAwo9U6qbbpjVHo3sz0res82ANEBgPBYf/qfMICbFbH5UQLj
rBUuPpgeA9SQdhSG9ZgF8S51/zsXGVDnMBuiet4FPZPx6Lu5qI4rJiNTKhqsgTMuOxRmvDmA4c5e
eu1WxuJTB/N2ZioUutroZPl4cwVjIBJYwJUGzXytGE9jGwiICouuyqLJxOdwJpQ61ATAnjIJC9dX
GBjISF66GidGw5p0w33fqgICMN4hFmX/fQM/11gP6LT/nIx/Xr6R+EtHAP90im9dhEs9DBIc4PbG
4SNQ5uzXix9lVojiHFfi1a/rmW3CEuYvBoQZf0upDUDPM7h1/2J9IAQyUX85wJvt8T3H6gLvM2kc
qTx8NxCRvo10e0LMfHfin8s2xcUtSUAL1I8flcf1IBQzd39Ra9vJG9W26KJcPvQF0q6TewQRj8V5
bMt2D4WXTsgx3MIp9TGoYcKG+LXEy8fpgM8vyhfoXHq5yPtvoItOkaP2CS3tHf/E7/WLjHFQMolY
Yw==
`pragma protect end_protected
