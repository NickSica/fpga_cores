`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1584)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5HeicKNw6vVu0avX3B/XrF1BeqBJt9ZeDgW5CDxoyofZURzRzprtod2+
c6hsydZ665B3vQsmD0m+fIOuN1WawwjUzkvozH7JrwIp43DvJIAeTrk4M9SZBHAprWHhPX9nMCw8
gIA2ticIyNoZ3WkA9RTQzFO8UqvyTfnemB/7dQQYRr7r6xKoIFzVXmVfn5QqnZfXoG7S9zs/lWHq
6TISzKeeJHuKF0v/PooVp73td2EUjOuBn58uzeRwWNkdFBW65gTuqVkqi+ffuj6nE/B6W2W7KMuS
GxmX/5uWaqhiTGGdNGDkpRSt4MdXcOIkGvxAiKQDboPa/PFKqcQhqQUcGU/YCfF7OplE/NBN1i9C
Uw4m5Y/6gzEVmdMAG6bUxRKHRd/mXYfeZMsTwgyrztyzDlGiiMk8K4MqmjRf+3ktYuETr6XEYun3
mLZvOqVug4x0kcTWqYK5/00or6hwyG1NETWSdyXOS1+ZczQPmX9SwXB84/lcR41Els7jgd89gJnI
0ZeL23l3Frd5uoQjslM98X/mLTBLRAJ6ZMuSJG4iUVh7jkzHrD/0Ah9KqWSzbrFxYEIBNZpZUTaV
Y6DD5Kxkc+WWPleOYwkqbYFBzrEFtRfsjbgtbobCzzfEyZT8P2piglbwKfHyONH0Pt4qfJrOYSsc
3MLNZ7EldS63EXv0doUXQzU/tHNCmcqEGx6y0jdOxqaXAN86DlP7/CTgdZKNPbIT5rYSJh5Tv0Ts
TvMHAoahAAC1TzfW2zfICbfv8mZ47NoatiUqo9FMABWhvpt/EW3fEGHsbJ5EzIvQ+H5tTmX1154D
kUlDZd/jmM40g5glPjU5MOrCmdcYvE5GeQwMZ1Dv2O7XyX7HvhIYQ4vqJkA7TbywgH3unW5/hieW
znCAihXZX3yLj+QCtUFWP8t+8F3yhN4OYXfLTyeChjVT5fPE3GTrnGwhHRv20QIGRzCWvTrOTxUb
gBD+uxQeThY+GOAZ5ldeTdf9oI3ksoGb/nbzMLWEVrQcg5URMw2pDrvCK6TOAZvbskPWyNeHVPlx
3hmSkTT+BFHyGu2aW5lIXYno/IXC8LPd9QIGOgnxMG+fAoSYou0p1ls9Qe59nijvJEaPl8L2T8cO
BTPj0jADG/UOrUFc7uoTqlwAOBiA427rr2yI4BsbwiuRa0JGDmf6juHJZ7NBuv/XFTiYU5YkBjwH
4Amvb6/wwwPIcN3I5s3wbDskxT80mHSryl/FgTGXGp+JXbvIG9QcPf3u7hP+SaPzhvMJZRidxFjo
qTiWD9G4r2z/QHQ6bQWld3l/bg5xekih3IR5ppqf6jcGz/tfkKMfI3a/5OXMIuz3ec7PvRKp7qXt
0YMO1C6PSgjxItD75NqmiCdOH11dKl+FqA4C75YoV18HvlxjuehqM8yFRfNvDbs+SOt1l1TSY7GU
vosZTNlMx81FukV9ndCIRcz+a417MicOwa+VedYrWfkzH0u+zETujZoohEKAWwukArIIdC+zl74A
ctTCrEIf04X6m6lVcRPSjpxsdI0wGEDMa92etTX9dkU9vpSRoRPGo1EqcFcEOeJHM5w7McmijAhz
iRut2BMOvo07Agx90UyL9zBk4YjbJexVOC8Z1l06NvlELEYcEFB+yJe1RLQC6YMSnv1uqWNOapeD
QB3o685duE320av9pgl1RPLt9njgAujCiEZQiOimkhj+ThYLJIYtqqbufKreMR3hpsCwBvmMwLGv
RSW9AtSD4/TTJYo56UHETrq2nLlKFKzjAnSaJYWXxboW0EEujTn4G5+Rydxj8tTumZA5+N+rfwY8
oQ9DaYBxLghkFv2K28DCsiocAJ9O/Ruf4y21pRhACHP6x7HjLkXSRg3EVP4zY3lSrParKAE57zPG
8eL2AL8zGVFdj+x0GsnDcJQvERN8oinkIGIA4cGJVCmrc92WBQ4+FIpgiZEhg3bukghVaEdC/CyK
ULZNXx28cecsVbVA5S1+RIb3t0G3xw+ihFbZ/7//EUW55dLAxT6rJxUELSxI8pqqeqSY3jfMHZdq
osvJngOWXTBMisqwrJpCl6nvJlTLenr7j8NW6M2KGfB6NMX6zweONzXVVCDV
`pragma protect end_protected
