`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
R1WqgqFekyFBf+R1EmSjRCQxUuOx6MT9aQyodTNNebOe0CK13nDxh2Wir1luIC2E+1RiIa720P7G
30ynEHVRjA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KNMY+1Jln0fE2Hw6EJV59uwRAjQ2BHIWVdMuSpeAltv11pWP/JZCrd4z/uZcVTngSRY8jZzhCZTQ
WJ4MxCfVaXUWBZm7mY0qLw6qcMnyzincQFakqwRdOx84IckfsGjNGJ3OEjUVkf7dW/J0o6KJvGRq
A/P9gVOYmGcnWb2CkLI=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
sL7gG3oizEXkzDHancu7/45cwKfdv4EnXAdeK54QMEX/eoc5P95Q2IxqcI+tnVljSH1drXWj0Eb6
Of0W/iXPKZ8OP77HA72GpMs5rDnQtlgP3rECZlxuTJ9RMJVfJzzO19m/vMWeqMysX1t8PW29rrsf
0Tqwcs84OG2uxBTuyDEWCBSCU7Yk0aBYU4VmF2rkELqh6jo2Q/udlKIUXrwoYSdX0O9uon++5ahv
mjzu8SGK6zkA4uqzG9ghLIe8qBE6KYXQuzvdlMdTVdy8eHbCbzVTNoB6j51Qlq+S5oMMSQvxBaRz
DIAN76FuevwCbX/XKHESsvee5Sen235LJDeW6Q==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NTwqMfOwske0aroynepwGO4Lz00SLylJkTISN8LAcq5uE8ZoeT6aFHS3yIuZsI6EEE3s5mQQ8Cob
RXh00Ler2BvOA4K7lNGJUpMzGqJI7MZao2GijCVpdWL1r0vSvaacAIY9nlusgQmU63NqWs7cQx1t
7NMmVlpgPTHr3KxO5lMNWR2EuXJ0I0zOxQbbrTneEEip68PBGwJFyFdSjQNe3iwSj7O0u1NlI0nF
01F/RGHelGngznubnZikT85LEu94GTbx+WNlMlaxWaxuIaRvhH8UG7MPhsxH6x7sS5ZS9GHBkFDK
gyo/ARDW7a6331M9HUgGOcgw3trs1/Klf0nskg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
F0eZzxJQxbI/Xk9S9oAxZw5Tpi91CrcqL3BrQB2lyqn9Vl25Garq+8JIOwcSUfEju0nEdI9Cvd5l
ooe0NMs4K3iY8tnE+FiNZhFGnmyV5djhXaAeRPiaySzeXAc0nSnoahW36RgdEHyPbHBrMfq1pT3d
S/0aa8cloJNV0EZcGFq/QrhQOhscPpDi8uk4IV75ihx4K3Y6D/SPBsIijokh2lVOyPsWt72NbpFl
R1J6iXczzSEND79HNenePfXgQ1Sr+h8Z2ujGHirxn/++xFCAHxWZmhGcFFwVO7AI15b3pfNiyQF1
2SACCg7/b/5q/JpHGBLoFY5e10UGMoGkaXNq2g==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eShHfvBzKaZ/Wp/QUxGlK7/6Td59dAgzaJsrKOgtjc73r+sFOocLpKUK8YR7XmM0pkfLOBkjrXYq
jGiy10qSwBo8l2eE17VZo8T9nQ0IB2FFGgVl0zNGiZaKSzE4a7K5so8c5gtUyyVlyHWXKqYAj6Ro
NzUEnqMqJPppbTPQbvI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
VtDvfrNdg+YlmytFZV1nO9Ch/hNzGllGY3c+wOLUGxBvYhloxzDDcAB/7/ljwrwghZilvxZm/DJg
2fzdltt6rugwiyCDZPTj9bYqZhAAM0bSdp5YpZP0gTz8EvbCxUo8+Op+ufZee7A2QX4lG973f4tu
FbV42AkOjECD3RCU/zC8zhB5kCMonmYQSEe1sGWBe2+Ga49sur53s1VC1GSUOY3PQLHNqtwSq2Ra
owo+cSlmwu7mHpq7nDvHG8vWLm58VKt4pglBRfC9BYdbhmSQeWT4IcMsVz3wzwUMY4HmFkj+0Htu
JAA3fKLFH4/svF3ilwX+klAmiEhOn+ftw2QOyw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HHgo2A7au8S1PE/PLf9TgssZhqFUk1LyRHoBPoQd7KZOhYH8iTwJV9W8hjvxzC2Na0peqSJ5zF18
7DRfKJ++XfNw8OtnyxfjOhMGRjIzpk9/xlZOxoCpZPFsl6WTW8CoN0RLlh22HuIAeiFQu4jBiY8s
f/eG3F7z8aDUIS222+2y8Lc0ifWDx1YbNoJritsavlDA9L9WOwq+EXi3pvUCyXszhqfkMn1JVCVR
qUhUx37i3M4UJEKXpk5rfAol3dwNa+jlOtqwiBj8/VnhZxY2i53S+bX3OP8N1Zx5wRoa1UkpaXLd
9XQOggc4VKKTgU9CJZPlRk8FrwN41qv2G8xfRQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16736)
`pragma protect data_block
eeCl3Hcc/V4mGRBHBrnlVKP4yhCz5zwFqZyK1LMRDWNokFHL1R0AV+Xt07jE/v4WEVNKL6BkzYsk
yQ/FPwT4uZH0Zk3sdjF1YjE0wvrNTAEPInzcF4TyR/LAJkNOc2jzF5Afl/lbRQgFgaaKnM8GyDQ8
+MmkSOGV+xrNIKx5FPoAuesHkpVtr9O+YHexKjZnFP0N5SsJci6c/e1tghPdvWIrShbe0VgllpiG
UBjsaFjtl02kpxwy5bX1PElcNUyU5GYvGzZb0JncjVDuU01XoOJp1LbV6G4tf7vVsr7DnIRSZUhj
4/1rEpJNt9AVEAO52IYYlNIDCbz0aG9mtAlqL2A+oUBh8ajoqTWAetMHpTUbknAbIb8nt4QdT4Ei
y6PK0mhcIUivnRs8WAVYWMIyUGBgToZvVJLMwrMmGypQvn7TvNOM3BzttfSJb6btIrza6/ZL3fLc
s2cvJbvon1MySM/mNFJoBbFhuLoAEWPmuAnJus/ozYr21/+r8aaUn+KBkkLg8ObhDzlOjZesR2VW
mAaLtUfyaB387XusiLZl2K+w1cGkhUP+Q5ezKdHRCoQL3HD+XTPlJvHwBY7PuPKcFfcbRz2I5Cbd
lJs+vlOpSDoYGO0yAqjE7LwMzlA+Le6N9Jb+Yxk6cJc7VIRKHg7akAtpGL+JkEMHj54lawbPYrIG
12l/FKZb3cwnBHGjlJn/jPf5cBcokQa4vMenbG6JFb09/sw9Pe48lOVgvlQZSCU9jvxLWnYwiFHO
oBl1uN9iOEoyvXckQ0yJHfTfZu5egB1OG0b6Uet+gVRVJGyq7BtWgmnfNmfbnCgS+A4lGgHJyo5h
Vellq8BG61whbdvJ3UEiKFqru/rt/HUYLlDBsJqGjth3VAPqEiUHlX0sus4E+Zcz4z60+CBmxh7r
A5wrfC/SddGftHSDcrCvNOLo5c2D2Eqc/g96BhRJvf6THx5wShZ1u6ugUnQ6IHRqi2F7/n+nHiku
A+VXfGQGMuQb7VbM0agyK//W9BXe71vZTnepbl3wvUh/S0LVDqlbY4exz3SQ56ANycjqNiQ9hplK
ndKLkzpIJOTvB191YrwCzYd+Eg4UXCCzvKr3rNcKnlYiWluMO3SgN2sDzNOXRvxNme9fOFXdGZVl
BhkmIQQfI60u+TKu9xnHBy3b3oetO5SYYGMVHxSSOn2gJ/maLJ/Xr6gNHtS4ee7r2QLMHPaZ0e2j
+cAcEb1sknPMXhR00wcDuRYCz8JvDWvg7u1ljNTSjB20Vmit+m2t/b/K/tgUzzdWvAvPoiK9StIr
w4/Ns+pCFR9iE1OlVNItc44YvHPBe+Ld/u1NjnKfd6dg+aOi2ExZfp2KzZu1VEbrJ77uv3JixeqZ
pPSohrbT6MWzbXPwze1Fq37AnQa9Qf8v5XnxhCyqcNSG3o0tATSQqIrSybG/J/GEkfdDGWma8Ect
68fB3ea8PrKMS3rLE9DXZ9vgDyR92OVwOrl5OXXUdY/s/HIn7nw/exxksdygDmsaI6vW6GKoWng6
bCmR2g3bJf50yFN3lO2E+xeZfSg6ScB57dW4B6RJ0O1LqTmJd2r4EoOB9SlU6fHSTmMC31R1TbMu
PK8GVFsKCvi/tDQQSIprVPPvjcShCvlYUHIyX5fxrGB2a+5V8YmxunaRdOg0LxIDFxSRzV3iJAg2
tPgHTAe6A66tLervjurU2ZOfG27UHdg/ZYoKz97cEXjq6yB0JwtniS38z4n99lOSXKkc6illasdf
i9+zk6OZewZ4sBgQ538VhILy7oSHnvs2AkoMHTxhIc5yg+p1TtV8WFcgSJKyahcZ9AvCJd8/RHah
IEKF9c93dBih48o1X/a4Ymeg1icgKQ8UHMX2pATO8fwOmlBv4OAkhFSlOw5xWt6Na1IXLoXydDh4
NhMDxktHRC98qkhsUOMcUdyZceQkQbpNx+Nhn4qWrPoa1PKJTD4j9HkFreljr828T2Yn8gQGHILy
fqAiS6SpWorDMeL56fX/8kOeNZLwqVBZfb4uj+68i+WGzb3R6JS4WOnjQMogqHGT2DSozUrbJb5n
b9u9rfwkU0inrIUwqymu/muJp8Cu8+0TckpGu+8RKHpMImqsYM6xCinrFOWIqSpJxXW9pLPAjSEp
P5NJG5Utsg2QS6S4eFo6CHm+lTarMOUbBEqGDrIhp1G0O1WHIZvw5xglvU7OWu0arlTkB30QKNzB
MalIydLfCzI2L2eW9SYLuAQ5DUd3aSbc8YmgZnZ/oOiLXyaZxJoZPkDTYNHTeG5cPyMp+VdRMrS7
ce/1peRtU+9uYKBZgyP+QCmteCnQ0fgJutT4O0gpG7uExBZ0g2IFoCr7ZV9tCj2HVtl4fr1Ej9Mf
qi0IN67cqhbkL+CQJg9wVsWPamnlubwMGNqJ6NdGlcPh+Aev5+kKltB92MYfB2KBUEXMHzay1WCF
MZfxDbHj2TTDtGTAkXDcgdzJdWJeTw1pPgtfUEnN40PrIIqrIb54dHTV8nzlWvungME0SREqOqKZ
8pzVHZMH3vtNG1MQ5UKThuukBt5mc87SWJIfBdx/bmyyfgV9rJ/HJx98tcThU3jz2GEH6pfZgE52
irimyYdcnz1rvvpj7HAlJOtjPjDEtTG0etEO9Qn95djgQ1FoamftAzicl+1CWwtQP0mPNsKEY/4h
PGlmuYc3FifUhXhXEv3uWpI+TVDmawylc8F1Kkn6mOnPvHNJI/vpRV0qkmkEIl6TA4JvQtz1oT5F
kS6wsEt1tCUzeXABWjtUiogcYZb5vl5/NLpPkIi3vGGJFEZ+P2oyxaU4XUVzZfW4B9msBytPBEsr
SovaK1wWABUwjO7wHWuGaX3/L+Tx5/mu84ZhzuDhVS0X8by48Zk4i2Y/8F9MGGVVJLkh5uFklzxC
9lsLBqd4pxrnQndp5Rr5bDwY2iqdYZ0F+N7gUgAn0tzuDgRkH7SSxRjqtgkqOvma7pOcV9Hq/A0I
m7idqkQEWVzU8UY61fJz11MRu5D7wsA93r1VODY5z//yRAn+JtAto2deJB5iSjLjUyrnbUiZ7KQP
U60iQgixgu9cnfMK3m+qjwwKucnCKIHu+3lbv1ity2INNAkslccaknhlGiCMUsuFFCauzAbDOQfo
RNYJvIgfnyLwJZpP2bVx8+1pUn+Cf2beZxGJNgiDf3IbQvHtVFYjvr0Hgn4d2Mp8vOPZU9L1gI8s
EFWOI1L0mgaN4MZp2jl8OIJplSFm/YOZHpy/Jx3l2bhh7AHubBKvxXkZLklORJV/Th/xzyV63WcW
w6SQQv3/nXcVgovMTPXrUVxOz6EmamrgJ3+6qjCY1aGPC9t+kSlyOxgbW/j9FagBdwMejvLA+p9P
5ItqAyYymidsY/bqFXhPKw44DRmK5L3OQ3S2GS/ZQLz3KNpiEVgP0tyt0O698xP+wZHIVSMAzyTj
3kDMIybbbs1tt0gpdZTeUDz+cToU5EAn9YIgHA/xwAr0jiX/+zqjehQhG7wGv253/4yAF0j2Z8WJ
nK6KpgLiluF/yiBpoXPk6O3MRRP5t5I4Jrj9fSkEY0foozuFpZxIUbrR3rRsHPFwY9gvGJ6ZBlQJ
YZXi/6qPSbpgTJNjtDsnZ6I//eCymveQyt178/25F+taPJ5zBacZV/1Zrs5Gn1ty7uMm47gGRd02
IIMjUyQebwK7r1GssdL7IhDSdg7gvHV87Py/1emp4yz06sdgkkxlYI9Z4I2nKu+84cvu/h4Z07+O
TNdG2NGLMyQWr5vLWJiI1U6orkklRtDnYeboDJkzak7LNbgCLF/jqcKdzLnbZz8Ledcvd1meXsgN
gh9m5oP3yCUNHv5VPs/OUfxvTED5L0G2zt8PTMFyhgClJb7P7aWedtXEIG3701rTuQvemGyIcHlC
ngr/8oicH+K9QT88gt+Y7AKZtUfOt+PjMlgRdDBU04ZlxBkKGRjFao1eULi27NEIuGmjOHD2Dbn9
nUlDhj8DG4RhVS9Rqmw4HbnSj0WPtmquYVf4VgT0av+wbx6e1fM6jSNanAv6GsHEcySEwj2oBaSS
1Ax6M4OuwX4mOVXVH9BScuHviPS83vHdFmkB+hL9OsUNrD1d9udW4joReTnMfPpcotxO6qsPKrmE
MDW1AB9xj53ooYO3aIdBY9rIfuAE8Ih+F0Q0flqpPmvjdUIgFxGnQxw6+ciJZGKoYhRQu7czN1SC
dVrqe/AIehExQdRI6VXtK1ovQc6AHMTMW6v+FulyimYu1zvoENrc6VCIRwgAbFJAtxxo6FmES7D9
pA8s6GXA/lt9TcAxiB0bElCtcBitjZVP9JEGFy31G8ntZ43Bfvp/4Fq7MsGD2jPhTOcpqFTFCH9K
QiUZcITt142U9YxSCaeVI1LyetHE2ShcUUPifCmUrwjke4SffnvxqAvulGSjVX84aa7Gi05CDrca
RX7USYLD9RTkrZGl5AJU/I2umrWR2/eyJqFwqaXnDDzIoR9JXBldb+Ea3AI2ddIYRxiYDEiGUsCP
4GRKXSmjHAC9gnA/12mc25Eq/mwGaPz5ETSlJy5OqP+VqVU5y8iqLDadV5PhVS5FF0R5vgNodB4s
ZCTRK0Oq1Gbh3gG9UImgT4hI66AzggS3VyKALihByt6whyjdohLyOWhLthZ/iV59otucGzmjuIcZ
te5Dn7cKSdoHgEfj37uk3wF3PCZSlP2ZR8jMReDceB/K17I8iRud8idfNvFlFXtbJSnWhBkfEV/O
6WwuDxKfHxKvSM62PGSbGHqVfoFYpZSostUIY+7WWYWbgynS9N1zsYaM85c85iLvDqqvxYWpIJ5q
hPdKJDuSFaMUXhMv8RIapn/AOYCT5lZqKLEUNYBgaaaRmks6V7HLtCwOAWKnr/wFWrNdXiXvj7vr
nrbzQQ9NxN3ijVVi0q1Xu9F1S/f/SbTcA2DCjT9H6YFQf3MJMwRpxL3QgFwEJTXcvXEPFooQPBqQ
n8lKQKS+9MX1dENmCuG9qj8/pJ7I7mmNSaXuSXOmszkhMnyWKf67ihLFBPFIzWofl8kfeuVx4kbq
tihTRQFuWRoFfIomk5FCTe/DO2dusEhSQZpzVUI5nIDturyOD+mahdFed24qE3CMjha5bTwDkLAs
0a1WwmM6WfFDSZeZRKOlUTL/UB5U1AZTb20absqc3Z2LN/SWzlWMDKIrIkm5db0QmA0atqJ0UVEp
s01ivMbe0eYSZKYAQIwINk84qKKtutTgVaRJrglz01lKo8sjAquOUzX2ON7DZg3NSiVbaht7fguq
byaixwJdJ4YYnC07gkyWEZxWby+Zv6vFyH/g5GAOwFVrwNvf+Lf/EB1JHeF9X9Pk2eyEqD5CoPDB
EgMeYHU28jhmfCkxN9AHDxm5s75anCbWCWDrinq8eB2M1RP3ToJIOQCaEzFPjKgWxGUyZLD2Eo55
GeONx8fyr9Tl1xcEYD/O71TYg/DI0wYQFyUnwetjxOMMzf8YdTz7WvMZRmIhBSVODHBue2tovTiC
PWzNX83FP/eT9bBmNzHZrSynn/jXfMj3pilZ2yakWhc+LGXGPI7biJoz2E5n2ejs9+L5MLZ+6oTt
2y2mi3/66Ury1oeoB2bg71kcfU78OAeXyOEabhK8x+AWAt02r6mF4aSt064Avt42AQuZv37vDJrs
+kCNEv4znCZu/cvzW+2CImYKit7HC7S7uU9gWn0b1mTpMXD8kOgP9QYX109lkViGyD36FUPMNY0k
x2vx6DzsNb5wfoNujN98DHf49QTHDf6elQX8aiSa+P8wCS4DW8YTgT9dXV4HhoP5+bf4y+HFeIKj
wsoQ0jQEGVdy6bOmpHkvW2SVfCRg+4slyGoDL7AffMdXPuWIkv8kdrzhZRpH5dGevlaDoY7tWul9
7qDoH1fNGR0YnL1nsqk9xn7CbNF+RVw5m3v8zcQpt0yXnxd0uGJYyD0CxvAamwYzC5eLxR+e5PPd
cxi5207mSjtF/1TgpmmrM2cOYIIzGKkW4DQEsvO3PZfYlMcaTQENUOf5AeV659eqUYecCtIHawzj
TLkTBoPbpj+C5DpohGMOWQydg+hm46BC3iA3PU18nQ2KUl4IR4XhH8BkAyRgvDcmUErqQkpiA5lt
Y836Wy/ZyhPs1iu/XDAQ5vSHeExN9D38Fz5vzs/TKfmSX/DSCE60VF9i0Np3BNkYGiuK72HZc/GK
6K4nMnCn2aWOrI3xrg4aC0WgJlOg81U3sNbSi6hqfFGrSoQiTQQ0ldv6vIly/bscgN5yv1q7WuBQ
csJZn7uxRs2dQ2QOU5SzYAHrl2tSvQPJl+aujrlgBPs3A4ZdubIt2KFA/1RVxdSbfm33kUPn8pOo
dykBS2xsFTsvhmfpT8s7eX56ST3Eqov0jKLfDsLwRFJ+R5nTlzoSzNCRkXpCMIFF873Dn1tNJkr3
/DDjk6CpJvxtfOTG9pEGMpVkPrB6Xp69z7NLX/EWDUXf/PoQoJWtYg7niE2RtI4HZ4TKhj+a1utU
LzhlnoB5POlrYF0VJhEquFAoZwyNZbhRmZ93GUqT1UQ5pgGGGAIAtZ74XQ0SJ51x+Z0UwoDm48MZ
eXrLH2Asqp0jANLGIJF0S6QP/jIgkeLuG8Cn0xPR0GPp4bon3a+bAt+9oZyRoAGejxjtQMdX59ig
gUTnCF0p/Soa3j4dlUZnwJOVt64CpagWbDc/oGT07JzFEswRl5h0ModY8LHpG4aG+kTD54mjgxvB
s3AyERsH0FM48l+4K8PsQrxPK5zFo/h0dp5I1sxAzoVbzAbDyuZZxMA0/fWYtEiIpzLkvh2o4pVS
TJcTqgRrQ9uYMp+aR1Qbnj1plfVKNikxwywoTHKsTla7Mf3bQ3jOeoJQFc7wJF3dEByCeo4IQjow
ABEAtI7hvMjVkDlNggB7gWyFWmpl6d/ziX/qMJ6HmP2g9gOCjti37G2msVoQwpdBxsbeZ37pWkFo
WthFAQJy92Xbn+SnJ2SusXII6x3KmCr47JOns9gOePredHKyQn5xhqLmlMoelA0fHJTeZb2PU45+
E0vmLlbdld01cXQ/cmSdallkSUjMzzNmuO8zYQE58hJiheydtzKSN5C42nlhFmKaM3behKx++9JK
+jx5HevSJL+p7+k8PW+PY7pjpoePY/YnuCAgesL+zQRN3mdc+e0LPmllEnSay0g/BIUYvJryqEZk
i+DsOuwERp+nyvxUDkoByKBAi9QGHJrVuDIDh1UgOLXRAGi6zKrzV7fsIzvjT3vf/CMI1Fhf0E7u
C1mLPU1sZULa15r1JiTBGxrwiSZWJHurBP+QQkhk4b+zatZeitHns93H5K7PG86+y+OVR7XhV6gi
BxTLvm+yTKnYIMt1vlvBwdZFUs7dp9B9P0xZ+cIefOSqnNB/cFU1d5D08CTWlIAfWFQsHnoPLEjf
xAYpPEezohxeUbf/ypDQPvGeK6YKblgIxsYkbeSe4N8h9uREaHHmwlIu5LpX0xwC7W2a4FVQfLH/
YHTL24IAvzXgARzEl8lYlfX0apvJF9MtWnj9owjEi4AtzdZxBqvBoLAqmT9ji7odMCzqUnV/3guU
1QBr/eSCwrq109+y6I2VjOzxCPt2lkcDjCSapaa6Jhkzc+YxaVRhl3DyiUIwo56iiqaJqy0gF7zE
nJh/3Usenv1IRBpQXLttuuYwqoHBmsCiYlqBkCnVBEcJ2Z0lIXp8pdVl33ksFrNnR0RKm/TV/33y
BaDxlxh6E4UINLKNeQXNLvNoRU0t5hDvLjZaXmEd/N4eLrqdftvckvNDx9E9xgcDcCvkQPtJGQBq
rOnzLn5wLqOtD1vXvI13vZ+UwSBD9oEHHEhzl/3kpfb+ZeLmg597J7hfPbEe9hLrIND732M6rXMr
yAVIZ42ecJUNgsG4cXQ0pnF8s4CDdvpfhbl88QmpCgVfIqxGWY4P3WDylvPgv6syj//AF1hryv+Y
5rHYdMRynySRQW7zK7kamMOQt2cHesuTvvkwNBWAW7ZA274icND+tsrcLWJl88b4KI4WFjzPzkD7
uhYBtkk+OtoGqLJ4givthd5uOB65RuYatXegvxnYqC0MAKpW1cL9Nr0Z1XkgPg9XlspDkp/3T55R
wMkw59M9xd2nhy0afWulYKtRLgrAgnnuPXAg5EImmprP1RCdu/BkMy49EKgaEqKWQnY4VZPPI69T
ujgzNocnwCrAgbJ+Y979qe5QfePZcs3G91k2WueNqXhXK2/ThN2YIUT4NPvm3Wj72EMGwRg5lboY
1uzDCuTMnwszhctFMDDsy1wlUl0V9Jo0KWYPBMyeFUdX88suMp2iUdWDfgRMwiCcV6QsnbjuSlh/
mvv+Ih3nusuzL2GRfXB3U1W86jsqQ7Nhq07SIkx5ACc4eA9pEX/BwqfQ/J/H8j/aoJ7YpteMyl7A
SuyM2TuDY9zSKQL0pODMRP/dTWICeMTHbRbXdaWKWydF+8h3V8fJAvVIcpl6O4pk/NfyeT3uuO/E
rhoOn1MT96EM7sqz1t6I46YOyUwDYPDVXx6CaafLAD0q4Qm8RQDRoOC9NTSygo7OnyeHKwbNNsZ3
KR4dreyy4fTJjB8DYMeBIvTv88t9BlV8SnzF2lXCekPvKUNf5FsXAOO3OFgr9BeypGtLNZnI3C+J
UvFZ5cU2r0bbga0vEy+k+Hgi32O3OYMPUG81mAfgvfGgcW5enj1rTbiaq5vYjqLn4T3+g45HJUYZ
ZpUmUMNHe09Ay/4YyEoK+jpxMS6LjEjxMBoKS75jROM4F8VeNvfckiF241TplrFC+QzWiIABoTzE
s/K0hBL3eAqX8S+Qd+sFy5VXVdbv79FTkqL0+Uuqni01Oh/sSRnX6r/wLH62/2NkRPIjnSFBuD+v
8pZYb2zazYgvbRy9DULYWI7A+96iPizDzPS/qfv5shB1rSx+UkKd8MtgJDWpZ0EARbsnONL+hPT5
FkfrMuyK5JMY6UmQka/NqS1ESjo9P06mCXxKIeyxbItgSDnkmwIVHzhFvwsTskFlm0JsvJ8LfTWm
HL2SCgrQEo/2BPb/PRsxGm/9vBDef5hjSVABBDyZcEnVadJQYViWc8gJrIzTcPACHfTULZQHrP4i
R4SOrUkXbPenCZqDx0OrA1SHg+tF2QCKixykmt1sppdgJwdYhcspxu5Wzbs4AGAqCBYHHOir3IB4
pQxJMdJBzbI4d2Ir2t9Y4FVrTTCOap5ggD8RIhIBsqwovWEWUDwJ89WssR0tej/zNjONnmHiNqzA
/crGuXFXxte5HxeyUD0dtGoW6eMsxmvvz/vxwlSPSCyUSHU5WvsTKIi+1tpaqOCjJnEPtnW/gnz7
/m1loXVehdLfLoj/gxazgfzM8cozn7FMaw0BLr1FI5QIb9rdrPZgcK+61f7BDuIROMohcU/bVZbU
WBHegYmtJNiOIzYYXGbh948nhUQmL/fel7Iidq2wHxbClXWepU0BRw9kVKww+E1K6b7g3oHdW/8x
1oDNJhJ01jrsY85PKIXwSHzZ/kT2ZoyK5Ext6RHaYmeUTkPqXoFWPrv7awRO7MC/aXV9zF+8Kpdv
w/bkZ390NplL5a/fBodyMOjoD23of10Rg2K9ptNVs7QWgxDUoDYMqBjp1qE+4Eqgbi7Gn6RUBPmh
cnqzqertpC8svTnO47S/YDvXGRo16CwIDm0aBdryOHvp1iJTvc+4akim+rGXC8od88yxV43KNzgn
yfX68FfjUnB3O7rX4tsPSWbT27JuXZBsC1mAhK4vfyVrN8xrSCgqf2OIa3cfQwBRuMdoJeA8ienT
2YdlISCelhYFDn37HHPwi7ZLhz0Pjh4zRMkLX79mrcBIS6zJnslQb+qFiD9Zp22R91FDq/j5xTeS
MocBWjVwwxIhRIzF7IC4vHI8x5xsCfJA191iEDDt9vBEjAAk6GM/Nk48SJ2nH93pYB8yCEQL2w4x
hzBi0pfQ0Mj9p1JS1TSI1s/66f6K5XQoIriFy0NAG2Rsb5DdhNMpm34mrn2IdiXFz2mhqOTN4y3a
9khQqsV74OLAwmAE4pqZdQSerqtFblUNharcMY8eONd/5iWHSP8NkrPLIHEOKUMykWhcJL+wftXj
+4P0W/vzmthjqGhTqC5ApH8S/uD2J9mYqE+bulj5EtW7en6wGGobcs/AbXXFitbYo1cJ7F6sfZJ1
T2an4CvS0IwFiVOXA5/yVdtM4Zt9Zc4YN9dSA3MV1/t0GyVx2Ov0quGGe4TwmeD31naT3mkBEL24
vqGBJRTfAsi5lv7IxMq/Ce61qaLPSDeNsN+GFML9VWSV4jOOIUyqbH/FEj5BOTF9UylRI7a9QySI
8+/lEL4P3lPoRti2EEqqyormcxHxmabmWnH2joGKsqC3OMeMLUNgzrg5i5K5xMf5M46tF2fVVX8t
K8vt0+Hn3dwc/S1aOgR/40npEGtdflaJU5OdZ4CDhAynSpMVrIMBTR/H2P0Hyy3cU/itQw1+41FK
D4Rdm3V1gk9c+q9/bVykbwLhmJUt6Co0fm0CtedOIHcBvPs5Lx1+wjHFCaKisUSBH7AukYxdy4+N
UYkXgnfXD8nt+/a0jjG0Y9qBvcrM3JDzu/fOGt9REyurjDgRQrjVfAqa3bE7ZQRqT2k+YPyjq6qh
WE6DLKEyYSFVUJjwjLVMQCYW+KE9jWMVdL9kiX+/kkma+8HUr1KmiN5Ltw5tb8fSALPB8mlUmdAj
pI2JqXm4V228sMf+NuZSxQx+5DzNpm0FuUap67QlrszZxuEcV575dzchCJ2YYZNBArqYumdZsBZT
6O9GVOxfx5gIVTc9t4gZElkP89UJa7O6jU4z6D48zNU/BHXz0kbWeX9k8wPZn5eJ083fGDfsyPLF
mA0mUknIbLkyk24V8erjAXobvKzvpBaJkS3lC5AIDBfV8/qYfDRi29QzvRTkag+dXTZ4QGeSsmBQ
NbGMRPWZ0j7qVtCwCVTYqiGClzBoY2GJNrvvEOZ/3GubCp85k3vjts7QFTRtyqvF724cJ8chcXQg
KCUpMfju2h9ABl6EMBPEgyeW8vN1Vb7SQjZWl29jIo9c2LitC6r40V5pNqipO54bNYKmuWiM56xp
OS/g5++YKKVNPmpK6ULqii0vUjAyZnMNGRZKDnHZNsgbOAg9fXEcAHT78kb6t/untxgW7TtfrSq6
DPB0WACG+1kdE9DlOVFZH00lrwon/YotFwkfL8HSwrqBnPFvgLGCVXGLYyZshOGS1jRNzwp8cGby
YnJ05EAWqR3qP2awpei9YHBmNPQYmel/enUVxwsTbU0JznY5on9jbDuBfSRvJ7+WprdazJ7vRL16
APKXSt1ockYyzUX4109S/HWlDsbOO+ezGohDXKP3BpqP3ce2q45QWPWFOZpdXY9nJTPcD/CuQh3W
vyjG3Z4X4NmzDiIhpxeqDcjNG1A+ubG901bXtPs2XmelEcmlt1gJCGHTmCg6rQtT9NvI90AWK/6n
kZLiaOSc4+2QP/KeeEt1HIuKPy1u/lKfL7qeqMr11RQi+Ztld8jvWBDWaVHILdFjSDMIPomQzina
A1Vy37RTOxcsq5U9Rahs5FhBmC0RuLed0Zq3QOcZD2Ct807aTqif3sZcIgGMsu8OsNo1toD/w44H
ha2OLunia4+RB+QKYzNBzv8EO6wgGt/hGdDnBGlyfxrz7Bkq1VX37r48Ex733Y4W5Cu+zlHKooS9
WWcvf6VF60Sab3UcPDsU145d2yJgqHH7fquCCe4NRMHqa1orhZLh7O9/Zd2UKxR+pyYCiRwvxzQo
TerroMCp3+0iun87NXX0qi9LWlT5Lu9692moCO4iVsyHpmZV4x5JcZ7MCKDVGEF+5khol41KGlat
PCTcshJ1JaaBJrMD0pAPBMrpqqrCABpm0qU7j4Ry49E+hzzOANgAExxeuc8spJsHew0RYdkoN1Ci
Lh+s+8P+ljUtpNY3Atx4RWNi6htBvKpPLCBHUkOr7+bd9oMbssOPpmOy5IGsNieec/u6l4/KdH2g
8CKhmYO4rZlmTp+dYKMp5vvrAwgXrVQ/p3KAl/TUa1BGbXoihsnyFAXVn2BHLFVwbJch+e36696e
shY1GA9xph5Qpc+Mne4S/Ve3OvgNnQHbbPPR5EApAEU8WibmBkblErAZPKBIBC90PjU2t7rminlZ
oNCk0uAmeycDMoEAbqNfOAtpZ/4b/+xUBp5xS3CURWCspQFURnNvoMn0P6Mogq+ewlALdfKZOpCc
isqMGtwVPzCEO41m70J67LzmprQHQfkS0RJjX3f+SBKtL2zNFJ8Jxk9GmbmhFURm61nygMD6IRVl
SWo0g0KQJ9eDfIIbvCWkP2PzmmKFRYFmA6uxWTtEKd+lw5SNz8GolOwpJF1cDBV+BtIBgojfXeOj
L/Vpo4d0vyixAPttFkwgQVKGDKo8fGz02j7rEHeOgJKaTWYUs5Lg2Wfv235aZCjg6EJqQYRNdVu1
Ui2iat8qcVM3LXSeoD5/6y9Pg0RCRH85VkIOcR5g22pQrrBES73jKQSfQEq5V7eFLZyk1jmR7H7B
ae8/ryKkfIeo5VfaND8NP1aC2wl5j2Bj6N7N1WdhpKDU5dGIlfyP3BghVQ6/lGGJA0vCEPx16aTl
LalzHtK5Q7mKKSVJVCepQ3rzARmuvsNUENxUkqJ4DKdsXefpLyfc3wiJeUSwBumt/ewaxrcFcBOH
IEXqtdiUKbiPbZFffXdfnTZEZnBEeeKCtCp/NyMpbQAWNJFRxELAGChVaZkLy5AmdJkxbgL5ZbYF
ym6kEx4rMKXmEAhet1V7WKE5xEaDzgWkeZBwVUXxUeOMWcGJCeIVYWC4P1D9zhqh9BCzzd5em281
/vEJ4aovh9IMg+mZbU1MPyVI6jk/QQv4XspC6lh8gaBjz+yKYWo3sxgZEhfpnbE2vgrtLihpSP0y
MA3jzFUro8ST8lA0sniEq43mJ8Q2eXiTDGLmaMkT2hPpTwA7i9loigvj/PnzfTIohPCGlwGrF8CY
4T05I+Yfgg4TZx0Tf+NXBiuNNvIEzm+CfZPGw3YfoSw9r2IcG/1PayvhMOIGAFz04hNXhmMifPt4
PYabiMTc88mJBE4g9PCzXurWI+cJB+VkHipRx2YXwmSfxjdnru4DUBap0r1PWtYHdBBnaQgGEMO+
hIjNiq265QrmR/BWrmyzSrdgzTPmQQkc6EjvtrAW/WzNZTpidTizivzv7p9EJ72boajvbOdmj6ni
FktYltBXtS4QyHEHBsbOppDRk5R1NasWzSeT/KqDjqDmGnVhefrWhVRWIOt9MtzjbvHv4c1cxjIE
xLkNaiSlUpE1vCQPhIuoL4Rqtxm2CNqqR0BmgU92YZV5V/U0+6U/wwox2pL/5iOBeRkGr5HMPvxe
+FgUmJiu1LFDzYNN6wInCVGTncdtcqSJ4OTfpOhUquPqmrXlENw4pXMXVHFpApune1R0DMNhM4yW
9s1K+TnvHTBggpQw/Fwu8zlNT2EHqwDIhUC+YdJ2VjeQNnl9cgAqvSQAofxozA13UynQNVtNZ630
bOG3k66rzkgWQn0iEqyf3RuTM0fl7KKpveyhB8U3hfUv0NfDxnm/y1VBeL2NjzXDTNO3qkhNTbsS
1Kh3mC0sTnJmJeAVzulz4WZXR0v+WfvQneNlX8BaE7Ay3ioNOKi6iyTUK7JrtQwQtk376ItamRqw
wRnfY5wuOtAY3yNBXn0TWCP/o4/2Omk3cxg+9u6gLBJ8vAU05giuQ8HF4uQb07PNIHrSHjkXR3i2
KtVwV3f+bLE8bK7A+837CHEwZgusAgghDuOOq8WwWu731Ntu2H6663Bnc6TPCG5F5YEmNW91GtjE
WxBpsMc2AHCiF8bl22vhvURCUvyUPsLtlEVDiIVYAuDJUG8eBEQ147yR+JtfnX8xdthc02GjLCeb
cYzTq9X8P1hrqv1c5rpb57nkZaCNd34ZOsnRFmIu/68t2tR0BNv+xpqTLxUB+ztsEwAgP0Z43rQN
ZlPK+oJ3C3eEeSOPXaE5aQCq8B4waFQShT8gvTUy3eoMKUMP9meILyxygAeVncHFYZYH+sBq8gmi
+pGzj4aAppEGI5omSZGgX82hDsTR1g53MMX5WMpnPVxxmVJwdTrFeqCdrsmHGlVkcuBgynXefNEU
yGtZXwLl7UnWXKNAd9jhv/ThS59NeI6aij3POrkKTHmbW0S3FP6ndDnLtT62e31xBWHV8jN9ke3m
L1tjkELN9OJBb/zY60ifN/Px+yrEjgYAOZiKlRywsyAAz4Hc3/9+44mOOIZ+OlEmAu8qqe+5nq8r
nET09qS1tvC9Zrs7iLAX9nupdcbFKCf7Eo/u9gYZMtFRpH8yu51FPSTulK4t4IJm0kwEDklc2NUq
WukjFMq93hxnH+f8g0b0kqRHkaOzWJPwo0UJ+XmH1N4OV3YJvBV+t+BLgFxxNFpTI5hZbdLAbh4K
zuebPuRvuwfZvKZ3h2ALAskI8tcKU9SP/kbR7IhC0CrVJNrWA6aJ6J3vaZMmS6cA5DHI7LwpJTTj
rQsi8wORsqT0elEu1F+zKjOh5Nh9toamRdSGgHF2DUf5j+C9yal7qn5J+40vknRBGj3PrhwtICJC
UTxMopU27DsXlyjOABXB1F6krWHyTNpZWqrSltsgkVJAGT0M+aLlD06cVsJvBMuE3ZVR3tXSy9Fp
cj05RbbN+uiqyE6E4TR0b8F29g5rIvdxdD4xzvACFhMm0bNGtzLFVaqrMK3PaVIpZiGtQBH0rdpC
ghnfwrchbXUd1ddSlKoA8z034lXfJzIAJ0e9On4vOz1Ew3QF8p545fWpupHN76LrYL8zn127cPt+
OcAyjZacvrRSMzcEOPBjJze4XdmMyoIjXT/kFbs3L6mGjkIf/rT8DinIL/SeARkYZoKDWDuBB42H
xvNmdDfAY4SvgpX6iUua6F+h2VCtzVnbHfC1PslyT4D0gGGuCrVREIMqdEC+588OMP5ZVQccFLaN
MKs7mW2WGl+5pY0NL9AKB5ZhXgWviGa40mp7rHeNOr18pIGDrLUiezYA3UEAWfnAz86t4HnjW6it
YIOnDDsVHjvuLjwS3aMCgJy/N12S3xFMcMi+KAgrr7tA422lgvHcSLWBvn7Ll0aatr82N4GUCFtY
WYSuxRyx7iQB6xoz6X/gN8tm8KLbe2NmXq+77XUDJ2cnHq5lKp39x1aiInXu5udGi8zattaQ4+g1
mc6jiVmsfboMNeEl82mCskNMOvFThXk5W6ZuxrAYc2vuz7U7jt+woDQnFVfU1d/OXnRmN2rfotUr
EqxCl3xI2lgYXRRbPSxEaXGc6ntoqcxoFZDiHcMXLgIzCWyCUYijeHmjxrQ931lHCMkPCE70MUCz
T5HpZfbt7wz4ZbNzwpfZnXD9vP2wtpqVmUcASTGigD7yQFuvV37MrNAySTVqeiI21Ayv0fMIQQvq
4ur94qnEXl3OACRZR/sVl644NEXvIsBpIFrXWDB7eQmJcy06vgqS1cGicyWc4ms6zMftT1Ik3SDZ
Oo5USRmMzvOITvEliMTGri65rkqvIzC+ZEwGc2n03rmDMmSCAPPk+ideA7dSEoys5uWXUb6GJOF2
DFlU+BDEbY18JNjw+M1sWJpFT67Ya18nBGM2Deuex4FP7qejHgx7lG/ecCfmmdJnQcfFLidOu4Fd
U/XmxyZ0CtBRf51pO1m/mYR/wKMsM5qwMCG46zWFuTO2erpEm4PZCCY5tWVCqORLNF4kXmcai5vi
SEjY9gHp+vYmKCX+NGUTuPre+EcXt/hx6pqvXctJMaKc5gReFWEMr1VCCfrtIc5X5eq/abRSJnWJ
cScOMdwT2GvIh/LxClMKtN28M/nFEb7ErdVtLZ7uzDQ7wG9jhihvV5biZTEM6cmHNhMAq07zgiAx
uh7WNwq3g9f+E8SMUQBQtxSBQwtZ4McHS8M6GtAJYOIF6lxuoCSNL8+lf6xn4vZg1sL8sAvKRmjd
i2Y94yo+PY6JJ6wb84sK/6Svr2ie4KtJfwd1YpY01H0ToQdLZki8JCL3Co8jVCrBUuRQhKRu3clD
lMhVHnxg01f+ikStSYeYUXDczKcmXlIVSJvrL39ZfVH1Y5qBlg1t0weYF1C0FicwVlPt+Nlax38y
iTdif99QxFTezJk1W67GQ8dkzN54uFANM4algGG8N3a7mYhw7FjDv5bxXIInktmK53nj9fiJreYp
3+oNOVrZtE6twq0KG/XBPnKPAa55dHX6D2nTMzN24C/RPk9M+cl2M0KOAlsITVC3LQwVDCsScbon
BWwgiUuo8wzRvcTmLEROByMgJ+Px8KnoE1k2PrT7v+ycq+ytduT1xKb5d0CaHuTARcQADI+Osruj
XRvny2LjETAovkGJA2PJh/aNWbsHaUiQH8HhaBJhgqdYYmt0QEj25OwWpMPmnKU6Mqfz16FQXJfW
jWokqX2ublGza0T1xWPHVQe2RnNl6mRobEBWoTSGIJrnvD6W1AAg1oHf4NRbApfu+dY8gCgoF7u2
v1iB9O4nwXz4cPSh1JI8eimHxKi8Lk5B4ohMaXui3zi8kF1wMKbIeF6rkxkNPLqolKIcStDfmTNS
u9+re7QAicu62coClYbx5LuaXLbNlW3fdSm526OfWJEAevAeIpEUzqQNQAj/UIyoFeQdISej17yS
v/YVKu3Kke9MlrwuUtdfZCddU2LpEala1uaP/GBhMhqyNZ2fDtr5ABNookofRx2OUJ0gghaKaK0l
+lZpmsGFFaAWamzU2Nkq5XMOIqm073kJA1JVeeP33btNfYwiUExkXCalRZjCiK+M6kqfCbakZMP2
G2DPEDCDfcUndaDzVNksNC+Oo3ssLW9ovOH2w5ZSOsFQUz5Fx43HMd6DQ4CMswQRnAxDEXS3qoma
Zv+bUl66zJCXwiafwSKiungWko/79KCCGHymQbocMHPL8iRLcB7YIdh4MJU2LZC59qfEDRtV098F
j3ehNX8CcYys0ZB8k5KtuF5mkFnDRL0hJ7T9Gs4UrjBZpRkrGSJt9fT17WOxhP0LXPffUMH1O9kM
QMgsgN6xFRDe5Wx413FKFXwR7RLTYf5L6FUbaNs7N9vnZEy2yXHN0QCWJRIgK+O1mLEhdHtkAJO8
UTOI7a7qsWXsZVakpQnDkHJp+sOKrFhprh30pbDMTWOZXUoHQyp5ZNmeuYRMEwP1148Zss5yIcgm
xFxVgiHY426Ml519gvtQPeBDUvv1GMNzixCrOvT3+1kmg0E/+s4LcCgO+qnv7nJpZzpmq2brr6Xk
wDaMmkrnEv2FDqpip8QnX2f32tRDWVuGuY1/410u2b5TGI2R7YiOB94cSIS6GMiu+cJNQKhP4T9r
u8MAEOQNRilpHhehw+Dvo81ZR57Q6R9IZCT/hDoFnIv0qDFlMGCSiUZN2mQMZ1sn9etFlSMj1+6i
Nh1AOLnFZkqWsnlNk6zT99laGWKFj2EErOw9/+2GsoaDl5PxhOsU3EzcUjAsWY1CaEYI2ovktvLv
nIDrDE7XCjtQapq2PitetkkxQc7FMOococBkZTndmEQyY4N71pqtr/reMoIewI3z2/nRjP0r6Wtl
AGECa9AYBYE3V4qQwZdtqX8wCtVISdvKfK/mmqWYaOs2yf373Rd3nhIvFJ0yda/Bs6LPo8Z01DJE
brGCIGi+joVRZKMmHcJPdEgji2kueaQ4889spDk7xDF+67ebPaj7Y4/3CEEOWaKoQ58El8lupVJS
rKekfNmEgoeySVtSCCrx7RHbggAP0w/0UDSHKBVYPkBKmfgpwK5vTD9BgwK8yneqVW1q9BkVBx/s
sV//4z8IFt6Hx9LSh5OY6YQTlG/4SO59N7cRvj3570VHWcQgLMRfbSLCQYsFimOg6Og812vxYbKs
FpZSX/Y6AjnnJ+c3GrhlHHeu3MED0tDBSh+DGhnb7eIvhcI9BcviIFbgOEDxphfho5cm+gXf8dNm
0pOI0ky+DYfxTs0S0mv0kEcdu+L58pbJSPnruRBaAEYWJeY6zMy2Iz5rENumbkaloRZ85LZ7WQNl
0/xjRSQjOL8jFHpcA28pMhnMBiTbmI1w5z4KmUKZIP3bqXOroY3O1Qh9nOCOQwiAS6svYXvjU6Cm
eWUZRYJNP/kGOUCZfvQ7mwQoy4TqxwlpxkLBgKTI7auwHPQxQNqoXibvmGxk7G3iDrsM1BoVB+b+
bM06g+bxa2lPN2D0Ho2Xz/cEh9GEASswo89xB6uVLDUFZtoB32r/2K2RgvOJPjdqSrTFtqfqXuXD
D/7sEjd+qrNs0UD08t6dlenU7a+RDyhIGN2+RZfcu2i6UlY0iN2RYUNvMH+Uc6bEqCMDU9Jldzms
MksMg1WpYtTETQXhKIZe+M//eAYp7Ic8D2u/RKwkHBRl96y45xTef+WoN+gdrPZd4W5MsVAUUxNk
6gdcf+y2uty4vXvGpbHGtWIl2BbX2k1YJXCAQ+UyHcfxPDfqJfxHhBjYDcVbvdTYoptMDVYPNoKf
8/mPl/k35/tO37Mrn+WWzMUJ54bUbRtUoMIk+ywM8FoO8rAseMxiXcfw2lftVUmLA67HSV9U/D8e
fVDhCK8yeWqU8oFzGu8EUrgLN5kT42jwElFE2qGUqcxCs5TzewGEnahBBbFquMELVyh9by7Ll+NJ
BQwVMtbXe5+M1c7i/Q4hnQQ3sSkoTroOvoycx0qcLTgSFtVHMOYqKw4NYqP3HBfW/K6WtpnJA11s
EhV4SfOTpCbGGSAuXcT9qAlkVijpw9R4hZTouPy87DZmmdHbzsablse8uY3PWj9mhgBW8FwLo1xF
AzC2cAsvMOb135N//XWL3GicoOBNJwUH+b2G5GssysUUCP4Z6GjnbVNYEuLd2srnjDuB6tocJzii
sj6rgMShKY/pND/e6To1iKVZ1ur7e1u7oBqx7rvDmv8r3tF07YLmPS0iVhXrD67nh1ufZTNZNCC/
9DiSjdj2/aGDFwYMKqmr1zBIeGWLC+cTr5uUvDUu8Cw84Mu89CZXdogOow5LCgJx/G7xHBArtOP3
pY2sIY22gvHQMIz7CTbxIXfs5/bKIPbBSiVktr/taaKFwgjJgaaqVCjLxTbJgluPvHB/nktzuBa5
r6xS19QxpPnPXZa6fdqq1KqLePHoZ4qGqYaEK4U7aG0vEJhkpo17DM9u05Sc6xz3knUTtZ2n142H
iW4s8SVSwVsMwYSiUeprGU+u5jUwPDrWEMjYaWXSq2cN/nQUk77fPUTJ16OvcNL474UcXAdosVOT
qLEJxAiRGiZd6eMqQlXGxv/uq/Vle4GqPqpK972s0ymNrvBAo3eCx/rIxOTPVHYwLO0DI7eBpPpO
jHC3LzbD/YVMHyVWuCWJoNFaDwPJVvYpARymOBMrGXooCEg1YOghWQS5s13emFlFwY0k2tmN/VlC
kjt32jEawE4zfe/Wn/rNSxVNaBuP5jOtzgyy+hq7NFMxfiOUxo8rMlFasSBDdSnocSzR7x6LZHRE
o0C3pLeqVDXSHkwfcgo1Lquho4gGVy/NL8ythYRHqR1V1PRot4nx4V6oLV4VmyMYwU3J90HaZ0o3
D82Sa2dwnXE6wtGaydj4EwI0Bd9R2h+DmsVwlejrQNpM05bMMEMDORJxsvdvoxINa33W2a7IUxVo
wh0wIEepkm3e4w+fZrzN98CESwi2GZRfotsSQI1sGaJkvr6q+++qCJzWNEYi7MR+Zz+7i2xN09e1
hW9O03EzwwRGUXOmKwSJNyCwV+aobxeJahBVMxei4rEm+72btkOHguZUWcakjSIDBviq/FfLvrsm
9zrYPwtS6O5vB9IOZeHMQbWw9cRswhittXufGcSY6ByFb6PTUuz2C0h2k72IgWgsPtRCnrQjCTeA
wNoaf0jcJzxjNo9QtKRiPtikyyD6lHgCsOaPrkb+o92/97r7KPVE8dIwHh5Sk0unJBC14eyhMWR4
0Wson3znbh1nRXZpzFxWIEA9MUOywjTp3NptQQlBeBryUX84qfiY07jjkeOulBUcfWlRJeJc9EiV
P73uZC0+iDPHIjDI9SgjAApvoUtNqQ7gVt+pmnsbmJvd3WlcPgBRFCyCSRgV5p9YRoaZRvFN+ABa
/mbBKrp5qf0APwjt1p1omYLlKxlpV6pfM7MG++pbPeoo3vjdMOs2RwOH5nHBZtAPs7ODtZvOsISA
SCAdCuO2PuAG8ntUuboXj7yWWsJJUhX3KaIVxxyifhE04xxDhNZBl/EGZMrXYGB3xBaUaF1ACIaF
Jkvmc+HQuy4JLILvls62TuOWfQm2X8SRNJwS0ldAqIFDuvSI+3RiiM3W+qYdESuiTfbCD1UtrT+/
Rb+pc8/1Tog2lYgwS3gPahs5c/Uj+BjI2RlCxhDHD0LfEhMeSySCmCc18bThnkBqr79VWXIbmpqJ
bFI11KMelVKZxwq26fYfAFjWmRUs8DLKeSUhqpP0G67yoi6zPxpEqrBKg9oTToahLMPX4E1NlsYM
PbP9oYMLqVNdPXwOhW++oKA31GjJDmD2G93x4Vn3GnEBOMgfUKYgpdSncwMLXCrZCsdOd6hbPgSf
BQRuBmz4Jp5XlTjUyWy0xF/9/zC2EWAKj8WaX5Hm/gjLoz0muy+/PX3AsqOgeYuBpV1lBTLVymta
nu73BiWsN5REAqEiero+rQyGmWXuw+6aTBhU/tHxhRd/VZhMRhygibl7g5mSrQz+Yt6ytCvI/xiV
H0Snt4SX4Hc/+1FZTVCP0lZJ8nSU1Ek1GfxNSZyg3PmkAEgPiu0fXdZkaIFP5N/PmZv2u6YNajb1
Y4BWK4QRbTsXRXtU4/JN9590yKMTFZiL9in1J0AqK07YQ585WpTItUxkzQGPTRbKCKwvK7irbB51
geNv+rOsGSAPZ2gCKpVLa5d1OJcLh3+1it3hHbNp0cqOrrYyLGAfaMrsY5FAoBN+IHj/ihn8vPMK
VsX0AHigQmmhbbo4KJtHI1Y/TUaDqV6ps0oaaCiibAiTyOJpZJhzskFQ4NO/RarISbbBRbfghAeK
JOZBFEEMqIvSML01UX7ml4HyoSPuh/BHw6OUQ0wC5o+UaAPE4SR59UVLyI4fIuoqgK4eC7HK3GQZ
X/ZB/ZRBYBXvwTmal5gNcb1iOGprgXIjyuIxIvw9DUSCMVAsUj2qDK/bBMyzKjBmprztfkANpxRu
vYHaVOp4EHwMRkJza/z6XnA0NwlgGzCwVbr0Nvx55CJU0sTfmSEb2z3NydoxNIEBH1Sc3O+DvldC
Xc7J7U+rUq7LbOqLvCtGQZLe5JFIao8WRPiHWtVYxhnd/uALg58MMgol8gOHF1dfljA+CDTG0JE5
S8LUSynyh3BUkHpdIxQ+ulNyDopKeN6Gx0wxTDNepOZWIJ+g9AOw7tzRtzppwCL08eVl5lx7y5bW
GPb63AOVmfYcewWxRv6k+UjR6gqU5o7cSRLzKiJ6YLZwprKnZbdRRRsBJregReYvFV4iZT6oymWV
aKIovaqFvfh9VOlY34LlU4hYFQUxQWKaBelPekDA1RchyDEAM14Iv0sKAZkImZ8U0t/VIZvFvyLe
Q6fIRD5FlpIcDylPyQu0prSc2Ott+ejlmiZMxYO+g7uuxLj9CBzhiE0+Bnletpcn2ECbqmVNTr/j
zbZc5g7LOTWQJqpfiniaSqYPhQGm+WpO5Tn01ZJ5UBNkL3vi3kpnmGYKOGAuPo7S4QgW5OTmbCtd
pJwcyl9bkVE7eV41iQMOptiuwhc1O1b5ogWv3J+NrF9aYgRkc/aEzVDdcVLUi1PC9XsHl0i3jqO7
blyR0vnQEthBUEdGDtfni/m0lY6aJbf5P8y1bRmCwg+GWJxrOM6+ySdRs+vk0roGuGRAIVg7Uf7Z
DRJ2ieuyvz/SteONMrAdPsSp+pjQEkaxSzWIusHWLt/eNKifq79pZc4nGRLapzFKxElJjSJpJT00
Wu0PCYr6MepSXC5o0oHwrDb+A1EAbSUKxjhBpt1eWGCeyF8LiD3DRflSOlsuC6TXlM1y5pwjnpGJ
lP46+FgalWlrx7Th0VU+JE9sB7QFXAi2LB70PVFG5H2q+d/n6eXOHZE3SG+F6UxdwsgDB2ZcSYIF
Q+Q6FY9kErAW/ASKDOQ/C66FOidykT4P8LUe0qj04GYrIZAtF/+aXzPjHIPd5VgKIH07Y7wn4BN/
oV0OoM0bHlhdgsKd1rz1dRpO2H9c6jc6IQpogAWKqRSuw2BI77OPBiSHPbo3v0r79wmAl7fMBW3f
BrV7r/vWTdKgT1NGNXZlIlF9EYGEuMG3giLVKqdH7EXhhS4KOcCEX92ijh8zomVBtsvg6JP3Rrsu
3V+QYjrfGuwiI5Y04cIKbKOsfX4FmwUrj+2J22jdZw715Mtg9cU1z9NIOTtVnczqLLT3ifzm/Pav
p1UwTPJQFJd0qV69R+rm0OWh6Eficpim8QLAjt0itu5JeXg=
`pragma protect end_protected
