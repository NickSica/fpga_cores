  localparam LC_TOTAL_PROBE_IN_WIDTH  = (
        C_PROBE_IN255_WIDTH + C_PROBE_IN254_WIDTH + C_PROBE_IN253_WIDTH +
        C_PROBE_IN252_WIDTH + C_PROBE_IN251_WIDTH + C_PROBE_IN250_WIDTH +
        C_PROBE_IN249_WIDTH + C_PROBE_IN248_WIDTH + C_PROBE_IN247_WIDTH +
        C_PROBE_IN246_WIDTH + C_PROBE_IN245_WIDTH + C_PROBE_IN244_WIDTH + 
        C_PROBE_IN243_WIDTH + C_PROBE_IN242_WIDTH + C_PROBE_IN241_WIDTH +
        C_PROBE_IN240_WIDTH + C_PROBE_IN239_WIDTH + C_PROBE_IN238_WIDTH +
        C_PROBE_IN237_WIDTH + C_PROBE_IN236_WIDTH + C_PROBE_IN235_WIDTH +
        C_PROBE_IN234_WIDTH + C_PROBE_IN233_WIDTH + C_PROBE_IN232_WIDTH +
        C_PROBE_IN231_WIDTH + C_PROBE_IN230_WIDTH + C_PROBE_IN229_WIDTH +
        C_PROBE_IN228_WIDTH + C_PROBE_IN227_WIDTH + C_PROBE_IN226_WIDTH +
        C_PROBE_IN225_WIDTH + C_PROBE_IN224_WIDTH + C_PROBE_IN223_WIDTH + 
        C_PROBE_IN222_WIDTH + C_PROBE_IN221_WIDTH + C_PROBE_IN220_WIDTH +
        C_PROBE_IN219_WIDTH + C_PROBE_IN218_WIDTH + C_PROBE_IN217_WIDTH +
        C_PROBE_IN216_WIDTH + C_PROBE_IN215_WIDTH + C_PROBE_IN214_WIDTH +
        C_PROBE_IN213_WIDTH + C_PROBE_IN212_WIDTH + C_PROBE_IN211_WIDTH +
        C_PROBE_IN210_WIDTH + C_PROBE_IN209_WIDTH + C_PROBE_IN208_WIDTH +
        C_PROBE_IN207_WIDTH + C_PROBE_IN206_WIDTH + C_PROBE_IN205_WIDTH +
        C_PROBE_IN204_WIDTH + C_PROBE_IN203_WIDTH + C_PROBE_IN202_WIDTH +
        C_PROBE_IN201_WIDTH + C_PROBE_IN200_WIDTH + C_PROBE_IN199_WIDTH +
        C_PROBE_IN198_WIDTH + C_PROBE_IN197_WIDTH + C_PROBE_IN196_WIDTH +
        C_PROBE_IN195_WIDTH + C_PROBE_IN194_WIDTH + C_PROBE_IN193_WIDTH +
        C_PROBE_IN192_WIDTH + C_PROBE_IN191_WIDTH + C_PROBE_IN190_WIDTH +
        C_PROBE_IN189_WIDTH + C_PROBE_IN188_WIDTH + C_PROBE_IN187_WIDTH +
        C_PROBE_IN186_WIDTH + C_PROBE_IN185_WIDTH + C_PROBE_IN184_WIDTH +
        C_PROBE_IN183_WIDTH + C_PROBE_IN182_WIDTH + C_PROBE_IN181_WIDTH +
        C_PROBE_IN180_WIDTH + C_PROBE_IN179_WIDTH + C_PROBE_IN178_WIDTH +
        C_PROBE_IN177_WIDTH + C_PROBE_IN176_WIDTH + C_PROBE_IN175_WIDTH +
        C_PROBE_IN174_WIDTH + C_PROBE_IN173_WIDTH + C_PROBE_IN172_WIDTH +
        C_PROBE_IN171_WIDTH + C_PROBE_IN170_WIDTH + C_PROBE_IN169_WIDTH +
        C_PROBE_IN168_WIDTH + C_PROBE_IN167_WIDTH + C_PROBE_IN166_WIDTH +
        C_PROBE_IN165_WIDTH + C_PROBE_IN164_WIDTH + C_PROBE_IN163_WIDTH +
        C_PROBE_IN162_WIDTH + C_PROBE_IN161_WIDTH + C_PROBE_IN160_WIDTH +
        C_PROBE_IN159_WIDTH + C_PROBE_IN158_WIDTH + C_PROBE_IN157_WIDTH +
        C_PROBE_IN156_WIDTH + C_PROBE_IN155_WIDTH + C_PROBE_IN154_WIDTH +
        C_PROBE_IN153_WIDTH + C_PROBE_IN152_WIDTH + C_PROBE_IN151_WIDTH +
        C_PROBE_IN150_WIDTH + C_PROBE_IN149_WIDTH + C_PROBE_IN148_WIDTH +
        C_PROBE_IN147_WIDTH + C_PROBE_IN146_WIDTH + C_PROBE_IN145_WIDTH + 
        C_PROBE_IN144_WIDTH + C_PROBE_IN143_WIDTH + C_PROBE_IN142_WIDTH +
        C_PROBE_IN141_WIDTH + C_PROBE_IN140_WIDTH + C_PROBE_IN139_WIDTH +
        C_PROBE_IN138_WIDTH + C_PROBE_IN137_WIDTH + C_PROBE_IN136_WIDTH +
        C_PROBE_IN135_WIDTH + C_PROBE_IN134_WIDTH + C_PROBE_IN133_WIDTH +
        C_PROBE_IN132_WIDTH + C_PROBE_IN131_WIDTH + C_PROBE_IN130_WIDTH +
        C_PROBE_IN129_WIDTH + C_PROBE_IN128_WIDTH + C_PROBE_IN127_WIDTH +
        C_PROBE_IN126_WIDTH + C_PROBE_IN125_WIDTH + C_PROBE_IN124_WIDTH +
        C_PROBE_IN123_WIDTH + C_PROBE_IN122_WIDTH + C_PROBE_IN121_WIDTH + 
        C_PROBE_IN120_WIDTH + C_PROBE_IN119_WIDTH + C_PROBE_IN118_WIDTH +
        C_PROBE_IN117_WIDTH + C_PROBE_IN116_WIDTH + C_PROBE_IN115_WIDTH +
        C_PROBE_IN114_WIDTH + C_PROBE_IN113_WIDTH + C_PROBE_IN112_WIDTH +
        C_PROBE_IN111_WIDTH + C_PROBE_IN110_WIDTH + C_PROBE_IN109_WIDTH +
        C_PROBE_IN108_WIDTH + C_PROBE_IN107_WIDTH + C_PROBE_IN106_WIDTH +
        C_PROBE_IN105_WIDTH + C_PROBE_IN104_WIDTH + C_PROBE_IN103_WIDTH +
        C_PROBE_IN102_WIDTH + C_PROBE_IN101_WIDTH + C_PROBE_IN100_WIDTH +
        C_PROBE_IN99_WIDTH  + C_PROBE_IN98_WIDTH  + C_PROBE_IN97_WIDTH  +
        C_PROBE_IN96_WIDTH  + C_PROBE_IN95_WIDTH  + C_PROBE_IN94_WIDTH  +
        C_PROBE_IN93_WIDTH  + C_PROBE_IN92_WIDTH  + C_PROBE_IN91_WIDTH  +
        C_PROBE_IN90_WIDTH  + C_PROBE_IN89_WIDTH  + C_PROBE_IN88_WIDTH  +
        C_PROBE_IN87_WIDTH  + C_PROBE_IN86_WIDTH  + C_PROBE_IN85_WIDTH  +
        C_PROBE_IN84_WIDTH  + C_PROBE_IN83_WIDTH  + C_PROBE_IN82_WIDTH  +
        C_PROBE_IN81_WIDTH  + C_PROBE_IN80_WIDTH  + C_PROBE_IN79_WIDTH  +
        C_PROBE_IN78_WIDTH  + C_PROBE_IN77_WIDTH  + C_PROBE_IN76_WIDTH  +
        C_PROBE_IN75_WIDTH  + C_PROBE_IN74_WIDTH  + C_PROBE_IN73_WIDTH  +
        C_PROBE_IN72_WIDTH  + C_PROBE_IN71_WIDTH  + C_PROBE_IN70_WIDTH  +
        C_PROBE_IN69_WIDTH  + C_PROBE_IN68_WIDTH  + C_PROBE_IN67_WIDTH  +
        C_PROBE_IN66_WIDTH  + C_PROBE_IN65_WIDTH  + C_PROBE_IN64_WIDTH  +
        C_PROBE_IN63_WIDTH  + C_PROBE_IN62_WIDTH  + C_PROBE_IN61_WIDTH  +
        C_PROBE_IN60_WIDTH  + C_PROBE_IN59_WIDTH  + C_PROBE_IN58_WIDTH  +
        C_PROBE_IN57_WIDTH  + C_PROBE_IN56_WIDTH  + C_PROBE_IN55_WIDTH  +
        C_PROBE_IN54_WIDTH  + C_PROBE_IN53_WIDTH  + C_PROBE_IN52_WIDTH  +
        C_PROBE_IN51_WIDTH  + C_PROBE_IN50_WIDTH  + C_PROBE_IN49_WIDTH  +
        C_PROBE_IN48_WIDTH  + C_PROBE_IN47_WIDTH  + C_PROBE_IN46_WIDTH  +
        C_PROBE_IN45_WIDTH  + C_PROBE_IN44_WIDTH  + C_PROBE_IN43_WIDTH  +
        C_PROBE_IN42_WIDTH  + C_PROBE_IN41_WIDTH  + C_PROBE_IN40_WIDTH  +
        C_PROBE_IN39_WIDTH  + C_PROBE_IN38_WIDTH  + C_PROBE_IN37_WIDTH  +
        C_PROBE_IN36_WIDTH  + C_PROBE_IN35_WIDTH  + C_PROBE_IN34_WIDTH  +
        C_PROBE_IN33_WIDTH  + C_PROBE_IN32_WIDTH  + C_PROBE_IN31_WIDTH  +
        C_PROBE_IN30_WIDTH  + C_PROBE_IN29_WIDTH  + C_PROBE_IN28_WIDTH  +
        C_PROBE_IN27_WIDTH  + C_PROBE_IN26_WIDTH  + C_PROBE_IN25_WIDTH  +
        C_PROBE_IN24_WIDTH  + C_PROBE_IN23_WIDTH  + C_PROBE_IN22_WIDTH  +
        C_PROBE_IN21_WIDTH  + C_PROBE_IN20_WIDTH  + C_PROBE_IN19_WIDTH  +
        C_PROBE_IN18_WIDTH  + C_PROBE_IN17_WIDTH  + C_PROBE_IN16_WIDTH  +
        C_PROBE_IN15_WIDTH  + C_PROBE_IN14_WIDTH  + C_PROBE_IN13_WIDTH  +
        C_PROBE_IN12_WIDTH  + C_PROBE_IN11_WIDTH  + C_PROBE_IN10_WIDTH  +
        C_PROBE_IN9_WIDTH   + C_PROBE_IN8_WIDTH   + C_PROBE_IN7_WIDTH   +
        C_PROBE_IN6_WIDTH   + C_PROBE_IN5_WIDTH   + C_PROBE_IN4_WIDTH   +
        C_PROBE_IN3_WIDTH   + C_PROBE_IN2_WIDTH   + C_PROBE_IN1_WIDTH   +
        C_PROBE_IN0_WIDTH   - C_MAX_NUM_PROBE     + C_NUM_PROBE_IN
      );

  localparam [2047:0]LC_PROBE_IN_WIDTH_STRING = {
    f_bit8_width(C_PROBE_IN255_WIDTH-1, (C_NUM_PROBE_IN > 255), 0),
    f_bit8_width(C_PROBE_IN254_WIDTH-1, (C_NUM_PROBE_IN > 254), 0),
    f_bit8_width(C_PROBE_IN253_WIDTH-1, (C_NUM_PROBE_IN > 253), 0),
    f_bit8_width(C_PROBE_IN252_WIDTH-1, (C_NUM_PROBE_IN > 252), 0),
    f_bit8_width(C_PROBE_IN251_WIDTH-1, (C_NUM_PROBE_IN > 251), 0),
    f_bit8_width(C_PROBE_IN250_WIDTH-1, (C_NUM_PROBE_IN > 250), 0),
    f_bit8_width(C_PROBE_IN249_WIDTH-1, (C_NUM_PROBE_IN > 249), 0),
    f_bit8_width(C_PROBE_IN248_WIDTH-1, (C_NUM_PROBE_IN > 248), 0),
    f_bit8_width(C_PROBE_IN247_WIDTH-1, (C_NUM_PROBE_IN > 247), 0),
    f_bit8_width(C_PROBE_IN246_WIDTH-1, (C_NUM_PROBE_IN > 246), 0),
    f_bit8_width(C_PROBE_IN245_WIDTH-1, (C_NUM_PROBE_IN > 245), 0),
    f_bit8_width(C_PROBE_IN244_WIDTH-1, (C_NUM_PROBE_IN > 244), 0),
    f_bit8_width(C_PROBE_IN243_WIDTH-1, (C_NUM_PROBE_IN > 243), 0),
    f_bit8_width(C_PROBE_IN242_WIDTH-1, (C_NUM_PROBE_IN > 242), 0),
    f_bit8_width(C_PROBE_IN241_WIDTH-1, (C_NUM_PROBE_IN > 241), 0),
    f_bit8_width(C_PROBE_IN240_WIDTH-1, (C_NUM_PROBE_IN > 240), 0),
    f_bit8_width(C_PROBE_IN239_WIDTH-1, (C_NUM_PROBE_IN > 239), 0),
    f_bit8_width(C_PROBE_IN238_WIDTH-1, (C_NUM_PROBE_IN > 238), 0),
    f_bit8_width(C_PROBE_IN237_WIDTH-1, (C_NUM_PROBE_IN > 237), 0),
    f_bit8_width(C_PROBE_IN236_WIDTH-1, (C_NUM_PROBE_IN > 236), 0),
    f_bit8_width(C_PROBE_IN235_WIDTH-1, (C_NUM_PROBE_IN > 235), 0),
    f_bit8_width(C_PROBE_IN234_WIDTH-1, (C_NUM_PROBE_IN > 234), 0),
    f_bit8_width(C_PROBE_IN233_WIDTH-1, (C_NUM_PROBE_IN > 233), 0),
    f_bit8_width(C_PROBE_IN232_WIDTH-1, (C_NUM_PROBE_IN > 232), 0),
    f_bit8_width(C_PROBE_IN231_WIDTH-1, (C_NUM_PROBE_IN > 231), 0),
    f_bit8_width(C_PROBE_IN230_WIDTH-1, (C_NUM_PROBE_IN > 230), 0),
    f_bit8_width(C_PROBE_IN229_WIDTH-1, (C_NUM_PROBE_IN > 229), 0),
    f_bit8_width(C_PROBE_IN228_WIDTH-1, (C_NUM_PROBE_IN > 228), 0),
    f_bit8_width(C_PROBE_IN227_WIDTH-1, (C_NUM_PROBE_IN > 227), 0),
    f_bit8_width(C_PROBE_IN226_WIDTH-1, (C_NUM_PROBE_IN > 226), 0),
    f_bit8_width(C_PROBE_IN225_WIDTH-1, (C_NUM_PROBE_IN > 225), 0),
    f_bit8_width(C_PROBE_IN224_WIDTH-1, (C_NUM_PROBE_IN > 224), 0),
    f_bit8_width(C_PROBE_IN223_WIDTH-1, (C_NUM_PROBE_IN > 223), 0),
    f_bit8_width(C_PROBE_IN222_WIDTH-1, (C_NUM_PROBE_IN > 222), 0),
    f_bit8_width(C_PROBE_IN221_WIDTH-1, (C_NUM_PROBE_IN > 221), 0),
    f_bit8_width(C_PROBE_IN220_WIDTH-1, (C_NUM_PROBE_IN > 220), 0),
    f_bit8_width(C_PROBE_IN219_WIDTH-1, (C_NUM_PROBE_IN > 219), 0),
    f_bit8_width(C_PROBE_IN218_WIDTH-1, (C_NUM_PROBE_IN > 218), 0),
    f_bit8_width(C_PROBE_IN217_WIDTH-1, (C_NUM_PROBE_IN > 217), 0),
    f_bit8_width(C_PROBE_IN216_WIDTH-1, (C_NUM_PROBE_IN > 216), 0),
    f_bit8_width(C_PROBE_IN215_WIDTH-1, (C_NUM_PROBE_IN > 215), 0),
    f_bit8_width(C_PROBE_IN214_WIDTH-1, (C_NUM_PROBE_IN > 214), 0),
    f_bit8_width(C_PROBE_IN213_WIDTH-1, (C_NUM_PROBE_IN > 213), 0),
    f_bit8_width(C_PROBE_IN212_WIDTH-1, (C_NUM_PROBE_IN > 212), 0),
    f_bit8_width(C_PROBE_IN211_WIDTH-1, (C_NUM_PROBE_IN > 211), 0),
    f_bit8_width(C_PROBE_IN210_WIDTH-1, (C_NUM_PROBE_IN > 210), 0),
    f_bit8_width(C_PROBE_IN209_WIDTH-1, (C_NUM_PROBE_IN > 209), 0),
    f_bit8_width(C_PROBE_IN208_WIDTH-1, (C_NUM_PROBE_IN > 208), 0),
    f_bit8_width(C_PROBE_IN207_WIDTH-1, (C_NUM_PROBE_IN > 207), 0),
    f_bit8_width(C_PROBE_IN206_WIDTH-1, (C_NUM_PROBE_IN > 206), 0),
    f_bit8_width(C_PROBE_IN205_WIDTH-1, (C_NUM_PROBE_IN > 205), 0),
    f_bit8_width(C_PROBE_IN204_WIDTH-1, (C_NUM_PROBE_IN > 204), 0),
    f_bit8_width(C_PROBE_IN203_WIDTH-1, (C_NUM_PROBE_IN > 203), 0),
    f_bit8_width(C_PROBE_IN202_WIDTH-1, (C_NUM_PROBE_IN > 202), 0),
    f_bit8_width(C_PROBE_IN201_WIDTH-1, (C_NUM_PROBE_IN > 201), 0),
    f_bit8_width(C_PROBE_IN200_WIDTH-1, (C_NUM_PROBE_IN > 200), 0),
    f_bit8_width(C_PROBE_IN199_WIDTH-1, (C_NUM_PROBE_IN > 199), 0),
    f_bit8_width(C_PROBE_IN198_WIDTH-1, (C_NUM_PROBE_IN > 198), 0),
    f_bit8_width(C_PROBE_IN197_WIDTH-1, (C_NUM_PROBE_IN > 197), 0),
    f_bit8_width(C_PROBE_IN196_WIDTH-1, (C_NUM_PROBE_IN > 196), 0),
    f_bit8_width(C_PROBE_IN195_WIDTH-1, (C_NUM_PROBE_IN > 195), 0),
    f_bit8_width(C_PROBE_IN194_WIDTH-1, (C_NUM_PROBE_IN > 194), 0),
    f_bit8_width(C_PROBE_IN193_WIDTH-1, (C_NUM_PROBE_IN > 193), 0),
    f_bit8_width(C_PROBE_IN192_WIDTH-1, (C_NUM_PROBE_IN > 192), 0),
    f_bit8_width(C_PROBE_IN191_WIDTH-1, (C_NUM_PROBE_IN > 191), 0),
    f_bit8_width(C_PROBE_IN190_WIDTH-1, (C_NUM_PROBE_IN > 190), 0),
        f_bit8_width(C_PROBE_IN161_WIDTH-1, (C_NUM_PROBE_IN > 161), 0),
    f_bit8_width(C_PROBE_IN160_WIDTH-1, (C_NUM_PROBE_IN > 160), 0),
    f_bit8_width(C_PROBE_IN159_WIDTH-1, (C_NUM_PROBE_IN > 159), 0),
    f_bit8_width(C_PROBE_IN158_WIDTH-1, (C_NUM_PROBE_IN > 158), 0),
    f_bit8_width(C_PROBE_IN157_WIDTH-1, (C_NUM_PROBE_IN > 157), 0),
    f_bit8_width(C_PROBE_IN156_WIDTH-1, (C_NUM_PROBE_IN > 156), 0),
    f_bit8_width(C_PROBE_IN155_WIDTH-1, (C_NUM_PROBE_IN > 155), 0),
    f_bit8_width(C_PROBE_IN154_WIDTH-1, (C_NUM_PROBE_IN > 154), 0),
    f_bit8_width(C_PROBE_IN153_WIDTH-1, (C_NUM_PROBE_IN > 153), 0),
    f_bit8_width(C_PROBE_IN152_WIDTH-1, (C_NUM_PROBE_IN > 152), 0),
    f_bit8_width(C_PROBE_IN151_WIDTH-1, (C_NUM_PROBE_IN > 151), 0),
    f_bit8_width(C_PROBE_IN150_WIDTH-1, (C_NUM_PROBE_IN > 150), 0),
    f_bit8_width(C_PROBE_IN149_WIDTH-1, (C_NUM_PROBE_IN > 149), 0),
    f_bit8_width(C_PROBE_IN148_WIDTH-1, (C_NUM_PROBE_IN > 148), 0),
    f_bit8_width(C_PROBE_IN147_WIDTH-1, (C_NUM_PROBE_IN > 147), 0),
    f_bit8_width(C_PROBE_IN146_WIDTH-1, (C_NUM_PROBE_IN > 146), 0),
    f_bit8_width(C_PROBE_IN145_WIDTH-1, (C_NUM_PROBE_IN > 145), 0),
    f_bit8_width(C_PROBE_IN144_WIDTH-1, (C_NUM_PROBE_IN > 144), 0),
    f_bit8_width(C_PROBE_IN143_WIDTH-1, (C_NUM_PROBE_IN > 143), 0),
    f_bit8_width(C_PROBE_IN142_WIDTH-1, (C_NUM_PROBE_IN > 142), 0),
    f_bit8_width(C_PROBE_IN141_WIDTH-1, (C_NUM_PROBE_IN > 141), 0),
    f_bit8_width(C_PROBE_IN140_WIDTH-1, (C_NUM_PROBE_IN > 140), 0),
    f_bit8_width(C_PROBE_IN139_WIDTH-1, (C_NUM_PROBE_IN > 139), 0),
    f_bit8_width(C_PROBE_IN138_WIDTH-1, (C_NUM_PROBE_IN > 138), 0),
    f_bit8_width(C_PROBE_IN137_WIDTH-1, (C_NUM_PROBE_IN > 137), 0),
    f_bit8_width(C_PROBE_IN136_WIDTH-1, (C_NUM_PROBE_IN > 136), 0),
    f_bit8_width(C_PROBE_IN135_WIDTH-1, (C_NUM_PROBE_IN > 135), 0),
    f_bit8_width(C_PROBE_IN134_WIDTH-1, (C_NUM_PROBE_IN > 134), 0),
    f_bit8_width(C_PROBE_IN133_WIDTH-1, (C_NUM_PROBE_IN > 133), 0),
    f_bit8_width(C_PROBE_IN132_WIDTH-1, (C_NUM_PROBE_IN > 132), 0),
    f_bit8_width(C_PROBE_IN131_WIDTH-1, (C_NUM_PROBE_IN > 131), 0),
    f_bit8_width(C_PROBE_IN130_WIDTH-1, (C_NUM_PROBE_IN > 130), 0),
    f_bit8_width(C_PROBE_IN129_WIDTH-1, (C_NUM_PROBE_IN > 129), 0),
    f_bit8_width(C_PROBE_IN128_WIDTH-1, (C_NUM_PROBE_IN > 128), 0),
    f_bit8_width(C_PROBE_IN127_WIDTH-1, (C_NUM_PROBE_IN > 127), 0),
    f_bit8_width(C_PROBE_IN126_WIDTH-1, (C_NUM_PROBE_IN > 126), 0),
    f_bit8_width(C_PROBE_IN125_WIDTH-1, (C_NUM_PROBE_IN > 125), 0),
    f_bit8_width(C_PROBE_IN124_WIDTH-1, (C_NUM_PROBE_IN > 124), 0),
    f_bit8_width(C_PROBE_IN123_WIDTH-1, (C_NUM_PROBE_IN > 123), 0),
    f_bit8_width(C_PROBE_IN122_WIDTH-1, (C_NUM_PROBE_IN > 122), 0),
    f_bit8_width(C_PROBE_IN121_WIDTH-1, (C_NUM_PROBE_IN > 121), 0),
    f_bit8_width(C_PROBE_IN120_WIDTH-1, (C_NUM_PROBE_IN > 120), 0),
    f_bit8_width(C_PROBE_IN119_WIDTH-1, (C_NUM_PROBE_IN > 119), 0),
    f_bit8_width(C_PROBE_IN118_WIDTH-1, (C_NUM_PROBE_IN > 118), 0),
    f_bit8_width(C_PROBE_IN117_WIDTH-1, (C_NUM_PROBE_IN > 117), 0),
    f_bit8_width(C_PROBE_IN116_WIDTH-1, (C_NUM_PROBE_IN > 116), 0),
    f_bit8_width(C_PROBE_IN115_WIDTH-1, (C_NUM_PROBE_IN > 115), 0),
    f_bit8_width(C_PROBE_IN114_WIDTH-1, (C_NUM_PROBE_IN > 114), 0),
    f_bit8_width(C_PROBE_IN113_WIDTH-1, (C_NUM_PROBE_IN > 113), 0),
    f_bit8_width(C_PROBE_IN112_WIDTH-1, (C_NUM_PROBE_IN > 112), 0),
    f_bit8_width(C_PROBE_IN111_WIDTH-1, (C_NUM_PROBE_IN > 111), 0),
    f_bit8_width(C_PROBE_IN110_WIDTH-1, (C_NUM_PROBE_IN > 110), 0),
    f_bit8_width(C_PROBE_IN109_WIDTH-1, (C_NUM_PROBE_IN > 109), 0),
    f_bit8_width(C_PROBE_IN108_WIDTH-1, (C_NUM_PROBE_IN > 108), 0),
    f_bit8_width(C_PROBE_IN107_WIDTH-1, (C_NUM_PROBE_IN > 107), 0),
    f_bit8_width(C_PROBE_IN106_WIDTH-1, (C_NUM_PROBE_IN > 106), 0),
    f_bit8_width(C_PROBE_IN105_WIDTH-1, (C_NUM_PROBE_IN > 105), 0),
    f_bit8_width(C_PROBE_IN104_WIDTH-1, (C_NUM_PROBE_IN > 104), 0),
    f_bit8_width(C_PROBE_IN103_WIDTH-1, (C_NUM_PROBE_IN > 103), 0),
    f_bit8_width(C_PROBE_IN102_WIDTH-1, (C_NUM_PROBE_IN > 102), 0),
    f_bit8_width(C_PROBE_IN101_WIDTH-1, (C_NUM_PROBE_IN > 101), 0),
    f_bit8_width(C_PROBE_IN100_WIDTH-1, (C_NUM_PROBE_IN > 100), 0),
    f_bit8_width(C_PROBE_IN99_WIDTH-1 , (C_NUM_PROBE_IN > 99), 0),
    f_bit8_width(C_PROBE_IN98_WIDTH-1 , (C_NUM_PROBE_IN > 98), 0),
    f_bit8_width(C_PROBE_IN97_WIDTH-1 , (C_NUM_PROBE_IN > 97), 0),
    f_bit8_width(C_PROBE_IN96_WIDTH-1 , (C_NUM_PROBE_IN > 96), 0),
    f_bit8_width(C_PROBE_IN95_WIDTH-1 , (C_NUM_PROBE_IN > 95), 0),
    f_bit8_width(C_PROBE_IN94_WIDTH-1 , (C_NUM_PROBE_IN > 94), 0),
    f_bit8_width(C_PROBE_IN93_WIDTH-1 , (C_NUM_PROBE_IN > 93), 0),
    f_bit8_width(C_PROBE_IN92_WIDTH-1 , (C_NUM_PROBE_IN > 92), 0),
    f_bit8_width(C_PROBE_IN91_WIDTH-1 , (C_NUM_PROBE_IN > 91), 0),
    f_bit8_width(C_PROBE_IN90_WIDTH-1 , (C_NUM_PROBE_IN > 90), 0),
    f_bit8_width(C_PROBE_IN89_WIDTH-1 , (C_NUM_PROBE_IN > 89), 0),
    f_bit8_width(C_PROBE_IN88_WIDTH-1 , (C_NUM_PROBE_IN > 88), 0),
    f_bit8_width(C_PROBE_IN87_WIDTH-1 , (C_NUM_PROBE_IN > 87), 0),
    f_bit8_width(C_PROBE_IN86_WIDTH-1 , (C_NUM_PROBE_IN > 86), 0),
    f_bit8_width(C_PROBE_IN85_WIDTH-1 , (C_NUM_PROBE_IN > 85), 0),
    f_bit8_width(C_PROBE_IN84_WIDTH-1 , (C_NUM_PROBE_IN > 84), 0),
    f_bit8_width(C_PROBE_IN83_WIDTH-1 , (C_NUM_PROBE_IN > 83), 0),
    f_bit8_width(C_PROBE_IN82_WIDTH-1 , (C_NUM_PROBE_IN > 82), 0),
    f_bit8_width(C_PROBE_IN81_WIDTH-1 , (C_NUM_PROBE_IN > 81), 0),
    f_bit8_width(C_PROBE_IN80_WIDTH-1 , (C_NUM_PROBE_IN > 80), 0),
    f_bit8_width(C_PROBE_IN79_WIDTH-1 , (C_NUM_PROBE_IN > 79), 0),
    f_bit8_width(C_PROBE_IN78_WIDTH-1 , (C_NUM_PROBE_IN > 78), 0),
    f_bit8_width(C_PROBE_IN77_WIDTH-1 , (C_NUM_PROBE_IN > 77), 0),
    f_bit8_width(C_PROBE_IN76_WIDTH-1 , (C_NUM_PROBE_IN > 76), 0),
    f_bit8_width(C_PROBE_IN75_WIDTH-1 , (C_NUM_PROBE_IN > 75), 0),
    f_bit8_width(C_PROBE_IN74_WIDTH-1 , (C_NUM_PROBE_IN > 74), 0),
    f_bit8_width(C_PROBE_IN73_WIDTH-1 , (C_NUM_PROBE_IN > 73), 0),
    f_bit8_width(C_PROBE_IN72_WIDTH-1 , (C_NUM_PROBE_IN > 72), 0),
    f_bit8_width(C_PROBE_IN71_WIDTH-1 , (C_NUM_PROBE_IN > 71), 0),
    f_bit8_width(C_PROBE_IN70_WIDTH-1 , (C_NUM_PROBE_IN > 70), 0),
    f_bit8_width(C_PROBE_IN69_WIDTH-1 , (C_NUM_PROBE_IN > 69), 0),
    f_bit8_width(C_PROBE_IN68_WIDTH-1 , (C_NUM_PROBE_IN > 68), 0),
    f_bit8_width(C_PROBE_IN67_WIDTH-1 , (C_NUM_PROBE_IN > 67), 0),
    f_bit8_width(C_PROBE_IN66_WIDTH-1 , (C_NUM_PROBE_IN > 66), 0),
    f_bit8_width(C_PROBE_IN65_WIDTH-1 , (C_NUM_PROBE_IN > 65), 0),
    f_bit8_width(C_PROBE_IN64_WIDTH-1 , (C_NUM_PROBE_IN > 64), 0),
    f_bit8_width(C_PROBE_IN63_WIDTH-1 , (C_NUM_PROBE_IN > 63), 0),
    f_bit8_width(C_PROBE_IN62_WIDTH-1 , (C_NUM_PROBE_IN > 62), 0),
    f_bit8_width(C_PROBE_IN61_WIDTH-1 , (C_NUM_PROBE_IN > 61), 0),
    f_bit8_width(C_PROBE_IN60_WIDTH-1 , (C_NUM_PROBE_IN > 60), 0),
    f_bit8_width(C_PROBE_IN59_WIDTH-1 , (C_NUM_PROBE_IN > 59), 0),
    f_bit8_width(C_PROBE_IN58_WIDTH-1 , (C_NUM_PROBE_IN > 58), 0),
    f_bit8_width(C_PROBE_IN57_WIDTH-1 , (C_NUM_PROBE_IN > 57), 0),
    f_bit8_width(C_PROBE_IN56_WIDTH-1 , (C_NUM_PROBE_IN > 56), 0),
    f_bit8_width(C_PROBE_IN55_WIDTH-1 , (C_NUM_PROBE_IN > 55), 0),
    f_bit8_width(C_PROBE_IN54_WIDTH-1 , (C_NUM_PROBE_IN > 54), 0),
    f_bit8_width(C_PROBE_IN53_WIDTH-1 , (C_NUM_PROBE_IN > 53), 0),
    f_bit8_width(C_PROBE_IN52_WIDTH-1 , (C_NUM_PROBE_IN > 52), 0),
    f_bit8_width(C_PROBE_IN51_WIDTH-1 , (C_NUM_PROBE_IN > 51), 0),
    f_bit8_width(C_PROBE_IN50_WIDTH-1 , (C_NUM_PROBE_IN > 50), 0),
    f_bit8_width(C_PROBE_IN49_WIDTH-1 , (C_NUM_PROBE_IN > 49), 0),
    f_bit8_width(C_PROBE_IN48_WIDTH-1 , (C_NUM_PROBE_IN > 48), 0),
    f_bit8_width(C_PROBE_IN47_WIDTH-1 , (C_NUM_PROBE_IN > 47), 0),
    f_bit8_width(C_PROBE_IN46_WIDTH-1 , (C_NUM_PROBE_IN > 46), 0),
    f_bit8_width(C_PROBE_IN45_WIDTH-1 , (C_NUM_PROBE_IN > 45), 0),
    f_bit8_width(C_PROBE_IN44_WIDTH-1 , (C_NUM_PROBE_IN > 44), 0),
    f_bit8_width(C_PROBE_IN43_WIDTH-1 , (C_NUM_PROBE_IN > 43), 0),
    f_bit8_width(C_PROBE_IN42_WIDTH-1 , (C_NUM_PROBE_IN > 42), 0),
    f_bit8_width(C_PROBE_IN41_WIDTH-1 , (C_NUM_PROBE_IN > 41), 0),
    f_bit8_width(C_PROBE_IN40_WIDTH-1 , (C_NUM_PROBE_IN > 40), 0),
    f_bit8_width(C_PROBE_IN39_WIDTH-1 , (C_NUM_PROBE_IN > 39), 0),
    f_bit8_width(C_PROBE_IN38_WIDTH-1 , (C_NUM_PROBE_IN > 38), 0),
    f_bit8_width(C_PROBE_IN37_WIDTH-1 , (C_NUM_PROBE_IN > 37), 0),
    f_bit8_width(C_PROBE_IN36_WIDTH-1 , (C_NUM_PROBE_IN > 36), 0),
    f_bit8_width(C_PROBE_IN35_WIDTH-1 , (C_NUM_PROBE_IN > 35), 0),
    f_bit8_width(C_PROBE_IN34_WIDTH-1 , (C_NUM_PROBE_IN > 34), 0),
    f_bit8_width(C_PROBE_IN33_WIDTH-1 , (C_NUM_PROBE_IN > 33), 0),
    f_bit8_width(C_PROBE_IN32_WIDTH-1 , (C_NUM_PROBE_IN > 32), 0),
    f_bit8_width(C_PROBE_IN31_WIDTH-1 , (C_NUM_PROBE_IN > 31), 0),
    f_bit8_width(C_PROBE_IN30_WIDTH-1 , (C_NUM_PROBE_IN > 30), 0),
    f_bit8_width(C_PROBE_IN29_WIDTH-1 , (C_NUM_PROBE_IN > 29), 0),
    f_bit8_width(C_PROBE_IN28_WIDTH-1 , (C_NUM_PROBE_IN > 28), 0),
    f_bit8_width(C_PROBE_IN27_WIDTH-1 , (C_NUM_PROBE_IN > 27), 0),
    f_bit8_width(C_PROBE_IN26_WIDTH-1 , (C_NUM_PROBE_IN > 26), 0),
    f_bit8_width(C_PROBE_IN25_WIDTH-1 , (C_NUM_PROBE_IN > 25), 0),
    f_bit8_width(C_PROBE_IN24_WIDTH-1 , (C_NUM_PROBE_IN > 24), 0),
    f_bit8_width(C_PROBE_IN23_WIDTH-1 , (C_NUM_PROBE_IN > 23), 0),
    f_bit8_width(C_PROBE_IN22_WIDTH-1 , (C_NUM_PROBE_IN > 22), 0),
    f_bit8_width(C_PROBE_IN21_WIDTH-1 , (C_NUM_PROBE_IN > 21), 0),
    f_bit8_width(C_PROBE_IN20_WIDTH-1 , (C_NUM_PROBE_IN > 20), 0),
    f_bit8_width(C_PROBE_IN19_WIDTH-1 , (C_NUM_PROBE_IN > 19), 0),
    f_bit8_width(C_PROBE_IN18_WIDTH-1 , (C_NUM_PROBE_IN > 18), 0),
    f_bit8_width(C_PROBE_IN17_WIDTH-1 , (C_NUM_PROBE_IN > 17), 0),
    f_bit8_width(C_PROBE_IN16_WIDTH-1 , (C_NUM_PROBE_IN > 16), 0),
    f_bit8_width(C_PROBE_IN15_WIDTH-1 , (C_NUM_PROBE_IN > 15), 0),
    f_bit8_width(C_PROBE_IN14_WIDTH-1 , (C_NUM_PROBE_IN > 14), 0),
    f_bit8_width(C_PROBE_IN13_WIDTH-1 , (C_NUM_PROBE_IN > 13), 0),
    f_bit8_width(C_PROBE_IN12_WIDTH-1 , (C_NUM_PROBE_IN > 12), 0),
    f_bit8_width(C_PROBE_IN11_WIDTH-1 , (C_NUM_PROBE_IN > 11), 0),
    f_bit8_width(C_PROBE_IN10_WIDTH-1 , (C_NUM_PROBE_IN > 10), 0),
    f_bit8_width(C_PROBE_IN9_WIDTH-1  , (C_NUM_PROBE_IN >  9), 0),
    f_bit8_width(C_PROBE_IN8_WIDTH-1  , (C_NUM_PROBE_IN >  8), 0),
    f_bit8_width(C_PROBE_IN7_WIDTH-1  , (C_NUM_PROBE_IN >  7), 0),
    f_bit8_width(C_PROBE_IN6_WIDTH-1  , (C_NUM_PROBE_IN >  6), 0),
    f_bit8_width(C_PROBE_IN5_WIDTH-1  , (C_NUM_PROBE_IN >  5), 0),
    f_bit8_width(C_PROBE_IN4_WIDTH-1  , (C_NUM_PROBE_IN >  4), 0),
    f_bit8_width(C_PROBE_IN3_WIDTH-1  , (C_NUM_PROBE_IN >  3), 0),
    f_bit8_width(C_PROBE_IN2_WIDTH-1  , (C_NUM_PROBE_IN >  2), 0),
    f_bit8_width(C_PROBE_IN1_WIDTH-1  , (C_NUM_PROBE_IN >  1), 0),
    f_bit8_width(C_PROBE_IN0_WIDTH-1  , (C_NUM_PROBE_IN >  0), 0)
  };

  localparam LC_TOTAL_PROBE_OUT_WIDTH  = (
        C_PROBE_OUT255_WIDTH + C_PROBE_OUT254_WIDTH + C_PROBE_OUT253_WIDTH +
        C_PROBE_OUT252_WIDTH + C_PROBE_OUT251_WIDTH + C_PROBE_OUT250_WIDTH +
        C_PROBE_OUT249_WIDTH + C_PROBE_OUT248_WIDTH + C_PROBE_OUT247_WIDTH +
        C_PROBE_OUT246_WIDTH + C_PROBE_OUT245_WIDTH + C_PROBE_OUT244_WIDTH + 
        C_PROBE_OUT243_WIDTH + C_PROBE_OUT242_WIDTH + C_PROBE_OUT241_WIDTH +
        C_PROBE_OUT240_WIDTH + C_PROBE_OUT239_WIDTH + C_PROBE_OUT238_WIDTH +
        C_PROBE_OUT237_WIDTH + C_PROBE_OUT236_WIDTH + C_PROBE_OUT235_WIDTH +
        C_PROBE_OUT234_WIDTH + C_PROBE_OUT233_WIDTH + C_PROBE_OUT232_WIDTH +
        C_PROBE_OUT231_WIDTH + C_PROBE_OUT230_WIDTH + C_PROBE_OUT229_WIDTH +
        C_PROBE_OUT228_WIDTH + C_PROBE_OUT227_WIDTH + C_PROBE_OUT226_WIDTH +
        C_PROBE_OUT225_WIDTH + C_PROBE_OUT224_WIDTH + C_PROBE_OUT223_WIDTH + 
        C_PROBE_OUT222_WIDTH + C_PROBE_OUT221_WIDTH + C_PROBE_OUT220_WIDTH +
        C_PROBE_OUT219_WIDTH + C_PROBE_OUT218_WIDTH + C_PROBE_OUT217_WIDTH +
        C_PROBE_OUT216_WIDTH + C_PROBE_OUT215_WIDTH + C_PROBE_OUT214_WIDTH +
        C_PROBE_OUT213_WIDTH + C_PROBE_OUT212_WIDTH + C_PROBE_OUT211_WIDTH +
        C_PROBE_OUT210_WIDTH + C_PROBE_OUT209_WIDTH + C_PROBE_OUT208_WIDTH +
        C_PROBE_OUT207_WIDTH + C_PROBE_OUT206_WIDTH + C_PROBE_OUT205_WIDTH +
        C_PROBE_OUT204_WIDTH + C_PROBE_OUT203_WIDTH + C_PROBE_OUT202_WIDTH +
        C_PROBE_OUT201_WIDTH + C_PROBE_OUT200_WIDTH + C_PROBE_OUT199_WIDTH +
        C_PROBE_OUT198_WIDTH + C_PROBE_OUT197_WIDTH + C_PROBE_OUT196_WIDTH +
        C_PROBE_OUT195_WIDTH + C_PROBE_OUT194_WIDTH + C_PROBE_OUT193_WIDTH +
        C_PROBE_OUT192_WIDTH + C_PROBE_OUT191_WIDTH + C_PROBE_OUT190_WIDTH +
        C_PROBE_OUT189_WIDTH + C_PROBE_OUT188_WIDTH + C_PROBE_OUT187_WIDTH +
        C_PROBE_OUT186_WIDTH + C_PROBE_OUT185_WIDTH + C_PROBE_OUT184_WIDTH +
        C_PROBE_OUT183_WIDTH + C_PROBE_OUT182_WIDTH + C_PROBE_OUT181_WIDTH +
        C_PROBE_OUT180_WIDTH + C_PROBE_OUT179_WIDTH + C_PROBE_OUT178_WIDTH +
        C_PROBE_OUT177_WIDTH + C_PROBE_OUT176_WIDTH + C_PROBE_OUT175_WIDTH +
        C_PROBE_OUT174_WIDTH + C_PROBE_OUT173_WIDTH + C_PROBE_OUT172_WIDTH +
        C_PROBE_OUT171_WIDTH + C_PROBE_OUT170_WIDTH + C_PROBE_OUT169_WIDTH +
        C_PROBE_OUT168_WIDTH + C_PROBE_OUT167_WIDTH + C_PROBE_OUT166_WIDTH +
        C_PROBE_OUT165_WIDTH + C_PROBE_OUT164_WIDTH + C_PROBE_OUT163_WIDTH +
        C_PROBE_OUT162_WIDTH + C_PROBE_OUT161_WIDTH + C_PROBE_OUT160_WIDTH +
        C_PROBE_OUT159_WIDTH + C_PROBE_OUT158_WIDTH + C_PROBE_OUT157_WIDTH +
        C_PROBE_OUT156_WIDTH + C_PROBE_OUT155_WIDTH + C_PROBE_OUT154_WIDTH +
        C_PROBE_OUT153_WIDTH + C_PROBE_OUT152_WIDTH + C_PROBE_OUT151_WIDTH +
        C_PROBE_OUT150_WIDTH + C_PROBE_OUT149_WIDTH + C_PROBE_OUT148_WIDTH +
        C_PROBE_OUT147_WIDTH + C_PROBE_OUT146_WIDTH + C_PROBE_OUT145_WIDTH + 
        C_PROBE_OUT144_WIDTH + C_PROBE_OUT143_WIDTH + C_PROBE_OUT142_WIDTH +
        C_PROBE_OUT141_WIDTH + C_PROBE_OUT140_WIDTH + C_PROBE_OUT139_WIDTH +
        C_PROBE_OUT138_WIDTH + C_PROBE_OUT137_WIDTH + C_PROBE_OUT136_WIDTH +
        C_PROBE_OUT135_WIDTH + C_PROBE_OUT134_WIDTH + C_PROBE_OUT133_WIDTH +
        C_PROBE_OUT132_WIDTH + C_PROBE_OUT131_WIDTH + C_PROBE_OUT130_WIDTH +
        C_PROBE_OUT129_WIDTH + C_PROBE_OUT128_WIDTH + C_PROBE_OUT127_WIDTH +
        C_PROBE_OUT126_WIDTH + C_PROBE_OUT125_WIDTH + C_PROBE_OUT124_WIDTH +
        C_PROBE_OUT123_WIDTH + C_PROBE_OUT122_WIDTH + C_PROBE_OUT121_WIDTH + 
        C_PROBE_OUT120_WIDTH + C_PROBE_OUT119_WIDTH + C_PROBE_OUT118_WIDTH +
        C_PROBE_OUT117_WIDTH + C_PROBE_OUT116_WIDTH + C_PROBE_OUT115_WIDTH +
        C_PROBE_OUT114_WIDTH + C_PROBE_OUT113_WIDTH + C_PROBE_OUT112_WIDTH +
        C_PROBE_OUT111_WIDTH + C_PROBE_OUT110_WIDTH + C_PROBE_OUT109_WIDTH +
        C_PROBE_OUT108_WIDTH + C_PROBE_OUT107_WIDTH + C_PROBE_OUT106_WIDTH +
        C_PROBE_OUT105_WIDTH + C_PROBE_OUT104_WIDTH + C_PROBE_OUT103_WIDTH +
        C_PROBE_OUT102_WIDTH + C_PROBE_OUT101_WIDTH + C_PROBE_OUT100_WIDTH +
        C_PROBE_OUT99_WIDTH  + C_PROBE_OUT98_WIDTH  + C_PROBE_OUT97_WIDTH  +
        C_PROBE_OUT96_WIDTH  + C_PROBE_OUT95_WIDTH  + C_PROBE_OUT94_WIDTH  +
        C_PROBE_OUT93_WIDTH  + C_PROBE_OUT92_WIDTH  + C_PROBE_OUT91_WIDTH  +
        C_PROBE_OUT90_WIDTH  + C_PROBE_OUT89_WIDTH  + C_PROBE_OUT88_WIDTH  +
        C_PROBE_OUT87_WIDTH  + C_PROBE_OUT86_WIDTH  + C_PROBE_OUT85_WIDTH  +
        C_PROBE_OUT84_WIDTH  + C_PROBE_OUT83_WIDTH  + C_PROBE_OUT82_WIDTH  +
        C_PROBE_OUT81_WIDTH  + C_PROBE_OUT80_WIDTH  + C_PROBE_OUT79_WIDTH  +
        C_PROBE_OUT78_WIDTH  + C_PROBE_OUT77_WIDTH  + C_PROBE_OUT76_WIDTH  +
        C_PROBE_OUT75_WIDTH  + C_PROBE_OUT74_WIDTH  + C_PROBE_OUT73_WIDTH  +
        C_PROBE_OUT72_WIDTH  + C_PROBE_OUT71_WIDTH  + C_PROBE_OUT70_WIDTH  +
        C_PROBE_OUT69_WIDTH  + C_PROBE_OUT68_WIDTH  + C_PROBE_OUT67_WIDTH  +
        C_PROBE_OUT66_WIDTH  + C_PROBE_OUT65_WIDTH  + C_PROBE_OUT64_WIDTH  +
        C_PROBE_OUT63_WIDTH  + C_PROBE_OUT62_WIDTH  + C_PROBE_OUT61_WIDTH  +
        C_PROBE_OUT60_WIDTH  + C_PROBE_OUT59_WIDTH  + C_PROBE_OUT58_WIDTH  +
        C_PROBE_OUT57_WIDTH  + C_PROBE_OUT56_WIDTH  + C_PROBE_OUT55_WIDTH  +
        C_PROBE_OUT54_WIDTH  + C_PROBE_OUT53_WIDTH  + C_PROBE_OUT52_WIDTH  +
        C_PROBE_OUT51_WIDTH  + C_PROBE_OUT50_WIDTH  + C_PROBE_OUT49_WIDTH  +
        C_PROBE_OUT48_WIDTH  + C_PROBE_OUT47_WIDTH  + C_PROBE_OUT46_WIDTH  +
        C_PROBE_OUT45_WIDTH  + C_PROBE_OUT44_WIDTH  + C_PROBE_OUT43_WIDTH  +
        C_PROBE_OUT42_WIDTH  + C_PROBE_OUT41_WIDTH  + C_PROBE_OUT40_WIDTH  +
        C_PROBE_OUT39_WIDTH  + C_PROBE_OUT38_WIDTH  + C_PROBE_OUT37_WIDTH  +
        C_PROBE_OUT36_WIDTH  + C_PROBE_OUT35_WIDTH  + C_PROBE_OUT34_WIDTH  +
        C_PROBE_OUT33_WIDTH  + C_PROBE_OUT32_WIDTH  + C_PROBE_OUT31_WIDTH  +
        C_PROBE_OUT30_WIDTH  + C_PROBE_OUT29_WIDTH  + C_PROBE_OUT28_WIDTH  +
        C_PROBE_OUT27_WIDTH  + C_PROBE_OUT26_WIDTH  + C_PROBE_OUT25_WIDTH  +
        C_PROBE_OUT24_WIDTH  + C_PROBE_OUT23_WIDTH  + C_PROBE_OUT22_WIDTH  +
        C_PROBE_OUT21_WIDTH  + C_PROBE_OUT20_WIDTH  + C_PROBE_OUT19_WIDTH  +
        C_PROBE_OUT18_WIDTH  + C_PROBE_OUT17_WIDTH  + C_PROBE_OUT16_WIDTH  +
        C_PROBE_OUT15_WIDTH  + C_PROBE_OUT14_WIDTH  + C_PROBE_OUT13_WIDTH  +
        C_PROBE_OUT12_WIDTH  + C_PROBE_OUT11_WIDTH  + C_PROBE_OUT10_WIDTH  +
        C_PROBE_OUT9_WIDTH   + C_PROBE_OUT8_WIDTH   + C_PROBE_OUT7_WIDTH   +
        C_PROBE_OUT6_WIDTH   + C_PROBE_OUT5_WIDTH   + C_PROBE_OUT4_WIDTH   +
        C_PROBE_OUT3_WIDTH   + C_PROBE_OUT2_WIDTH   + C_PROBE_OUT1_WIDTH   +
        C_PROBE_OUT0_WIDTH   - C_MAX_NUM_PROBE      + C_NUM_PROBE_OUT
      );

  localparam [2047:0]LC_PROBE_OUT_WIDTH_STRING = {
    f_bit8_width(C_PROBE_OUT255_WIDTH-1, (C_NUM_PROBE_OUT > 255), 0),
    f_bit8_width(C_PROBE_OUT254_WIDTH-1, (C_NUM_PROBE_OUT > 254), 0),
    f_bit8_width(C_PROBE_OUT253_WIDTH-1, (C_NUM_PROBE_OUT > 253), 0),
    f_bit8_width(C_PROBE_OUT252_WIDTH-1, (C_NUM_PROBE_OUT > 252), 0),
    f_bit8_width(C_PROBE_OUT251_WIDTH-1, (C_NUM_PROBE_OUT > 251), 0),
    f_bit8_width(C_PROBE_OUT250_WIDTH-1, (C_NUM_PROBE_OUT > 250), 0),
    f_bit8_width(C_PROBE_OUT249_WIDTH-1, (C_NUM_PROBE_OUT > 249), 0),
    f_bit8_width(C_PROBE_OUT248_WIDTH-1, (C_NUM_PROBE_OUT > 248), 0),
    f_bit8_width(C_PROBE_OUT247_WIDTH-1, (C_NUM_PROBE_OUT > 247), 0),
    f_bit8_width(C_PROBE_OUT246_WIDTH-1, (C_NUM_PROBE_OUT > 246), 0),
    f_bit8_width(C_PROBE_OUT245_WIDTH-1, (C_NUM_PROBE_OUT > 245), 0),
    f_bit8_width(C_PROBE_OUT244_WIDTH-1, (C_NUM_PROBE_OUT > 244), 0),
    f_bit8_width(C_PROBE_OUT243_WIDTH-1, (C_NUM_PROBE_OUT > 243), 0),
    f_bit8_width(C_PROBE_OUT242_WIDTH-1, (C_NUM_PROBE_OUT > 242), 0),
    f_bit8_width(C_PROBE_OUT241_WIDTH-1, (C_NUM_PROBE_OUT > 241), 0),
    f_bit8_width(C_PROBE_OUT240_WIDTH-1, (C_NUM_PROBE_OUT > 240), 0),
    f_bit8_width(C_PROBE_OUT239_WIDTH-1, (C_NUM_PROBE_OUT > 239), 0),
    f_bit8_width(C_PROBE_OUT238_WIDTH-1, (C_NUM_PROBE_OUT > 238), 0),
    f_bit8_width(C_PROBE_OUT237_WIDTH-1, (C_NUM_PROBE_OUT > 237), 0),
    f_bit8_width(C_PROBE_OUT236_WIDTH-1, (C_NUM_PROBE_OUT > 236), 0),
    f_bit8_width(C_PROBE_OUT235_WIDTH-1, (C_NUM_PROBE_OUT > 235), 0),
    f_bit8_width(C_PROBE_OUT234_WIDTH-1, (C_NUM_PROBE_OUT > 234), 0),
    f_bit8_width(C_PROBE_OUT233_WIDTH-1, (C_NUM_PROBE_OUT > 233), 0),
    f_bit8_width(C_PROBE_OUT232_WIDTH-1, (C_NUM_PROBE_OUT > 232), 0),
    f_bit8_width(C_PROBE_OUT231_WIDTH-1, (C_NUM_PROBE_OUT > 231), 0),
    f_bit8_width(C_PROBE_OUT230_WIDTH-1, (C_NUM_PROBE_OUT > 230), 0),
    f_bit8_width(C_PROBE_OUT229_WIDTH-1, (C_NUM_PROBE_OUT > 229), 0),
    f_bit8_width(C_PROBE_OUT228_WIDTH-1, (C_NUM_PROBE_OUT > 228), 0),
    f_bit8_width(C_PROBE_OUT227_WIDTH-1, (C_NUM_PROBE_OUT > 227), 0),
    f_bit8_width(C_PROBE_OUT226_WIDTH-1, (C_NUM_PROBE_OUT > 226), 0),
    f_bit8_width(C_PROBE_OUT225_WIDTH-1, (C_NUM_PROBE_OUT > 225), 0),
    f_bit8_width(C_PROBE_OUT224_WIDTH-1, (C_NUM_PROBE_OUT > 224), 0),
    f_bit8_width(C_PROBE_OUT223_WIDTH-1, (C_NUM_PROBE_OUT > 223), 0),
    f_bit8_width(C_PROBE_OUT222_WIDTH-1, (C_NUM_PROBE_OUT > 222), 0),
    f_bit8_width(C_PROBE_OUT221_WIDTH-1, (C_NUM_PROBE_OUT > 221), 0),
    f_bit8_width(C_PROBE_OUT220_WIDTH-1, (C_NUM_PROBE_OUT > 220), 0),
    f_bit8_width(C_PROBE_OUT219_WIDTH-1, (C_NUM_PROBE_OUT > 219), 0),
    f_bit8_width(C_PROBE_OUT218_WIDTH-1, (C_NUM_PROBE_OUT > 218), 0),
    f_bit8_width(C_PROBE_OUT217_WIDTH-1, (C_NUM_PROBE_OUT > 217), 0),
    f_bit8_width(C_PROBE_OUT216_WIDTH-1, (C_NUM_PROBE_OUT > 216), 0),
    f_bit8_width(C_PROBE_OUT215_WIDTH-1, (C_NUM_PROBE_OUT > 215), 0),
    f_bit8_width(C_PROBE_OUT214_WIDTH-1, (C_NUM_PROBE_OUT > 214), 0),
    f_bit8_width(C_PROBE_OUT213_WIDTH-1, (C_NUM_PROBE_OUT > 213), 0),
    f_bit8_width(C_PROBE_OUT212_WIDTH-1, (C_NUM_PROBE_OUT > 212), 0),
    f_bit8_width(C_PROBE_OUT211_WIDTH-1, (C_NUM_PROBE_OUT > 211), 0),
    f_bit8_width(C_PROBE_OUT210_WIDTH-1, (C_NUM_PROBE_OUT > 210), 0),
    f_bit8_width(C_PROBE_OUT209_WIDTH-1, (C_NUM_PROBE_OUT > 209), 0),
    f_bit8_width(C_PROBE_OUT208_WIDTH-1, (C_NUM_PROBE_OUT > 208), 0),
    f_bit8_width(C_PROBE_OUT207_WIDTH-1, (C_NUM_PROBE_OUT > 207), 0),
    f_bit8_width(C_PROBE_OUT206_WIDTH-1, (C_NUM_PROBE_OUT > 206), 0),
    f_bit8_width(C_PROBE_OUT205_WIDTH-1, (C_NUM_PROBE_OUT > 205), 0),
    f_bit8_width(C_PROBE_OUT204_WIDTH-1, (C_NUM_PROBE_OUT > 204), 0),
    f_bit8_width(C_PROBE_OUT203_WIDTH-1, (C_NUM_PROBE_OUT > 203), 0),
    f_bit8_width(C_PROBE_OUT202_WIDTH-1, (C_NUM_PROBE_OUT > 202), 0),
    f_bit8_width(C_PROBE_OUT201_WIDTH-1, (C_NUM_PROBE_OUT > 201), 0),
    f_bit8_width(C_PROBE_OUT200_WIDTH-1, (C_NUM_PROBE_OUT > 200), 0),
    f_bit8_width(C_PROBE_OUT199_WIDTH-1, (C_NUM_PROBE_OUT > 199), 0),
    f_bit8_width(C_PROBE_OUT198_WIDTH-1, (C_NUM_PROBE_OUT > 198), 0),
    f_bit8_width(C_PROBE_OUT197_WIDTH-1, (C_NUM_PROBE_OUT > 197), 0),
    f_bit8_width(C_PROBE_OUT196_WIDTH-1, (C_NUM_PROBE_OUT > 196), 0),
    f_bit8_width(C_PROBE_OUT195_WIDTH-1, (C_NUM_PROBE_OUT > 195), 0),
    f_bit8_width(C_PROBE_OUT194_WIDTH-1, (C_NUM_PROBE_OUT > 194), 0),
    f_bit8_width(C_PROBE_OUT193_WIDTH-1, (C_NUM_PROBE_OUT > 193), 0),
    f_bit8_width(C_PROBE_OUT192_WIDTH-1, (C_NUM_PROBE_OUT > 192), 0),
    f_bit8_width(C_PROBE_OUT191_WIDTH-1, (C_NUM_PROBE_OUT > 191), 0),
    f_bit8_width(C_PROBE_OUT190_WIDTH-1, (C_NUM_PROBE_OUT > 190), 0),
    f_bit8_width(C_PROBE_OUT189_WIDTH-1, (C_NUM_PROBE_OUT > 189), 0),
    f_bit8_width(C_PROBE_OUT188_WIDTH-1, (C_NUM_PROBE_OUT > 188), 0),
    f_bit8_width(C_PROBE_OUT187_WIDTH-1, (C_NUM_PROBE_OUT > 187), 0),
    f_bit8_width(C_PROBE_OUT186_WIDTH-1, (C_NUM_PROBE_OUT > 186), 0),
    f_bit8_width(C_PROBE_OUT185_WIDTH-1, (C_NUM_PROBE_OUT > 185), 0),
    f_bit8_width(C_PROBE_OUT184_WIDTH-1, (C_NUM_PROBE_OUT > 184), 0),
    f_bit8_width(C_PROBE_OUT183_WIDTH-1, (C_NUM_PROBE_OUT > 183), 0),
    f_bit8_width(C_PROBE_OUT182_WIDTH-1, (C_NUM_PROBE_OUT > 182), 0),
    f_bit8_width(C_PROBE_OUT181_WIDTH-1, (C_NUM_PROBE_OUT > 181), 0),
    f_bit8_width(C_PROBE_OUT180_WIDTH-1, (C_NUM_PROBE_OUT > 180), 0),
    f_bit8_width(C_PROBE_OUT179_WIDTH-1, (C_NUM_PROBE_OUT > 179), 0),
    f_bit8_width(C_PROBE_OUT178_WIDTH-1, (C_NUM_PROBE_OUT > 178), 0),
    f_bit8_width(C_PROBE_OUT177_WIDTH-1, (C_NUM_PROBE_OUT > 177), 0),
    f_bit8_width(C_PROBE_OUT176_WIDTH-1, (C_NUM_PROBE_OUT > 176), 0),
    f_bit8_width(C_PROBE_OUT175_WIDTH-1, (C_NUM_PROBE_OUT > 175), 0),
    f_bit8_width(C_PROBE_OUT174_WIDTH-1, (C_NUM_PROBE_OUT > 174), 0),
    f_bit8_width(C_PROBE_OUT173_WIDTH-1, (C_NUM_PROBE_OUT > 173), 0),
    f_bit8_width(C_PROBE_OUT172_WIDTH-1, (C_NUM_PROBE_OUT > 172), 0),
    f_bit8_width(C_PROBE_OUT171_WIDTH-1, (C_NUM_PROBE_OUT > 171), 0),
    f_bit8_width(C_PROBE_OUT170_WIDTH-1, (C_NUM_PROBE_OUT > 170), 0),
    f_bit8_width(C_PROBE_OUT169_WIDTH-1, (C_NUM_PROBE_OUT > 169), 0),
    f_bit8_width(C_PROBE_OUT168_WIDTH-1, (C_NUM_PROBE_OUT > 168), 0),
    f_bit8_width(C_PROBE_OUT167_WIDTH-1, (C_NUM_PROBE_OUT > 167), 0),
    f_bit8_width(C_PROBE_OUT166_WIDTH-1, (C_NUM_PROBE_OUT > 166), 0),
    f_bit8_width(C_PROBE_OUT165_WIDTH-1, (C_NUM_PROBE_OUT > 165), 0),
    f_bit8_width(C_PROBE_OUT164_WIDTH-1, (C_NUM_PROBE_OUT > 164), 0),
    f_bit8_width(C_PROBE_OUT163_WIDTH-1, (C_NUM_PROBE_OUT > 163), 0),
    f_bit8_width(C_PROBE_OUT162_WIDTH-1, (C_NUM_PROBE_OUT > 162), 0),
    f_bit8_width(C_PROBE_OUT161_WIDTH-1, (C_NUM_PROBE_OUT > 161), 0),
    f_bit8_width(C_PROBE_OUT160_WIDTH-1, (C_NUM_PROBE_OUT > 160), 0),
    f_bit8_width(C_PROBE_OUT159_WIDTH-1, (C_NUM_PROBE_OUT > 159), 0),
    f_bit8_width(C_PROBE_OUT158_WIDTH-1, (C_NUM_PROBE_OUT > 158), 0),
    f_bit8_width(C_PROBE_OUT157_WIDTH-1, (C_NUM_PROBE_OUT > 157), 0),
    f_bit8_width(C_PROBE_OUT156_WIDTH-1, (C_NUM_PROBE_OUT > 156), 0),
    f_bit8_width(C_PROBE_OUT155_WIDTH-1, (C_NUM_PROBE_OUT > 155), 0),
    f_bit8_width(C_PROBE_OUT154_WIDTH-1, (C_NUM_PROBE_OUT > 154), 0),
    f_bit8_width(C_PROBE_OUT153_WIDTH-1, (C_NUM_PROBE_OUT > 153), 0),
    f_bit8_width(C_PROBE_OUT152_WIDTH-1, (C_NUM_PROBE_OUT > 152), 0),
    f_bit8_width(C_PROBE_OUT151_WIDTH-1, (C_NUM_PROBE_OUT > 151), 0),
    f_bit8_width(C_PROBE_OUT150_WIDTH-1, (C_NUM_PROBE_OUT > 150), 0),
    f_bit8_width(C_PROBE_OUT149_WIDTH-1, (C_NUM_PROBE_OUT > 149), 0),
    f_bit8_width(C_PROBE_OUT148_WIDTH-1, (C_NUM_PROBE_OUT > 148), 0),
    f_bit8_width(C_PROBE_OUT147_WIDTH-1, (C_NUM_PROBE_OUT > 147), 0),
    f_bit8_width(C_PROBE_OUT146_WIDTH-1, (C_NUM_PROBE_OUT > 146), 0),
    f_bit8_width(C_PROBE_OUT145_WIDTH-1, (C_NUM_PROBE_OUT > 145), 0),
    f_bit8_width(C_PROBE_OUT144_WIDTH-1, (C_NUM_PROBE_OUT > 144), 0),
    f_bit8_width(C_PROBE_OUT143_WIDTH-1, (C_NUM_PROBE_OUT > 143), 0),
    f_bit8_width(C_PROBE_OUT142_WIDTH-1, (C_NUM_PROBE_OUT > 142), 0),
    f_bit8_width(C_PROBE_OUT141_WIDTH-1, (C_NUM_PROBE_OUT > 141), 0),
    f_bit8_width(C_PROBE_OUT140_WIDTH-1, (C_NUM_PROBE_OUT > 140), 0),
    f_bit8_width(C_PROBE_OUT139_WIDTH-1, (C_NUM_PROBE_OUT > 139), 0),
    f_bit8_width(C_PROBE_OUT138_WIDTH-1, (C_NUM_PROBE_OUT > 138), 0),
    f_bit8_width(C_PROBE_OUT137_WIDTH-1, (C_NUM_PROBE_OUT > 137), 0),
    f_bit8_width(C_PROBE_OUT136_WIDTH-1, (C_NUM_PROBE_OUT > 136), 0),
    f_bit8_width(C_PROBE_OUT135_WIDTH-1, (C_NUM_PROBE_OUT > 135), 0),
    f_bit8_width(C_PROBE_OUT134_WIDTH-1, (C_NUM_PROBE_OUT > 134), 0),
    f_bit8_width(C_PROBE_OUT133_WIDTH-1, (C_NUM_PROBE_OUT > 133), 0),
    f_bit8_width(C_PROBE_OUT132_WIDTH-1, (C_NUM_PROBE_OUT > 132), 0),
    f_bit8_width(C_PROBE_OUT131_WIDTH-1, (C_NUM_PROBE_OUT > 131), 0),
    f_bit8_width(C_PROBE_OUT130_WIDTH-1, (C_NUM_PROBE_OUT > 130), 0),
    f_bit8_width(C_PROBE_OUT129_WIDTH-1, (C_NUM_PROBE_OUT > 129), 0),
    f_bit8_width(C_PROBE_OUT128_WIDTH-1, (C_NUM_PROBE_OUT > 128), 0),
    f_bit8_width(C_PROBE_OUT127_WIDTH-1, (C_NUM_PROBE_OUT > 127), 0),
    f_bit8_width(C_PROBE_OUT126_WIDTH-1, (C_NUM_PROBE_OUT > 126), 0),
    f_bit8_width(C_PROBE_OUT125_WIDTH-1, (C_NUM_PROBE_OUT > 125), 0),
    f_bit8_width(C_PROBE_OUT124_WIDTH-1, (C_NUM_PROBE_OUT > 124), 0),
    f_bit8_width(C_PROBE_OUT123_WIDTH-1, (C_NUM_PROBE_OUT > 123), 0),
    f_bit8_width(C_PROBE_OUT122_WIDTH-1, (C_NUM_PROBE_OUT > 122), 0),
    f_bit8_width(C_PROBE_OUT121_WIDTH-1, (C_NUM_PROBE_OUT > 121), 0),
    f_bit8_width(C_PROBE_OUT120_WIDTH-1, (C_NUM_PROBE_OUT > 120), 0),
    f_bit8_width(C_PROBE_OUT119_WIDTH-1, (C_NUM_PROBE_OUT > 119), 0),
    f_bit8_width(C_PROBE_OUT118_WIDTH-1, (C_NUM_PROBE_OUT > 118), 0),
    f_bit8_width(C_PROBE_OUT117_WIDTH-1, (C_NUM_PROBE_OUT > 117), 0),
    f_bit8_width(C_PROBE_OUT116_WIDTH-1, (C_NUM_PROBE_OUT > 116), 0),
    f_bit8_width(C_PROBE_OUT115_WIDTH-1, (C_NUM_PROBE_OUT > 115), 0),
    f_bit8_width(C_PROBE_OUT114_WIDTH-1, (C_NUM_PROBE_OUT > 114), 0),
    f_bit8_width(C_PROBE_OUT113_WIDTH-1, (C_NUM_PROBE_OUT > 113), 0),
    f_bit8_width(C_PROBE_OUT112_WIDTH-1, (C_NUM_PROBE_OUT > 112), 0),
    f_bit8_width(C_PROBE_OUT111_WIDTH-1, (C_NUM_PROBE_OUT > 111), 0),
    f_bit8_width(C_PROBE_OUT110_WIDTH-1, (C_NUM_PROBE_OUT > 110), 0),
    f_bit8_width(C_PROBE_OUT109_WIDTH-1, (C_NUM_PROBE_OUT > 109), 0),
    f_bit8_width(C_PROBE_OUT108_WIDTH-1, (C_NUM_PROBE_OUT > 108), 0),
    f_bit8_width(C_PROBE_OUT107_WIDTH-1, (C_NUM_PROBE_OUT > 107), 0),
    f_bit8_width(C_PROBE_OUT106_WIDTH-1, (C_NUM_PROBE_OUT > 106), 0),
    f_bit8_width(C_PROBE_OUT105_WIDTH-1, (C_NUM_PROBE_OUT > 105), 0),
    f_bit8_width(C_PROBE_OUT104_WIDTH-1, (C_NUM_PROBE_OUT > 104), 0),
    f_bit8_width(C_PROBE_OUT103_WIDTH-1, (C_NUM_PROBE_OUT > 103), 0),
    f_bit8_width(C_PROBE_OUT102_WIDTH-1, (C_NUM_PROBE_OUT > 102), 0),
    f_bit8_width(C_PROBE_OUT101_WIDTH-1, (C_NUM_PROBE_OUT > 101), 0),
    f_bit8_width(C_PROBE_OUT100_WIDTH-1, (C_NUM_PROBE_OUT > 100), 0),
    f_bit8_width(C_PROBE_OUT99_WIDTH-1 , (C_NUM_PROBE_OUT > 99), 0),
    f_bit8_width(C_PROBE_OUT98_WIDTH-1 , (C_NUM_PROBE_OUT > 98), 0),
    f_bit8_width(C_PROBE_OUT97_WIDTH-1 , (C_NUM_PROBE_OUT > 97), 0),
    f_bit8_width(C_PROBE_OUT96_WIDTH-1 , (C_NUM_PROBE_OUT > 96), 0),
    f_bit8_width(C_PROBE_OUT95_WIDTH-1 , (C_NUM_PROBE_OUT > 95), 0),
    f_bit8_width(C_PROBE_OUT94_WIDTH-1 , (C_NUM_PROBE_OUT > 94), 0),
    f_bit8_width(C_PROBE_OUT93_WIDTH-1 , (C_NUM_PROBE_OUT > 93), 0),
    f_bit8_width(C_PROBE_OUT92_WIDTH-1 , (C_NUM_PROBE_OUT > 92), 0),
    f_bit8_width(C_PROBE_OUT91_WIDTH-1 , (C_NUM_PROBE_OUT > 91), 0),
    f_bit8_width(C_PROBE_OUT90_WIDTH-1 , (C_NUM_PROBE_OUT > 90), 0),
    f_bit8_width(C_PROBE_OUT89_WIDTH-1 , (C_NUM_PROBE_OUT > 89), 0),
    f_bit8_width(C_PROBE_OUT88_WIDTH-1 , (C_NUM_PROBE_OUT > 88), 0),
    f_bit8_width(C_PROBE_OUT87_WIDTH-1 , (C_NUM_PROBE_OUT > 87), 0),
    f_bit8_width(C_PROBE_OUT86_WIDTH-1 , (C_NUM_PROBE_OUT > 86), 0),
    f_bit8_width(C_PROBE_OUT85_WIDTH-1 , (C_NUM_PROBE_OUT > 85), 0),
    f_bit8_width(C_PROBE_OUT84_WIDTH-1 , (C_NUM_PROBE_OUT > 84), 0),
    f_bit8_width(C_PROBE_OUT83_WIDTH-1 , (C_NUM_PROBE_OUT > 83), 0),
    f_bit8_width(C_PROBE_OUT82_WIDTH-1 , (C_NUM_PROBE_OUT > 82), 0),
    f_bit8_width(C_PROBE_OUT81_WIDTH-1 , (C_NUM_PROBE_OUT > 81), 0),
    f_bit8_width(C_PROBE_OUT80_WIDTH-1 , (C_NUM_PROBE_OUT > 80), 0),
    f_bit8_width(C_PROBE_OUT79_WIDTH-1 , (C_NUM_PROBE_OUT > 79), 0),
    f_bit8_width(C_PROBE_OUT78_WIDTH-1 , (C_NUM_PROBE_OUT > 78), 0),
    f_bit8_width(C_PROBE_OUT77_WIDTH-1 , (C_NUM_PROBE_OUT > 77), 0),
    f_bit8_width(C_PROBE_OUT76_WIDTH-1 , (C_NUM_PROBE_OUT > 76), 0),
    f_bit8_width(C_PROBE_OUT75_WIDTH-1 , (C_NUM_PROBE_OUT > 75), 0),
    f_bit8_width(C_PROBE_OUT74_WIDTH-1 , (C_NUM_PROBE_OUT > 74), 0),
    f_bit8_width(C_PROBE_OUT73_WIDTH-1 , (C_NUM_PROBE_OUT > 73), 0),
    f_bit8_width(C_PROBE_OUT72_WIDTH-1 , (C_NUM_PROBE_OUT > 72), 0),
    f_bit8_width(C_PROBE_OUT71_WIDTH-1 , (C_NUM_PROBE_OUT > 71), 0),
    f_bit8_width(C_PROBE_OUT70_WIDTH-1 , (C_NUM_PROBE_OUT > 70), 0),
    f_bit8_width(C_PROBE_OUT69_WIDTH-1 , (C_NUM_PROBE_OUT > 69), 0),
    f_bit8_width(C_PROBE_OUT68_WIDTH-1 , (C_NUM_PROBE_OUT > 68), 0),
    f_bit8_width(C_PROBE_OUT67_WIDTH-1 , (C_NUM_PROBE_OUT > 67), 0),
    f_bit8_width(C_PROBE_OUT66_WIDTH-1 , (C_NUM_PROBE_OUT > 66), 0),
    f_bit8_width(C_PROBE_OUT65_WIDTH-1 , (C_NUM_PROBE_OUT > 65), 0),
    f_bit8_width(C_PROBE_OUT64_WIDTH-1 , (C_NUM_PROBE_OUT > 64), 0),
    f_bit8_width(C_PROBE_OUT63_WIDTH-1 , (C_NUM_PROBE_OUT > 63), 0),
    f_bit8_width(C_PROBE_OUT62_WIDTH-1 , (C_NUM_PROBE_OUT > 62), 0),
    f_bit8_width(C_PROBE_OUT61_WIDTH-1 , (C_NUM_PROBE_OUT > 61), 0),
    f_bit8_width(C_PROBE_OUT60_WIDTH-1 , (C_NUM_PROBE_OUT > 60), 0),
    f_bit8_width(C_PROBE_OUT59_WIDTH-1 , (C_NUM_PROBE_OUT > 59), 0),
    f_bit8_width(C_PROBE_OUT58_WIDTH-1 , (C_NUM_PROBE_OUT > 58), 0),
    f_bit8_width(C_PROBE_OUT57_WIDTH-1 , (C_NUM_PROBE_OUT > 57), 0),
    f_bit8_width(C_PROBE_OUT56_WIDTH-1 , (C_NUM_PROBE_OUT > 56), 0),
    f_bit8_width(C_PROBE_OUT55_WIDTH-1 , (C_NUM_PROBE_OUT > 55), 0),
    f_bit8_width(C_PROBE_OUT54_WIDTH-1 , (C_NUM_PROBE_OUT > 54), 0),
    f_bit8_width(C_PROBE_OUT53_WIDTH-1 , (C_NUM_PROBE_OUT > 53), 0),
    f_bit8_width(C_PROBE_OUT52_WIDTH-1 , (C_NUM_PROBE_OUT > 52), 0),
    f_bit8_width(C_PROBE_OUT51_WIDTH-1 , (C_NUM_PROBE_OUT > 51), 0),
    f_bit8_width(C_PROBE_OUT50_WIDTH-1 , (C_NUM_PROBE_OUT > 50), 0),
    f_bit8_width(C_PROBE_OUT49_WIDTH-1 , (C_NUM_PROBE_OUT > 49), 0),
    f_bit8_width(C_PROBE_OUT48_WIDTH-1 , (C_NUM_PROBE_OUT > 48), 0),
    f_bit8_width(C_PROBE_OUT47_WIDTH-1 , (C_NUM_PROBE_OUT > 47), 0),
    f_bit8_width(C_PROBE_OUT46_WIDTH-1 , (C_NUM_PROBE_OUT > 46), 0),
    f_bit8_width(C_PROBE_OUT45_WIDTH-1 , (C_NUM_PROBE_OUT > 45), 0),
    f_bit8_width(C_PROBE_OUT44_WIDTH-1 , (C_NUM_PROBE_OUT > 44), 0),
    f_bit8_width(C_PROBE_OUT43_WIDTH-1 , (C_NUM_PROBE_OUT > 43), 0),
    f_bit8_width(C_PROBE_OUT42_WIDTH-1 , (C_NUM_PROBE_OUT > 42), 0),
    f_bit8_width(C_PROBE_OUT41_WIDTH-1 , (C_NUM_PROBE_OUT > 41), 0),
    f_bit8_width(C_PROBE_OUT40_WIDTH-1 , (C_NUM_PROBE_OUT > 40), 0),
    f_bit8_width(C_PROBE_OUT39_WIDTH-1 , (C_NUM_PROBE_OUT > 39), 0),
    f_bit8_width(C_PROBE_OUT38_WIDTH-1 , (C_NUM_PROBE_OUT > 38), 0),
    f_bit8_width(C_PROBE_OUT37_WIDTH-1 , (C_NUM_PROBE_OUT > 37), 0),
    f_bit8_width(C_PROBE_OUT36_WIDTH-1 , (C_NUM_PROBE_OUT > 36), 0),
    f_bit8_width(C_PROBE_OUT35_WIDTH-1 , (C_NUM_PROBE_OUT > 35), 0),
    f_bit8_width(C_PROBE_OUT34_WIDTH-1 , (C_NUM_PROBE_OUT > 34), 0),
    f_bit8_width(C_PROBE_OUT33_WIDTH-1 , (C_NUM_PROBE_OUT > 33), 0),
    f_bit8_width(C_PROBE_OUT32_WIDTH-1 , (C_NUM_PROBE_OUT > 32), 0),
    f_bit8_width(C_PROBE_OUT31_WIDTH-1 , (C_NUM_PROBE_OUT > 31), 0),
    f_bit8_width(C_PROBE_OUT30_WIDTH-1 , (C_NUM_PROBE_OUT > 30), 0),
    f_bit8_width(C_PROBE_OUT29_WIDTH-1 , (C_NUM_PROBE_OUT > 29), 0),
    f_bit8_width(C_PROBE_OUT28_WIDTH-1 , (C_NUM_PROBE_OUT > 28), 0),
    f_bit8_width(C_PROBE_OUT27_WIDTH-1 , (C_NUM_PROBE_OUT > 27), 0),
    f_bit8_width(C_PROBE_OUT26_WIDTH-1 , (C_NUM_PROBE_OUT > 26), 0),
    f_bit8_width(C_PROBE_OUT25_WIDTH-1 , (C_NUM_PROBE_OUT > 25), 0),
    f_bit8_width(C_PROBE_OUT24_WIDTH-1 , (C_NUM_PROBE_OUT > 24), 0),
    f_bit8_width(C_PROBE_OUT23_WIDTH-1 , (C_NUM_PROBE_OUT > 23), 0),
    f_bit8_width(C_PROBE_OUT22_WIDTH-1 , (C_NUM_PROBE_OUT > 22), 0),
    f_bit8_width(C_PROBE_OUT21_WIDTH-1 , (C_NUM_PROBE_OUT > 21), 0),
    f_bit8_width(C_PROBE_OUT20_WIDTH-1 , (C_NUM_PROBE_OUT > 20), 0),
    f_bit8_width(C_PROBE_OUT19_WIDTH-1 , (C_NUM_PROBE_OUT > 19), 0),
    f_bit8_width(C_PROBE_OUT18_WIDTH-1 , (C_NUM_PROBE_OUT > 18), 0),
    f_bit8_width(C_PROBE_OUT17_WIDTH-1 , (C_NUM_PROBE_OUT > 17), 0),
    f_bit8_width(C_PROBE_OUT16_WIDTH-1 , (C_NUM_PROBE_OUT > 16), 0),
    f_bit8_width(C_PROBE_OUT15_WIDTH-1 , (C_NUM_PROBE_OUT > 15), 0),
    f_bit8_width(C_PROBE_OUT14_WIDTH-1 , (C_NUM_PROBE_OUT > 14), 0),
    f_bit8_width(C_PROBE_OUT13_WIDTH-1 , (C_NUM_PROBE_OUT > 13), 0),
    f_bit8_width(C_PROBE_OUT12_WIDTH-1 , (C_NUM_PROBE_OUT > 12), 0),
    f_bit8_width(C_PROBE_OUT11_WIDTH-1 , (C_NUM_PROBE_OUT > 11), 0),
    f_bit8_width(C_PROBE_OUT10_WIDTH-1 , (C_NUM_PROBE_OUT > 10), 0),
    f_bit8_width(C_PROBE_OUT9_WIDTH-1  , (C_NUM_PROBE_OUT >  9), 0),
    f_bit8_width(C_PROBE_OUT8_WIDTH-1  , (C_NUM_PROBE_OUT >  8), 0),
    f_bit8_width(C_PROBE_OUT7_WIDTH-1  , (C_NUM_PROBE_OUT >  7), 0),
    f_bit8_width(C_PROBE_OUT6_WIDTH-1  , (C_NUM_PROBE_OUT >  6), 0),
    f_bit8_width(C_PROBE_OUT5_WIDTH-1  , (C_NUM_PROBE_OUT >  5), 0),
    f_bit8_width(C_PROBE_OUT4_WIDTH-1  , (C_NUM_PROBE_OUT >  4), 0),
    f_bit8_width(C_PROBE_OUT3_WIDTH-1  , (C_NUM_PROBE_OUT >  3), 0),
    f_bit8_width(C_PROBE_OUT2_WIDTH-1  , (C_NUM_PROBE_OUT >  2), 0),
    f_bit8_width(C_PROBE_OUT1_WIDTH-1  , (C_NUM_PROBE_OUT >  1), 0),
    f_bit8_width(C_PROBE_OUT0_WIDTH-1  , (C_NUM_PROBE_OUT >  0), 0)
  };

  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT0   = C_PROBE_OUT0_WIDTH           - 1                   ;	        
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT1   = LC_HIGH_BIT_POS_PROBE_OUT0   + C_PROBE_OUT1_WIDTH  ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT2   = LC_HIGH_BIT_POS_PROBE_OUT1   + C_PROBE_OUT2_WIDTH  ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT3   = LC_HIGH_BIT_POS_PROBE_OUT2   + C_PROBE_OUT3_WIDTH  ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT4   = LC_HIGH_BIT_POS_PROBE_OUT3   + C_PROBE_OUT4_WIDTH  ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT5   = LC_HIGH_BIT_POS_PROBE_OUT4   + C_PROBE_OUT5_WIDTH  ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT6   = LC_HIGH_BIT_POS_PROBE_OUT5   + C_PROBE_OUT6_WIDTH  ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT7   = LC_HIGH_BIT_POS_PROBE_OUT6   + C_PROBE_OUT7_WIDTH  ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT8   = LC_HIGH_BIT_POS_PROBE_OUT7   + C_PROBE_OUT8_WIDTH  ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT9   = LC_HIGH_BIT_POS_PROBE_OUT8   + C_PROBE_OUT9_WIDTH  ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT10  = LC_HIGH_BIT_POS_PROBE_OUT9   + C_PROBE_OUT10_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT11  = LC_HIGH_BIT_POS_PROBE_OUT10  + C_PROBE_OUT11_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT12  = LC_HIGH_BIT_POS_PROBE_OUT11  + C_PROBE_OUT12_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT13  = LC_HIGH_BIT_POS_PROBE_OUT12  + C_PROBE_OUT13_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT14  = LC_HIGH_BIT_POS_PROBE_OUT13  + C_PROBE_OUT14_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT15  = LC_HIGH_BIT_POS_PROBE_OUT14  + C_PROBE_OUT15_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT16  = LC_HIGH_BIT_POS_PROBE_OUT15  + C_PROBE_OUT16_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT17  = LC_HIGH_BIT_POS_PROBE_OUT16  + C_PROBE_OUT17_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT18  = LC_HIGH_BIT_POS_PROBE_OUT17  + C_PROBE_OUT18_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT19  = LC_HIGH_BIT_POS_PROBE_OUT18  + C_PROBE_OUT19_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT20  = LC_HIGH_BIT_POS_PROBE_OUT19  + C_PROBE_OUT20_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT21  = LC_HIGH_BIT_POS_PROBE_OUT20  + C_PROBE_OUT21_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT22  = LC_HIGH_BIT_POS_PROBE_OUT21  + C_PROBE_OUT22_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT23  = LC_HIGH_BIT_POS_PROBE_OUT22  + C_PROBE_OUT23_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT24  = LC_HIGH_BIT_POS_PROBE_OUT23  + C_PROBE_OUT24_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT25  = LC_HIGH_BIT_POS_PROBE_OUT24  + C_PROBE_OUT25_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT26  = LC_HIGH_BIT_POS_PROBE_OUT25  + C_PROBE_OUT26_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT27  = LC_HIGH_BIT_POS_PROBE_OUT26  + C_PROBE_OUT27_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT28  = LC_HIGH_BIT_POS_PROBE_OUT27  + C_PROBE_OUT28_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT29  = LC_HIGH_BIT_POS_PROBE_OUT28  + C_PROBE_OUT29_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT30  = LC_HIGH_BIT_POS_PROBE_OUT29  + C_PROBE_OUT30_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT31  = LC_HIGH_BIT_POS_PROBE_OUT30  + C_PROBE_OUT31_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT32  = LC_HIGH_BIT_POS_PROBE_OUT31  + C_PROBE_OUT32_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT33  = LC_HIGH_BIT_POS_PROBE_OUT32  + C_PROBE_OUT33_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT34  = LC_HIGH_BIT_POS_PROBE_OUT33  + C_PROBE_OUT34_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT35  = LC_HIGH_BIT_POS_PROBE_OUT34  + C_PROBE_OUT35_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT36  = LC_HIGH_BIT_POS_PROBE_OUT35  + C_PROBE_OUT36_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT37  = LC_HIGH_BIT_POS_PROBE_OUT36  + C_PROBE_OUT37_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT38  = LC_HIGH_BIT_POS_PROBE_OUT37  + C_PROBE_OUT38_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT39  = LC_HIGH_BIT_POS_PROBE_OUT38  + C_PROBE_OUT39_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT40  = LC_HIGH_BIT_POS_PROBE_OUT39  + C_PROBE_OUT40_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT41  = LC_HIGH_BIT_POS_PROBE_OUT40  + C_PROBE_OUT41_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT42  = LC_HIGH_BIT_POS_PROBE_OUT41  + C_PROBE_OUT42_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT43  = LC_HIGH_BIT_POS_PROBE_OUT42  + C_PROBE_OUT43_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT44  = LC_HIGH_BIT_POS_PROBE_OUT43  + C_PROBE_OUT44_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT45  = LC_HIGH_BIT_POS_PROBE_OUT44  + C_PROBE_OUT45_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT46  = LC_HIGH_BIT_POS_PROBE_OUT45  + C_PROBE_OUT46_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT47  = LC_HIGH_BIT_POS_PROBE_OUT46  + C_PROBE_OUT47_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT48  = LC_HIGH_BIT_POS_PROBE_OUT47  + C_PROBE_OUT48_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT49  = LC_HIGH_BIT_POS_PROBE_OUT48  + C_PROBE_OUT49_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT50  = LC_HIGH_BIT_POS_PROBE_OUT49  + C_PROBE_OUT50_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT51  = LC_HIGH_BIT_POS_PROBE_OUT50  + C_PROBE_OUT51_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT52  = LC_HIGH_BIT_POS_PROBE_OUT51  + C_PROBE_OUT52_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT53  = LC_HIGH_BIT_POS_PROBE_OUT52  + C_PROBE_OUT53_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT54  = LC_HIGH_BIT_POS_PROBE_OUT53  + C_PROBE_OUT54_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT55  = LC_HIGH_BIT_POS_PROBE_OUT54  + C_PROBE_OUT55_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT56  = LC_HIGH_BIT_POS_PROBE_OUT55  + C_PROBE_OUT56_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT57  = LC_HIGH_BIT_POS_PROBE_OUT56  + C_PROBE_OUT57_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT58  = LC_HIGH_BIT_POS_PROBE_OUT57  + C_PROBE_OUT58_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT59  = LC_HIGH_BIT_POS_PROBE_OUT58  + C_PROBE_OUT59_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT60  = LC_HIGH_BIT_POS_PROBE_OUT59  + C_PROBE_OUT60_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT61  = LC_HIGH_BIT_POS_PROBE_OUT60  + C_PROBE_OUT61_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT62  = LC_HIGH_BIT_POS_PROBE_OUT61  + C_PROBE_OUT62_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT63  = LC_HIGH_BIT_POS_PROBE_OUT62  + C_PROBE_OUT63_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT64  = LC_HIGH_BIT_POS_PROBE_OUT63  + C_PROBE_OUT64_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT65  = LC_HIGH_BIT_POS_PROBE_OUT64  + C_PROBE_OUT65_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT66  = LC_HIGH_BIT_POS_PROBE_OUT65  + C_PROBE_OUT66_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT67  = LC_HIGH_BIT_POS_PROBE_OUT66  + C_PROBE_OUT67_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT68  = LC_HIGH_BIT_POS_PROBE_OUT67  + C_PROBE_OUT68_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT69  = LC_HIGH_BIT_POS_PROBE_OUT68  + C_PROBE_OUT69_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT70  = LC_HIGH_BIT_POS_PROBE_OUT69  + C_PROBE_OUT70_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT71  = LC_HIGH_BIT_POS_PROBE_OUT70  + C_PROBE_OUT71_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT72  = LC_HIGH_BIT_POS_PROBE_OUT71  + C_PROBE_OUT72_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT73  = LC_HIGH_BIT_POS_PROBE_OUT72  + C_PROBE_OUT73_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT74  = LC_HIGH_BIT_POS_PROBE_OUT73  + C_PROBE_OUT74_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT75  = LC_HIGH_BIT_POS_PROBE_OUT74  + C_PROBE_OUT75_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT76  = LC_HIGH_BIT_POS_PROBE_OUT75  + C_PROBE_OUT76_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT77  = LC_HIGH_BIT_POS_PROBE_OUT76  + C_PROBE_OUT77_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT78  = LC_HIGH_BIT_POS_PROBE_OUT77  + C_PROBE_OUT78_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT79  = LC_HIGH_BIT_POS_PROBE_OUT78  + C_PROBE_OUT79_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT80  = LC_HIGH_BIT_POS_PROBE_OUT79  + C_PROBE_OUT80_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT81  = LC_HIGH_BIT_POS_PROBE_OUT80  + C_PROBE_OUT81_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT82  = LC_HIGH_BIT_POS_PROBE_OUT81  + C_PROBE_OUT82_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT83  = LC_HIGH_BIT_POS_PROBE_OUT82  + C_PROBE_OUT83_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT84  = LC_HIGH_BIT_POS_PROBE_OUT83  + C_PROBE_OUT84_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT85  = LC_HIGH_BIT_POS_PROBE_OUT84  + C_PROBE_OUT85_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT86  = LC_HIGH_BIT_POS_PROBE_OUT85  + C_PROBE_OUT86_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT87  = LC_HIGH_BIT_POS_PROBE_OUT86  + C_PROBE_OUT87_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT88  = LC_HIGH_BIT_POS_PROBE_OUT87  + C_PROBE_OUT88_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT89  = LC_HIGH_BIT_POS_PROBE_OUT88  + C_PROBE_OUT89_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT90  = LC_HIGH_BIT_POS_PROBE_OUT89  + C_PROBE_OUT90_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT91  = LC_HIGH_BIT_POS_PROBE_OUT90  + C_PROBE_OUT91_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT92  = LC_HIGH_BIT_POS_PROBE_OUT91  + C_PROBE_OUT92_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT93  = LC_HIGH_BIT_POS_PROBE_OUT92  + C_PROBE_OUT93_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT94  = LC_HIGH_BIT_POS_PROBE_OUT93  + C_PROBE_OUT94_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT95  = LC_HIGH_BIT_POS_PROBE_OUT94  + C_PROBE_OUT95_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT96  = LC_HIGH_BIT_POS_PROBE_OUT95  + C_PROBE_OUT96_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT97  = LC_HIGH_BIT_POS_PROBE_OUT96  + C_PROBE_OUT97_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT98  = LC_HIGH_BIT_POS_PROBE_OUT97  + C_PROBE_OUT98_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT99  = LC_HIGH_BIT_POS_PROBE_OUT98  + C_PROBE_OUT99_WIDTH ;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT100 = LC_HIGH_BIT_POS_PROBE_OUT99  + C_PROBE_OUT100_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT101 = LC_HIGH_BIT_POS_PROBE_OUT100 + C_PROBE_OUT101_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT102 = LC_HIGH_BIT_POS_PROBE_OUT101 + C_PROBE_OUT102_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT103 = LC_HIGH_BIT_POS_PROBE_OUT102 + C_PROBE_OUT103_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT104 = LC_HIGH_BIT_POS_PROBE_OUT103 + C_PROBE_OUT104_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT105 = LC_HIGH_BIT_POS_PROBE_OUT104 + C_PROBE_OUT105_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT106 = LC_HIGH_BIT_POS_PROBE_OUT105 + C_PROBE_OUT106_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT107 = LC_HIGH_BIT_POS_PROBE_OUT106 + C_PROBE_OUT107_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT108 = LC_HIGH_BIT_POS_PROBE_OUT107 + C_PROBE_OUT108_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT109 = LC_HIGH_BIT_POS_PROBE_OUT108 + C_PROBE_OUT109_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT110 = LC_HIGH_BIT_POS_PROBE_OUT109 + C_PROBE_OUT110_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT111 = LC_HIGH_BIT_POS_PROBE_OUT110 + C_PROBE_OUT111_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT112 = LC_HIGH_BIT_POS_PROBE_OUT111 + C_PROBE_OUT112_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT113 = LC_HIGH_BIT_POS_PROBE_OUT112 + C_PROBE_OUT113_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT114 = LC_HIGH_BIT_POS_PROBE_OUT113 + C_PROBE_OUT114_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT115 = LC_HIGH_BIT_POS_PROBE_OUT114 + C_PROBE_OUT115_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT116 = LC_HIGH_BIT_POS_PROBE_OUT115 + C_PROBE_OUT116_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT117 = LC_HIGH_BIT_POS_PROBE_OUT116 + C_PROBE_OUT117_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT118 = LC_HIGH_BIT_POS_PROBE_OUT117 + C_PROBE_OUT118_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT119 = LC_HIGH_BIT_POS_PROBE_OUT118 + C_PROBE_OUT119_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT120 = LC_HIGH_BIT_POS_PROBE_OUT119 + C_PROBE_OUT120_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT121 = LC_HIGH_BIT_POS_PROBE_OUT120 + C_PROBE_OUT121_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT122 = LC_HIGH_BIT_POS_PROBE_OUT121 + C_PROBE_OUT122_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT123 = LC_HIGH_BIT_POS_PROBE_OUT122 + C_PROBE_OUT123_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT124 = LC_HIGH_BIT_POS_PROBE_OUT123 + C_PROBE_OUT124_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT125 = LC_HIGH_BIT_POS_PROBE_OUT124 + C_PROBE_OUT125_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT126 = LC_HIGH_BIT_POS_PROBE_OUT125 + C_PROBE_OUT126_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT127 = LC_HIGH_BIT_POS_PROBE_OUT126 + C_PROBE_OUT127_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT128 = LC_HIGH_BIT_POS_PROBE_OUT127 + C_PROBE_OUT128_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT129 = LC_HIGH_BIT_POS_PROBE_OUT128 + C_PROBE_OUT129_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT130 = LC_HIGH_BIT_POS_PROBE_OUT129 + C_PROBE_OUT130_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT131 = LC_HIGH_BIT_POS_PROBE_OUT130 + C_PROBE_OUT131_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT132 = LC_HIGH_BIT_POS_PROBE_OUT131 + C_PROBE_OUT132_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT133 = LC_HIGH_BIT_POS_PROBE_OUT132 + C_PROBE_OUT133_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT134 = LC_HIGH_BIT_POS_PROBE_OUT133 + C_PROBE_OUT134_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT135 = LC_HIGH_BIT_POS_PROBE_OUT134 + C_PROBE_OUT135_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT136 = LC_HIGH_BIT_POS_PROBE_OUT135 + C_PROBE_OUT136_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT137 = LC_HIGH_BIT_POS_PROBE_OUT136 + C_PROBE_OUT137_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT138 = LC_HIGH_BIT_POS_PROBE_OUT137 + C_PROBE_OUT138_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT139 = LC_HIGH_BIT_POS_PROBE_OUT138 + C_PROBE_OUT139_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT140 = LC_HIGH_BIT_POS_PROBE_OUT139 + C_PROBE_OUT140_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT141 = LC_HIGH_BIT_POS_PROBE_OUT140 + C_PROBE_OUT141_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT142 = LC_HIGH_BIT_POS_PROBE_OUT141 + C_PROBE_OUT142_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT143 = LC_HIGH_BIT_POS_PROBE_OUT142 + C_PROBE_OUT143_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT144 = LC_HIGH_BIT_POS_PROBE_OUT143 + C_PROBE_OUT144_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT145 = LC_HIGH_BIT_POS_PROBE_OUT144 + C_PROBE_OUT145_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT146 = LC_HIGH_BIT_POS_PROBE_OUT145 + C_PROBE_OUT146_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT147 = LC_HIGH_BIT_POS_PROBE_OUT146 + C_PROBE_OUT147_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT148 = LC_HIGH_BIT_POS_PROBE_OUT147 + C_PROBE_OUT148_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT149 = LC_HIGH_BIT_POS_PROBE_OUT148 + C_PROBE_OUT149_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT150 = LC_HIGH_BIT_POS_PROBE_OUT149 + C_PROBE_OUT150_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT151 = LC_HIGH_BIT_POS_PROBE_OUT150 + C_PROBE_OUT151_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT152 = LC_HIGH_BIT_POS_PROBE_OUT151 + C_PROBE_OUT152_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT153 = LC_HIGH_BIT_POS_PROBE_OUT152 + C_PROBE_OUT153_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT154 = LC_HIGH_BIT_POS_PROBE_OUT153 + C_PROBE_OUT154_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT155 = LC_HIGH_BIT_POS_PROBE_OUT154 + C_PROBE_OUT155_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT156 = LC_HIGH_BIT_POS_PROBE_OUT155 + C_PROBE_OUT156_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT157 = LC_HIGH_BIT_POS_PROBE_OUT156 + C_PROBE_OUT157_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT158 = LC_HIGH_BIT_POS_PROBE_OUT157 + C_PROBE_OUT158_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT159 = LC_HIGH_BIT_POS_PROBE_OUT158 + C_PROBE_OUT159_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT160 = LC_HIGH_BIT_POS_PROBE_OUT159 + C_PROBE_OUT160_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT161 = LC_HIGH_BIT_POS_PROBE_OUT160 + C_PROBE_OUT161_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT162 = LC_HIGH_BIT_POS_PROBE_OUT161 + C_PROBE_OUT162_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT163 = LC_HIGH_BIT_POS_PROBE_OUT162 + C_PROBE_OUT163_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT164 = LC_HIGH_BIT_POS_PROBE_OUT163 + C_PROBE_OUT164_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT165 = LC_HIGH_BIT_POS_PROBE_OUT164 + C_PROBE_OUT165_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT166 = LC_HIGH_BIT_POS_PROBE_OUT165 + C_PROBE_OUT166_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT167 = LC_HIGH_BIT_POS_PROBE_OUT166 + C_PROBE_OUT167_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT168 = LC_HIGH_BIT_POS_PROBE_OUT167 + C_PROBE_OUT168_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT169 = LC_HIGH_BIT_POS_PROBE_OUT168 + C_PROBE_OUT169_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT170 = LC_HIGH_BIT_POS_PROBE_OUT169 + C_PROBE_OUT170_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT171 = LC_HIGH_BIT_POS_PROBE_OUT170 + C_PROBE_OUT171_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT172 = LC_HIGH_BIT_POS_PROBE_OUT171 + C_PROBE_OUT172_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT173 = LC_HIGH_BIT_POS_PROBE_OUT172 + C_PROBE_OUT173_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT174 = LC_HIGH_BIT_POS_PROBE_OUT173 + C_PROBE_OUT174_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT175 = LC_HIGH_BIT_POS_PROBE_OUT174 + C_PROBE_OUT175_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT176 = LC_HIGH_BIT_POS_PROBE_OUT175 + C_PROBE_OUT176_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT177 = LC_HIGH_BIT_POS_PROBE_OUT176 + C_PROBE_OUT177_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT178 = LC_HIGH_BIT_POS_PROBE_OUT177 + C_PROBE_OUT178_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT179 = LC_HIGH_BIT_POS_PROBE_OUT178 + C_PROBE_OUT179_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT180 = LC_HIGH_BIT_POS_PROBE_OUT179 + C_PROBE_OUT180_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT181 = LC_HIGH_BIT_POS_PROBE_OUT180 + C_PROBE_OUT181_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT182 = LC_HIGH_BIT_POS_PROBE_OUT181 + C_PROBE_OUT182_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT183 = LC_HIGH_BIT_POS_PROBE_OUT182 + C_PROBE_OUT183_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT184 = LC_HIGH_BIT_POS_PROBE_OUT183 + C_PROBE_OUT184_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT185 = LC_HIGH_BIT_POS_PROBE_OUT184 + C_PROBE_OUT185_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT186 = LC_HIGH_BIT_POS_PROBE_OUT185 + C_PROBE_OUT186_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT187 = LC_HIGH_BIT_POS_PROBE_OUT186 + C_PROBE_OUT187_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT188 = LC_HIGH_BIT_POS_PROBE_OUT187 + C_PROBE_OUT188_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT189 = LC_HIGH_BIT_POS_PROBE_OUT188 + C_PROBE_OUT189_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT190 = LC_HIGH_BIT_POS_PROBE_OUT189 + C_PROBE_OUT190_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT191 = LC_HIGH_BIT_POS_PROBE_OUT190 + C_PROBE_OUT191_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT192 = LC_HIGH_BIT_POS_PROBE_OUT191 + C_PROBE_OUT192_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT193 = LC_HIGH_BIT_POS_PROBE_OUT192 + C_PROBE_OUT193_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT194 = LC_HIGH_BIT_POS_PROBE_OUT193 + C_PROBE_OUT194_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT195 = LC_HIGH_BIT_POS_PROBE_OUT194 + C_PROBE_OUT195_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT196 = LC_HIGH_BIT_POS_PROBE_OUT195 + C_PROBE_OUT196_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT197 = LC_HIGH_BIT_POS_PROBE_OUT196 + C_PROBE_OUT197_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT198 = LC_HIGH_BIT_POS_PROBE_OUT197 + C_PROBE_OUT198_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT199 = LC_HIGH_BIT_POS_PROBE_OUT198 + C_PROBE_OUT199_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT200 = LC_HIGH_BIT_POS_PROBE_OUT199 + C_PROBE_OUT200_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT201 = LC_HIGH_BIT_POS_PROBE_OUT200 + C_PROBE_OUT201_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT202 = LC_HIGH_BIT_POS_PROBE_OUT201 + C_PROBE_OUT202_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT203 = LC_HIGH_BIT_POS_PROBE_OUT202 + C_PROBE_OUT203_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT204 = LC_HIGH_BIT_POS_PROBE_OUT203 + C_PROBE_OUT204_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT205 = LC_HIGH_BIT_POS_PROBE_OUT204 + C_PROBE_OUT205_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT206 = LC_HIGH_BIT_POS_PROBE_OUT205 + C_PROBE_OUT206_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT207 = LC_HIGH_BIT_POS_PROBE_OUT206 + C_PROBE_OUT207_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT208 = LC_HIGH_BIT_POS_PROBE_OUT207 + C_PROBE_OUT208_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT209 = LC_HIGH_BIT_POS_PROBE_OUT208 + C_PROBE_OUT209_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT210 = LC_HIGH_BIT_POS_PROBE_OUT209 + C_PROBE_OUT210_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT211 = LC_HIGH_BIT_POS_PROBE_OUT210 + C_PROBE_OUT211_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT212 = LC_HIGH_BIT_POS_PROBE_OUT211 + C_PROBE_OUT212_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT213 = LC_HIGH_BIT_POS_PROBE_OUT212 + C_PROBE_OUT213_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT214 = LC_HIGH_BIT_POS_PROBE_OUT213 + C_PROBE_OUT214_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT215 = LC_HIGH_BIT_POS_PROBE_OUT214 + C_PROBE_OUT215_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT216 = LC_HIGH_BIT_POS_PROBE_OUT215 + C_PROBE_OUT216_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT217 = LC_HIGH_BIT_POS_PROBE_OUT216 + C_PROBE_OUT217_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT218 = LC_HIGH_BIT_POS_PROBE_OUT217 + C_PROBE_OUT218_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT219 = LC_HIGH_BIT_POS_PROBE_OUT218 + C_PROBE_OUT219_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT220 = LC_HIGH_BIT_POS_PROBE_OUT219 + C_PROBE_OUT220_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT221 = LC_HIGH_BIT_POS_PROBE_OUT220 + C_PROBE_OUT221_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT222 = LC_HIGH_BIT_POS_PROBE_OUT221 + C_PROBE_OUT222_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT223 = LC_HIGH_BIT_POS_PROBE_OUT222 + C_PROBE_OUT223_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT224 = LC_HIGH_BIT_POS_PROBE_OUT223 + C_PROBE_OUT224_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT225 = LC_HIGH_BIT_POS_PROBE_OUT224 + C_PROBE_OUT225_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT226 = LC_HIGH_BIT_POS_PROBE_OUT225 + C_PROBE_OUT226_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT227 = LC_HIGH_BIT_POS_PROBE_OUT226 + C_PROBE_OUT227_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT228 = LC_HIGH_BIT_POS_PROBE_OUT227 + C_PROBE_OUT228_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT229 = LC_HIGH_BIT_POS_PROBE_OUT228 + C_PROBE_OUT229_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT230 = LC_HIGH_BIT_POS_PROBE_OUT229 + C_PROBE_OUT230_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT231 = LC_HIGH_BIT_POS_PROBE_OUT230 + C_PROBE_OUT231_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT232 = LC_HIGH_BIT_POS_PROBE_OUT231 + C_PROBE_OUT232_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT233 = LC_HIGH_BIT_POS_PROBE_OUT232 + C_PROBE_OUT233_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT234 = LC_HIGH_BIT_POS_PROBE_OUT233 + C_PROBE_OUT234_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT235 = LC_HIGH_BIT_POS_PROBE_OUT234 + C_PROBE_OUT235_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT236 = LC_HIGH_BIT_POS_PROBE_OUT235 + C_PROBE_OUT236_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT237 = LC_HIGH_BIT_POS_PROBE_OUT236 + C_PROBE_OUT237_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT238 = LC_HIGH_BIT_POS_PROBE_OUT237 + C_PROBE_OUT238_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT239 = LC_HIGH_BIT_POS_PROBE_OUT238 + C_PROBE_OUT239_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT240 = LC_HIGH_BIT_POS_PROBE_OUT239 + C_PROBE_OUT240_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT241 = LC_HIGH_BIT_POS_PROBE_OUT240 + C_PROBE_OUT241_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT242 = LC_HIGH_BIT_POS_PROBE_OUT241 + C_PROBE_OUT242_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT243 = LC_HIGH_BIT_POS_PROBE_OUT242 + C_PROBE_OUT243_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT244 = LC_HIGH_BIT_POS_PROBE_OUT243 + C_PROBE_OUT244_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT245 = LC_HIGH_BIT_POS_PROBE_OUT244 + C_PROBE_OUT245_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT246 = LC_HIGH_BIT_POS_PROBE_OUT245 + C_PROBE_OUT246_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT247 = LC_HIGH_BIT_POS_PROBE_OUT246 + C_PROBE_OUT247_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT248 = LC_HIGH_BIT_POS_PROBE_OUT247 + C_PROBE_OUT248_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT249 = LC_HIGH_BIT_POS_PROBE_OUT248 + C_PROBE_OUT249_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT250 = LC_HIGH_BIT_POS_PROBE_OUT249 + C_PROBE_OUT250_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT251 = LC_HIGH_BIT_POS_PROBE_OUT250 + C_PROBE_OUT251_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT252 = LC_HIGH_BIT_POS_PROBE_OUT251 + C_PROBE_OUT252_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT253 = LC_HIGH_BIT_POS_PROBE_OUT252 + C_PROBE_OUT253_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT254 = LC_HIGH_BIT_POS_PROBE_OUT253 + C_PROBE_OUT254_WIDTH;
  localparam [15:0]LC_HIGH_BIT_POS_PROBE_OUT255 = LC_HIGH_BIT_POS_PROBE_OUT254 + C_PROBE_OUT255_WIDTH;
    
  localparam [4095:0]LC_PROBE_OUT_HIGH_BIT_POS_STRING = {
    LC_HIGH_BIT_POS_PROBE_OUT255, LC_HIGH_BIT_POS_PROBE_OUT254, 
    LC_HIGH_BIT_POS_PROBE_OUT253, LC_HIGH_BIT_POS_PROBE_OUT252, 
    LC_HIGH_BIT_POS_PROBE_OUT251, LC_HIGH_BIT_POS_PROBE_OUT250, 
    LC_HIGH_BIT_POS_PROBE_OUT249, LC_HIGH_BIT_POS_PROBE_OUT248, 
    LC_HIGH_BIT_POS_PROBE_OUT247, LC_HIGH_BIT_POS_PROBE_OUT246, 
    LC_HIGH_BIT_POS_PROBE_OUT245, LC_HIGH_BIT_POS_PROBE_OUT244, 
    LC_HIGH_BIT_POS_PROBE_OUT243, LC_HIGH_BIT_POS_PROBE_OUT242, 
    LC_HIGH_BIT_POS_PROBE_OUT241, LC_HIGH_BIT_POS_PROBE_OUT240, 
    LC_HIGH_BIT_POS_PROBE_OUT239, LC_HIGH_BIT_POS_PROBE_OUT238, 
    LC_HIGH_BIT_POS_PROBE_OUT237, LC_HIGH_BIT_POS_PROBE_OUT236, 
    LC_HIGH_BIT_POS_PROBE_OUT235, LC_HIGH_BIT_POS_PROBE_OUT234, 
    LC_HIGH_BIT_POS_PROBE_OUT233, LC_HIGH_BIT_POS_PROBE_OUT232, 
    LC_HIGH_BIT_POS_PROBE_OUT231, LC_HIGH_BIT_POS_PROBE_OUT230, 
    LC_HIGH_BIT_POS_PROBE_OUT229, LC_HIGH_BIT_POS_PROBE_OUT228, 
    LC_HIGH_BIT_POS_PROBE_OUT227, LC_HIGH_BIT_POS_PROBE_OUT226, 
    LC_HIGH_BIT_POS_PROBE_OUT225, LC_HIGH_BIT_POS_PROBE_OUT224, 
    LC_HIGH_BIT_POS_PROBE_OUT223, LC_HIGH_BIT_POS_PROBE_OUT222, 
    LC_HIGH_BIT_POS_PROBE_OUT221, LC_HIGH_BIT_POS_PROBE_OUT220, 
    LC_HIGH_BIT_POS_PROBE_OUT219, LC_HIGH_BIT_POS_PROBE_OUT218, 
    LC_HIGH_BIT_POS_PROBE_OUT217, LC_HIGH_BIT_POS_PROBE_OUT216, 
    LC_HIGH_BIT_POS_PROBE_OUT215, LC_HIGH_BIT_POS_PROBE_OUT214, 
    LC_HIGH_BIT_POS_PROBE_OUT213, LC_HIGH_BIT_POS_PROBE_OUT212, 
    LC_HIGH_BIT_POS_PROBE_OUT211, LC_HIGH_BIT_POS_PROBE_OUT210, 
    LC_HIGH_BIT_POS_PROBE_OUT209, LC_HIGH_BIT_POS_PROBE_OUT208, 
    LC_HIGH_BIT_POS_PROBE_OUT207, LC_HIGH_BIT_POS_PROBE_OUT206, 
    LC_HIGH_BIT_POS_PROBE_OUT205, LC_HIGH_BIT_POS_PROBE_OUT204, 
    LC_HIGH_BIT_POS_PROBE_OUT203, LC_HIGH_BIT_POS_PROBE_OUT202, 
    LC_HIGH_BIT_POS_PROBE_OUT201, LC_HIGH_BIT_POS_PROBE_OUT200, 
    LC_HIGH_BIT_POS_PROBE_OUT199, LC_HIGH_BIT_POS_PROBE_OUT198, 
    LC_HIGH_BIT_POS_PROBE_OUT197, LC_HIGH_BIT_POS_PROBE_OUT196, 
    LC_HIGH_BIT_POS_PROBE_OUT195, LC_HIGH_BIT_POS_PROBE_OUT194, 
    LC_HIGH_BIT_POS_PROBE_OUT193, LC_HIGH_BIT_POS_PROBE_OUT192, 
    LC_HIGH_BIT_POS_PROBE_OUT191, LC_HIGH_BIT_POS_PROBE_OUT190, 
    LC_HIGH_BIT_POS_PROBE_OUT189, LC_HIGH_BIT_POS_PROBE_OUT188, 
    LC_HIGH_BIT_POS_PROBE_OUT187, LC_HIGH_BIT_POS_PROBE_OUT186, 
    LC_HIGH_BIT_POS_PROBE_OUT185, LC_HIGH_BIT_POS_PROBE_OUT184, 
    LC_HIGH_BIT_POS_PROBE_OUT183, LC_HIGH_BIT_POS_PROBE_OUT182, 
    LC_HIGH_BIT_POS_PROBE_OUT181, LC_HIGH_BIT_POS_PROBE_OUT180, 
    LC_HIGH_BIT_POS_PROBE_OUT179, LC_HIGH_BIT_POS_PROBE_OUT178, 
    LC_HIGH_BIT_POS_PROBE_OUT177, LC_HIGH_BIT_POS_PROBE_OUT176, 
    LC_HIGH_BIT_POS_PROBE_OUT175, LC_HIGH_BIT_POS_PROBE_OUT174, 
    LC_HIGH_BIT_POS_PROBE_OUT173, LC_HIGH_BIT_POS_PROBE_OUT172, 
    LC_HIGH_BIT_POS_PROBE_OUT171, LC_HIGH_BIT_POS_PROBE_OUT170, 
    LC_HIGH_BIT_POS_PROBE_OUT169, LC_HIGH_BIT_POS_PROBE_OUT168, 
    LC_HIGH_BIT_POS_PROBE_OUT167, LC_HIGH_BIT_POS_PROBE_OUT166, 
    LC_HIGH_BIT_POS_PROBE_OUT165, LC_HIGH_BIT_POS_PROBE_OUT164, 
    LC_HIGH_BIT_POS_PROBE_OUT163, LC_HIGH_BIT_POS_PROBE_OUT162, 
    LC_HIGH_BIT_POS_PROBE_OUT161, LC_HIGH_BIT_POS_PROBE_OUT160, 
    LC_HIGH_BIT_POS_PROBE_OUT159, LC_HIGH_BIT_POS_PROBE_OUT158, 
    LC_HIGH_BIT_POS_PROBE_OUT157, LC_HIGH_BIT_POS_PROBE_OUT156, 
    LC_HIGH_BIT_POS_PROBE_OUT155, LC_HIGH_BIT_POS_PROBE_OUT154, 
    LC_HIGH_BIT_POS_PROBE_OUT153, LC_HIGH_BIT_POS_PROBE_OUT152, 
    LC_HIGH_BIT_POS_PROBE_OUT151, LC_HIGH_BIT_POS_PROBE_OUT150, 
    LC_HIGH_BIT_POS_PROBE_OUT149, LC_HIGH_BIT_POS_PROBE_OUT148, 
    LC_HIGH_BIT_POS_PROBE_OUT147, LC_HIGH_BIT_POS_PROBE_OUT146, 
    LC_HIGH_BIT_POS_PROBE_OUT145, LC_HIGH_BIT_POS_PROBE_OUT144, 
    LC_HIGH_BIT_POS_PROBE_OUT143, LC_HIGH_BIT_POS_PROBE_OUT142, 
    LC_HIGH_BIT_POS_PROBE_OUT141, LC_HIGH_BIT_POS_PROBE_OUT140, 
    LC_HIGH_BIT_POS_PROBE_OUT139, LC_HIGH_BIT_POS_PROBE_OUT138, 
    LC_HIGH_BIT_POS_PROBE_OUT137, LC_HIGH_BIT_POS_PROBE_OUT136, 
    LC_HIGH_BIT_POS_PROBE_OUT135, LC_HIGH_BIT_POS_PROBE_OUT134, 
    LC_HIGH_BIT_POS_PROBE_OUT133, LC_HIGH_BIT_POS_PROBE_OUT132, 
    LC_HIGH_BIT_POS_PROBE_OUT131, LC_HIGH_BIT_POS_PROBE_OUT130, 
    LC_HIGH_BIT_POS_PROBE_OUT129, LC_HIGH_BIT_POS_PROBE_OUT128, 
    LC_HIGH_BIT_POS_PROBE_OUT127, LC_HIGH_BIT_POS_PROBE_OUT126, 
    LC_HIGH_BIT_POS_PROBE_OUT125, LC_HIGH_BIT_POS_PROBE_OUT124, 
    LC_HIGH_BIT_POS_PROBE_OUT123, LC_HIGH_BIT_POS_PROBE_OUT122, 
    LC_HIGH_BIT_POS_PROBE_OUT121, LC_HIGH_BIT_POS_PROBE_OUT120, 
    LC_HIGH_BIT_POS_PROBE_OUT119, LC_HIGH_BIT_POS_PROBE_OUT118, 
    LC_HIGH_BIT_POS_PROBE_OUT117, LC_HIGH_BIT_POS_PROBE_OUT116, 
    LC_HIGH_BIT_POS_PROBE_OUT115, LC_HIGH_BIT_POS_PROBE_OUT114, 
    LC_HIGH_BIT_POS_PROBE_OUT113, LC_HIGH_BIT_POS_PROBE_OUT112, 
    LC_HIGH_BIT_POS_PROBE_OUT111, LC_HIGH_BIT_POS_PROBE_OUT110, 
    LC_HIGH_BIT_POS_PROBE_OUT109, LC_HIGH_BIT_POS_PROBE_OUT108, 
    LC_HIGH_BIT_POS_PROBE_OUT107, LC_HIGH_BIT_POS_PROBE_OUT106, 
    LC_HIGH_BIT_POS_PROBE_OUT105, LC_HIGH_BIT_POS_PROBE_OUT104, 
    LC_HIGH_BIT_POS_PROBE_OUT103, LC_HIGH_BIT_POS_PROBE_OUT102, 
    LC_HIGH_BIT_POS_PROBE_OUT101, LC_HIGH_BIT_POS_PROBE_OUT100, 
    LC_HIGH_BIT_POS_PROBE_OUT99 , LC_HIGH_BIT_POS_PROBE_OUT98 , 
    LC_HIGH_BIT_POS_PROBE_OUT97 , LC_HIGH_BIT_POS_PROBE_OUT96 , 
    LC_HIGH_BIT_POS_PROBE_OUT95 , LC_HIGH_BIT_POS_PROBE_OUT94 , 
    LC_HIGH_BIT_POS_PROBE_OUT93 , LC_HIGH_BIT_POS_PROBE_OUT92 , 
    LC_HIGH_BIT_POS_PROBE_OUT91 , LC_HIGH_BIT_POS_PROBE_OUT90 , 
    LC_HIGH_BIT_POS_PROBE_OUT89 , LC_HIGH_BIT_POS_PROBE_OUT88 , 
    LC_HIGH_BIT_POS_PROBE_OUT87 , LC_HIGH_BIT_POS_PROBE_OUT86 , 
    LC_HIGH_BIT_POS_PROBE_OUT85 , LC_HIGH_BIT_POS_PROBE_OUT84 , 
    LC_HIGH_BIT_POS_PROBE_OUT83 , LC_HIGH_BIT_POS_PROBE_OUT82 , 
    LC_HIGH_BIT_POS_PROBE_OUT81 , LC_HIGH_BIT_POS_PROBE_OUT80 , 
    LC_HIGH_BIT_POS_PROBE_OUT79 , LC_HIGH_BIT_POS_PROBE_OUT78 , 
    LC_HIGH_BIT_POS_PROBE_OUT77 , LC_HIGH_BIT_POS_PROBE_OUT76 , 
    LC_HIGH_BIT_POS_PROBE_OUT75 , LC_HIGH_BIT_POS_PROBE_OUT74 , 
    LC_HIGH_BIT_POS_PROBE_OUT73 , LC_HIGH_BIT_POS_PROBE_OUT72 , 
    LC_HIGH_BIT_POS_PROBE_OUT71 , LC_HIGH_BIT_POS_PROBE_OUT70 , 
    LC_HIGH_BIT_POS_PROBE_OUT69 , LC_HIGH_BIT_POS_PROBE_OUT68 , 
    LC_HIGH_BIT_POS_PROBE_OUT67 , LC_HIGH_BIT_POS_PROBE_OUT66 , 
    LC_HIGH_BIT_POS_PROBE_OUT65 , LC_HIGH_BIT_POS_PROBE_OUT64 , 
    LC_HIGH_BIT_POS_PROBE_OUT63 , LC_HIGH_BIT_POS_PROBE_OUT62 , 
    LC_HIGH_BIT_POS_PROBE_OUT61 , LC_HIGH_BIT_POS_PROBE_OUT60 , 
    LC_HIGH_BIT_POS_PROBE_OUT59 , LC_HIGH_BIT_POS_PROBE_OUT58 , 
    LC_HIGH_BIT_POS_PROBE_OUT57 , LC_HIGH_BIT_POS_PROBE_OUT56 , 
    LC_HIGH_BIT_POS_PROBE_OUT55 , LC_HIGH_BIT_POS_PROBE_OUT54 , 
    LC_HIGH_BIT_POS_PROBE_OUT53 , LC_HIGH_BIT_POS_PROBE_OUT52 , 
    LC_HIGH_BIT_POS_PROBE_OUT51 , LC_HIGH_BIT_POS_PROBE_OUT50 , 
    LC_HIGH_BIT_POS_PROBE_OUT49 , LC_HIGH_BIT_POS_PROBE_OUT48 , 
    LC_HIGH_BIT_POS_PROBE_OUT47 , LC_HIGH_BIT_POS_PROBE_OUT46 , 
    LC_HIGH_BIT_POS_PROBE_OUT45 , LC_HIGH_BIT_POS_PROBE_OUT44 , 
    LC_HIGH_BIT_POS_PROBE_OUT43 , LC_HIGH_BIT_POS_PROBE_OUT42 , 
    LC_HIGH_BIT_POS_PROBE_OUT41 , LC_HIGH_BIT_POS_PROBE_OUT40 , 
    LC_HIGH_BIT_POS_PROBE_OUT39 , LC_HIGH_BIT_POS_PROBE_OUT38 , 
    LC_HIGH_BIT_POS_PROBE_OUT37 , LC_HIGH_BIT_POS_PROBE_OUT36 , 
    LC_HIGH_BIT_POS_PROBE_OUT35 , LC_HIGH_BIT_POS_PROBE_OUT34 , 
    LC_HIGH_BIT_POS_PROBE_OUT33 , LC_HIGH_BIT_POS_PROBE_OUT32 , 
    LC_HIGH_BIT_POS_PROBE_OUT31 , LC_HIGH_BIT_POS_PROBE_OUT30 , 
    LC_HIGH_BIT_POS_PROBE_OUT29 , LC_HIGH_BIT_POS_PROBE_OUT28 , 
    LC_HIGH_BIT_POS_PROBE_OUT27 , LC_HIGH_BIT_POS_PROBE_OUT26 , 
    LC_HIGH_BIT_POS_PROBE_OUT25 , LC_HIGH_BIT_POS_PROBE_OUT24 , 
    LC_HIGH_BIT_POS_PROBE_OUT23 , LC_HIGH_BIT_POS_PROBE_OUT22 , 
    LC_HIGH_BIT_POS_PROBE_OUT21 , LC_HIGH_BIT_POS_PROBE_OUT20 , 
    LC_HIGH_BIT_POS_PROBE_OUT19 , LC_HIGH_BIT_POS_PROBE_OUT18 , 
    LC_HIGH_BIT_POS_PROBE_OUT17 , LC_HIGH_BIT_POS_PROBE_OUT16 , 
    LC_HIGH_BIT_POS_PROBE_OUT15 , LC_HIGH_BIT_POS_PROBE_OUT14 , 
    LC_HIGH_BIT_POS_PROBE_OUT13 , LC_HIGH_BIT_POS_PROBE_OUT12 , 
    LC_HIGH_BIT_POS_PROBE_OUT11 , LC_HIGH_BIT_POS_PROBE_OUT10 , 
    LC_HIGH_BIT_POS_PROBE_OUT9  , LC_HIGH_BIT_POS_PROBE_OUT8  , 
    LC_HIGH_BIT_POS_PROBE_OUT7  , LC_HIGH_BIT_POS_PROBE_OUT6  , 
    LC_HIGH_BIT_POS_PROBE_OUT5  , LC_HIGH_BIT_POS_PROBE_OUT4  , 
    LC_HIGH_BIT_POS_PROBE_OUT3  , LC_HIGH_BIT_POS_PROBE_OUT2  , 
    LC_HIGH_BIT_POS_PROBE_OUT1  , LC_HIGH_BIT_POS_PROBE_OUT0
  };

  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT0   = 0                               ;	        
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT1   = LC_HIGH_BIT_POS_PROBE_OUT0   + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT2   = LC_HIGH_BIT_POS_PROBE_OUT1   + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT3   = LC_HIGH_BIT_POS_PROBE_OUT2   + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT4   = LC_HIGH_BIT_POS_PROBE_OUT3   + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT5   = LC_HIGH_BIT_POS_PROBE_OUT4   + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT6   = LC_HIGH_BIT_POS_PROBE_OUT5   + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT7   = LC_HIGH_BIT_POS_PROBE_OUT6   + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT8   = LC_HIGH_BIT_POS_PROBE_OUT7   + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT9   = LC_HIGH_BIT_POS_PROBE_OUT8   + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT10  = LC_HIGH_BIT_POS_PROBE_OUT9   + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT11  = LC_HIGH_BIT_POS_PROBE_OUT10  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT12  = LC_HIGH_BIT_POS_PROBE_OUT11  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT13  = LC_HIGH_BIT_POS_PROBE_OUT12  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT14  = LC_HIGH_BIT_POS_PROBE_OUT13  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT15  = LC_HIGH_BIT_POS_PROBE_OUT14  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT16  = LC_HIGH_BIT_POS_PROBE_OUT15  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT17  = LC_HIGH_BIT_POS_PROBE_OUT16  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT18  = LC_HIGH_BIT_POS_PROBE_OUT17  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT19  = LC_HIGH_BIT_POS_PROBE_OUT18  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT20  = LC_HIGH_BIT_POS_PROBE_OUT19  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT21  = LC_HIGH_BIT_POS_PROBE_OUT20  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT22  = LC_HIGH_BIT_POS_PROBE_OUT21  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT23  = LC_HIGH_BIT_POS_PROBE_OUT22  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT24  = LC_HIGH_BIT_POS_PROBE_OUT23  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT25  = LC_HIGH_BIT_POS_PROBE_OUT24  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT26  = LC_HIGH_BIT_POS_PROBE_OUT25  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT27  = LC_HIGH_BIT_POS_PROBE_OUT26  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT28  = LC_HIGH_BIT_POS_PROBE_OUT27  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT29  = LC_HIGH_BIT_POS_PROBE_OUT28  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT30  = LC_HIGH_BIT_POS_PROBE_OUT29  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT31  = LC_HIGH_BIT_POS_PROBE_OUT30  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT32  = LC_HIGH_BIT_POS_PROBE_OUT31  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT33  = LC_HIGH_BIT_POS_PROBE_OUT32  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT34  = LC_HIGH_BIT_POS_PROBE_OUT33  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT35  = LC_HIGH_BIT_POS_PROBE_OUT34  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT36  = LC_HIGH_BIT_POS_PROBE_OUT35  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT37  = LC_HIGH_BIT_POS_PROBE_OUT36  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT38  = LC_HIGH_BIT_POS_PROBE_OUT37  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT39  = LC_HIGH_BIT_POS_PROBE_OUT38  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT40  = LC_HIGH_BIT_POS_PROBE_OUT39  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT41  = LC_HIGH_BIT_POS_PROBE_OUT40  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT42  = LC_HIGH_BIT_POS_PROBE_OUT41  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT43  = LC_HIGH_BIT_POS_PROBE_OUT42  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT44  = LC_HIGH_BIT_POS_PROBE_OUT43  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT45  = LC_HIGH_BIT_POS_PROBE_OUT44  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT46  = LC_HIGH_BIT_POS_PROBE_OUT45  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT47  = LC_HIGH_BIT_POS_PROBE_OUT46  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT48  = LC_HIGH_BIT_POS_PROBE_OUT47  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT49  = LC_HIGH_BIT_POS_PROBE_OUT48  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT50  = LC_HIGH_BIT_POS_PROBE_OUT49  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT51  = LC_HIGH_BIT_POS_PROBE_OUT50  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT52  = LC_HIGH_BIT_POS_PROBE_OUT51  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT53  = LC_HIGH_BIT_POS_PROBE_OUT52  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT54  = LC_HIGH_BIT_POS_PROBE_OUT53  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT55  = LC_HIGH_BIT_POS_PROBE_OUT54  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT56  = LC_HIGH_BIT_POS_PROBE_OUT55  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT57  = LC_HIGH_BIT_POS_PROBE_OUT56  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT58  = LC_HIGH_BIT_POS_PROBE_OUT57  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT59  = LC_HIGH_BIT_POS_PROBE_OUT58  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT60  = LC_HIGH_BIT_POS_PROBE_OUT59  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT61  = LC_HIGH_BIT_POS_PROBE_OUT60  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT62  = LC_HIGH_BIT_POS_PROBE_OUT61  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT63  = LC_HIGH_BIT_POS_PROBE_OUT62  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT64  = LC_HIGH_BIT_POS_PROBE_OUT63  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT65  = LC_HIGH_BIT_POS_PROBE_OUT64  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT66  = LC_HIGH_BIT_POS_PROBE_OUT65  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT67  = LC_HIGH_BIT_POS_PROBE_OUT66  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT68  = LC_HIGH_BIT_POS_PROBE_OUT67  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT69  = LC_HIGH_BIT_POS_PROBE_OUT68  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT70  = LC_HIGH_BIT_POS_PROBE_OUT69  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT71  = LC_HIGH_BIT_POS_PROBE_OUT70  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT72  = LC_HIGH_BIT_POS_PROBE_OUT71  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT73  = LC_HIGH_BIT_POS_PROBE_OUT72  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT74  = LC_HIGH_BIT_POS_PROBE_OUT73  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT75  = LC_HIGH_BIT_POS_PROBE_OUT74  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT76  = LC_HIGH_BIT_POS_PROBE_OUT75  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT77  = LC_HIGH_BIT_POS_PROBE_OUT76  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT78  = LC_HIGH_BIT_POS_PROBE_OUT77  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT79  = LC_HIGH_BIT_POS_PROBE_OUT78  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT80  = LC_HIGH_BIT_POS_PROBE_OUT79  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT81  = LC_HIGH_BIT_POS_PROBE_OUT80  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT82  = LC_HIGH_BIT_POS_PROBE_OUT81  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT83  = LC_HIGH_BIT_POS_PROBE_OUT82  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT84  = LC_HIGH_BIT_POS_PROBE_OUT83  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT85  = LC_HIGH_BIT_POS_PROBE_OUT84  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT86  = LC_HIGH_BIT_POS_PROBE_OUT85  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT87  = LC_HIGH_BIT_POS_PROBE_OUT86  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT88  = LC_HIGH_BIT_POS_PROBE_OUT87  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT89  = LC_HIGH_BIT_POS_PROBE_OUT88  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT90  = LC_HIGH_BIT_POS_PROBE_OUT89  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT91  = LC_HIGH_BIT_POS_PROBE_OUT90  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT92  = LC_HIGH_BIT_POS_PROBE_OUT91  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT93  = LC_HIGH_BIT_POS_PROBE_OUT92  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT94  = LC_HIGH_BIT_POS_PROBE_OUT93  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT95  = LC_HIGH_BIT_POS_PROBE_OUT94  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT96  = LC_HIGH_BIT_POS_PROBE_OUT95  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT97  = LC_HIGH_BIT_POS_PROBE_OUT96  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT98  = LC_HIGH_BIT_POS_PROBE_OUT97  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT99  = LC_HIGH_BIT_POS_PROBE_OUT98  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT100 = LC_HIGH_BIT_POS_PROBE_OUT99  + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT101 = LC_HIGH_BIT_POS_PROBE_OUT100 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT102 = LC_HIGH_BIT_POS_PROBE_OUT101 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT103 = LC_HIGH_BIT_POS_PROBE_OUT102 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT104 = LC_HIGH_BIT_POS_PROBE_OUT103 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT105 = LC_HIGH_BIT_POS_PROBE_OUT104 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT106 = LC_HIGH_BIT_POS_PROBE_OUT105 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT107 = LC_HIGH_BIT_POS_PROBE_OUT106 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT108 = LC_HIGH_BIT_POS_PROBE_OUT107 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT109 = LC_HIGH_BIT_POS_PROBE_OUT108 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT110 = LC_HIGH_BIT_POS_PROBE_OUT109 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT111 = LC_HIGH_BIT_POS_PROBE_OUT110 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT112 = LC_HIGH_BIT_POS_PROBE_OUT111 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT113 = LC_HIGH_BIT_POS_PROBE_OUT112 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT114 = LC_HIGH_BIT_POS_PROBE_OUT113 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT115 = LC_HIGH_BIT_POS_PROBE_OUT114 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT116 = LC_HIGH_BIT_POS_PROBE_OUT115 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT117 = LC_HIGH_BIT_POS_PROBE_OUT116 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT118 = LC_HIGH_BIT_POS_PROBE_OUT117 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT119 = LC_HIGH_BIT_POS_PROBE_OUT118 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT120 = LC_HIGH_BIT_POS_PROBE_OUT119 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT121 = LC_HIGH_BIT_POS_PROBE_OUT120 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT122 = LC_HIGH_BIT_POS_PROBE_OUT121 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT123 = LC_HIGH_BIT_POS_PROBE_OUT122 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT124 = LC_HIGH_BIT_POS_PROBE_OUT123 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT125 = LC_HIGH_BIT_POS_PROBE_OUT124 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT126 = LC_HIGH_BIT_POS_PROBE_OUT125 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT127 = LC_HIGH_BIT_POS_PROBE_OUT126 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT128 = LC_HIGH_BIT_POS_PROBE_OUT127 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT129 = LC_HIGH_BIT_POS_PROBE_OUT128 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT130 = LC_HIGH_BIT_POS_PROBE_OUT129 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT131 = LC_HIGH_BIT_POS_PROBE_OUT130 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT132 = LC_HIGH_BIT_POS_PROBE_OUT131 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT133 = LC_HIGH_BIT_POS_PROBE_OUT132 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT134 = LC_HIGH_BIT_POS_PROBE_OUT133 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT135 = LC_HIGH_BIT_POS_PROBE_OUT134 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT136 = LC_HIGH_BIT_POS_PROBE_OUT135 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT137 = LC_HIGH_BIT_POS_PROBE_OUT136 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT138 = LC_HIGH_BIT_POS_PROBE_OUT137 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT139 = LC_HIGH_BIT_POS_PROBE_OUT138 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT140 = LC_HIGH_BIT_POS_PROBE_OUT139 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT141 = LC_HIGH_BIT_POS_PROBE_OUT140 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT142 = LC_HIGH_BIT_POS_PROBE_OUT141 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT143 = LC_HIGH_BIT_POS_PROBE_OUT142 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT144 = LC_HIGH_BIT_POS_PROBE_OUT143 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT145 = LC_HIGH_BIT_POS_PROBE_OUT144 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT146 = LC_HIGH_BIT_POS_PROBE_OUT145 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT147 = LC_HIGH_BIT_POS_PROBE_OUT146 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT148 = LC_HIGH_BIT_POS_PROBE_OUT147 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT149 = LC_HIGH_BIT_POS_PROBE_OUT148 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT150 = LC_HIGH_BIT_POS_PROBE_OUT149 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT151 = LC_HIGH_BIT_POS_PROBE_OUT150 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT152 = LC_HIGH_BIT_POS_PROBE_OUT151 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT153 = LC_HIGH_BIT_POS_PROBE_OUT152 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT154 = LC_HIGH_BIT_POS_PROBE_OUT153 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT155 = LC_HIGH_BIT_POS_PROBE_OUT154 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT156 = LC_HIGH_BIT_POS_PROBE_OUT155 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT157 = LC_HIGH_BIT_POS_PROBE_OUT156 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT158 = LC_HIGH_BIT_POS_PROBE_OUT157 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT159 = LC_HIGH_BIT_POS_PROBE_OUT158 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT160 = LC_HIGH_BIT_POS_PROBE_OUT159 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT161 = LC_HIGH_BIT_POS_PROBE_OUT160 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT162 = LC_HIGH_BIT_POS_PROBE_OUT161 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT163 = LC_HIGH_BIT_POS_PROBE_OUT162 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT164 = LC_HIGH_BIT_POS_PROBE_OUT163 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT165 = LC_HIGH_BIT_POS_PROBE_OUT164 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT166 = LC_HIGH_BIT_POS_PROBE_OUT165 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT167 = LC_HIGH_BIT_POS_PROBE_OUT166 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT168 = LC_HIGH_BIT_POS_PROBE_OUT167 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT169 = LC_HIGH_BIT_POS_PROBE_OUT168 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT170 = LC_HIGH_BIT_POS_PROBE_OUT169 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT171 = LC_HIGH_BIT_POS_PROBE_OUT170 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT172 = LC_HIGH_BIT_POS_PROBE_OUT171 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT173 = LC_HIGH_BIT_POS_PROBE_OUT172 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT174 = LC_HIGH_BIT_POS_PROBE_OUT173 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT175 = LC_HIGH_BIT_POS_PROBE_OUT174 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT176 = LC_HIGH_BIT_POS_PROBE_OUT175 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT177 = LC_HIGH_BIT_POS_PROBE_OUT176 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT178 = LC_HIGH_BIT_POS_PROBE_OUT177 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT179 = LC_HIGH_BIT_POS_PROBE_OUT178 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT180 = LC_HIGH_BIT_POS_PROBE_OUT179 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT181 = LC_HIGH_BIT_POS_PROBE_OUT180 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT182 = LC_HIGH_BIT_POS_PROBE_OUT181 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT183 = LC_HIGH_BIT_POS_PROBE_OUT182 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT184 = LC_HIGH_BIT_POS_PROBE_OUT183 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT185 = LC_HIGH_BIT_POS_PROBE_OUT184 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT186 = LC_HIGH_BIT_POS_PROBE_OUT185 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT187 = LC_HIGH_BIT_POS_PROBE_OUT186 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT188 = LC_HIGH_BIT_POS_PROBE_OUT187 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT189 = LC_HIGH_BIT_POS_PROBE_OUT188 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT190 = LC_HIGH_BIT_POS_PROBE_OUT189 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT191 = LC_HIGH_BIT_POS_PROBE_OUT190 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT192 = LC_HIGH_BIT_POS_PROBE_OUT191 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT193 = LC_HIGH_BIT_POS_PROBE_OUT192 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT194 = LC_HIGH_BIT_POS_PROBE_OUT193 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT195 = LC_HIGH_BIT_POS_PROBE_OUT194 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT196 = LC_HIGH_BIT_POS_PROBE_OUT195 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT197 = LC_HIGH_BIT_POS_PROBE_OUT196 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT198 = LC_HIGH_BIT_POS_PROBE_OUT197 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT199 = LC_HIGH_BIT_POS_PROBE_OUT198 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT200 = LC_HIGH_BIT_POS_PROBE_OUT199 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT201 = LC_HIGH_BIT_POS_PROBE_OUT200 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT202 = LC_HIGH_BIT_POS_PROBE_OUT201 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT203 = LC_HIGH_BIT_POS_PROBE_OUT202 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT204 = LC_HIGH_BIT_POS_PROBE_OUT203 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT205 = LC_HIGH_BIT_POS_PROBE_OUT204 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT206 = LC_HIGH_BIT_POS_PROBE_OUT205 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT207 = LC_HIGH_BIT_POS_PROBE_OUT206 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT208 = LC_HIGH_BIT_POS_PROBE_OUT207 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT209 = LC_HIGH_BIT_POS_PROBE_OUT208 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT210 = LC_HIGH_BIT_POS_PROBE_OUT209 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT211 = LC_HIGH_BIT_POS_PROBE_OUT210 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT212 = LC_HIGH_BIT_POS_PROBE_OUT211 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT213 = LC_HIGH_BIT_POS_PROBE_OUT212 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT214 = LC_HIGH_BIT_POS_PROBE_OUT213 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT215 = LC_HIGH_BIT_POS_PROBE_OUT214 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT216 = LC_HIGH_BIT_POS_PROBE_OUT215 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT217 = LC_HIGH_BIT_POS_PROBE_OUT216 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT218 = LC_HIGH_BIT_POS_PROBE_OUT217 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT219 = LC_HIGH_BIT_POS_PROBE_OUT218 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT220 = LC_HIGH_BIT_POS_PROBE_OUT219 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT221 = LC_HIGH_BIT_POS_PROBE_OUT220 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT222 = LC_HIGH_BIT_POS_PROBE_OUT221 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT223 = LC_HIGH_BIT_POS_PROBE_OUT222 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT224 = LC_HIGH_BIT_POS_PROBE_OUT223 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT225 = LC_HIGH_BIT_POS_PROBE_OUT224 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT226 = LC_HIGH_BIT_POS_PROBE_OUT225 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT227 = LC_HIGH_BIT_POS_PROBE_OUT226 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT228 = LC_HIGH_BIT_POS_PROBE_OUT227 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT229 = LC_HIGH_BIT_POS_PROBE_OUT228 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT230 = LC_HIGH_BIT_POS_PROBE_OUT229 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT231 = LC_HIGH_BIT_POS_PROBE_OUT230 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT232 = LC_HIGH_BIT_POS_PROBE_OUT231 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT233 = LC_HIGH_BIT_POS_PROBE_OUT232 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT234 = LC_HIGH_BIT_POS_PROBE_OUT233 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT235 = LC_HIGH_BIT_POS_PROBE_OUT234 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT236 = LC_HIGH_BIT_POS_PROBE_OUT235 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT237 = LC_HIGH_BIT_POS_PROBE_OUT236 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT238 = LC_HIGH_BIT_POS_PROBE_OUT237 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT239 = LC_HIGH_BIT_POS_PROBE_OUT238 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT240 = LC_HIGH_BIT_POS_PROBE_OUT239 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT241 = LC_HIGH_BIT_POS_PROBE_OUT240 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT242 = LC_HIGH_BIT_POS_PROBE_OUT241 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT243 = LC_HIGH_BIT_POS_PROBE_OUT242 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT244 = LC_HIGH_BIT_POS_PROBE_OUT243 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT245 = LC_HIGH_BIT_POS_PROBE_OUT244 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT246 = LC_HIGH_BIT_POS_PROBE_OUT245 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT247 = LC_HIGH_BIT_POS_PROBE_OUT246 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT248 = LC_HIGH_BIT_POS_PROBE_OUT247 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT249 = LC_HIGH_BIT_POS_PROBE_OUT248 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT250 = LC_HIGH_BIT_POS_PROBE_OUT249 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT251 = LC_HIGH_BIT_POS_PROBE_OUT250 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT252 = LC_HIGH_BIT_POS_PROBE_OUT251 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT253 = LC_HIGH_BIT_POS_PROBE_OUT252 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT254 = LC_HIGH_BIT_POS_PROBE_OUT253 + 1;
  localparam [15:0]LC_LOW_BIT_POS_PROBE_OUT255 = LC_HIGH_BIT_POS_PROBE_OUT254 + 1;
    
  localparam [4095:0]LC_PROBE_OUT_LOW_BIT_POS_STRING = {
    LC_LOW_BIT_POS_PROBE_OUT255, LC_LOW_BIT_POS_PROBE_OUT254, 
    LC_LOW_BIT_POS_PROBE_OUT253, LC_LOW_BIT_POS_PROBE_OUT252, 
    LC_LOW_BIT_POS_PROBE_OUT251, LC_LOW_BIT_POS_PROBE_OUT250, 
    LC_LOW_BIT_POS_PROBE_OUT249, LC_LOW_BIT_POS_PROBE_OUT248, 
    LC_LOW_BIT_POS_PROBE_OUT247, LC_LOW_BIT_POS_PROBE_OUT246, 
    LC_LOW_BIT_POS_PROBE_OUT245, LC_LOW_BIT_POS_PROBE_OUT244, 
    LC_LOW_BIT_POS_PROBE_OUT243, LC_LOW_BIT_POS_PROBE_OUT242, 
    LC_LOW_BIT_POS_PROBE_OUT241, LC_LOW_BIT_POS_PROBE_OUT240, 
    LC_LOW_BIT_POS_PROBE_OUT239, LC_LOW_BIT_POS_PROBE_OUT238, 
    LC_LOW_BIT_POS_PROBE_OUT237, LC_LOW_BIT_POS_PROBE_OUT236, 
    LC_LOW_BIT_POS_PROBE_OUT235, LC_LOW_BIT_POS_PROBE_OUT234, 
    LC_LOW_BIT_POS_PROBE_OUT233, LC_LOW_BIT_POS_PROBE_OUT232, 
    LC_LOW_BIT_POS_PROBE_OUT231, LC_LOW_BIT_POS_PROBE_OUT230, 
    LC_LOW_BIT_POS_PROBE_OUT229, LC_LOW_BIT_POS_PROBE_OUT228, 
    LC_LOW_BIT_POS_PROBE_OUT227, LC_LOW_BIT_POS_PROBE_OUT226, 
    LC_LOW_BIT_POS_PROBE_OUT225, LC_LOW_BIT_POS_PROBE_OUT224, 
    LC_LOW_BIT_POS_PROBE_OUT223, LC_LOW_BIT_POS_PROBE_OUT222, 
    LC_LOW_BIT_POS_PROBE_OUT221, LC_LOW_BIT_POS_PROBE_OUT220, 
    LC_LOW_BIT_POS_PROBE_OUT219, LC_LOW_BIT_POS_PROBE_OUT218, 
    LC_LOW_BIT_POS_PROBE_OUT217, LC_LOW_BIT_POS_PROBE_OUT216, 
    LC_LOW_BIT_POS_PROBE_OUT215, LC_LOW_BIT_POS_PROBE_OUT214, 
    LC_LOW_BIT_POS_PROBE_OUT213, LC_LOW_BIT_POS_PROBE_OUT212, 
    LC_LOW_BIT_POS_PROBE_OUT211, LC_LOW_BIT_POS_PROBE_OUT210, 
    LC_LOW_BIT_POS_PROBE_OUT209, LC_LOW_BIT_POS_PROBE_OUT208, 
    LC_LOW_BIT_POS_PROBE_OUT207, LC_LOW_BIT_POS_PROBE_OUT206, 
    LC_LOW_BIT_POS_PROBE_OUT205, LC_LOW_BIT_POS_PROBE_OUT204, 
    LC_LOW_BIT_POS_PROBE_OUT203, LC_LOW_BIT_POS_PROBE_OUT202, 
    LC_LOW_BIT_POS_PROBE_OUT201, LC_LOW_BIT_POS_PROBE_OUT200, 
    LC_LOW_BIT_POS_PROBE_OUT199, LC_LOW_BIT_POS_PROBE_OUT198, 
    LC_LOW_BIT_POS_PROBE_OUT197, LC_LOW_BIT_POS_PROBE_OUT196, 
    LC_LOW_BIT_POS_PROBE_OUT195, LC_LOW_BIT_POS_PROBE_OUT194, 
    LC_LOW_BIT_POS_PROBE_OUT193, LC_LOW_BIT_POS_PROBE_OUT192, 
    LC_LOW_BIT_POS_PROBE_OUT191, LC_LOW_BIT_POS_PROBE_OUT190, 
    LC_LOW_BIT_POS_PROBE_OUT189, LC_LOW_BIT_POS_PROBE_OUT188, 
    LC_LOW_BIT_POS_PROBE_OUT187, LC_LOW_BIT_POS_PROBE_OUT186, 
    LC_LOW_BIT_POS_PROBE_OUT185, LC_LOW_BIT_POS_PROBE_OUT184, 
    LC_LOW_BIT_POS_PROBE_OUT183, LC_LOW_BIT_POS_PROBE_OUT182, 
    LC_LOW_BIT_POS_PROBE_OUT181, LC_LOW_BIT_POS_PROBE_OUT180, 
    LC_LOW_BIT_POS_PROBE_OUT179, LC_LOW_BIT_POS_PROBE_OUT178, 
    LC_LOW_BIT_POS_PROBE_OUT177, LC_LOW_BIT_POS_PROBE_OUT176, 
    LC_LOW_BIT_POS_PROBE_OUT175, LC_LOW_BIT_POS_PROBE_OUT174, 
    LC_LOW_BIT_POS_PROBE_OUT173, LC_LOW_BIT_POS_PROBE_OUT172, 
    LC_LOW_BIT_POS_PROBE_OUT171, LC_LOW_BIT_POS_PROBE_OUT170, 
    LC_LOW_BIT_POS_PROBE_OUT169, LC_LOW_BIT_POS_PROBE_OUT168, 
    LC_LOW_BIT_POS_PROBE_OUT167, LC_LOW_BIT_POS_PROBE_OUT166, 
    LC_LOW_BIT_POS_PROBE_OUT165, LC_LOW_BIT_POS_PROBE_OUT164, 
    LC_LOW_BIT_POS_PROBE_OUT163, LC_LOW_BIT_POS_PROBE_OUT162, 
    LC_LOW_BIT_POS_PROBE_OUT161, LC_LOW_BIT_POS_PROBE_OUT160, 
    LC_LOW_BIT_POS_PROBE_OUT159, LC_LOW_BIT_POS_PROBE_OUT158, 
    LC_LOW_BIT_POS_PROBE_OUT157, LC_LOW_BIT_POS_PROBE_OUT156, 
    LC_LOW_BIT_POS_PROBE_OUT155, LC_LOW_BIT_POS_PROBE_OUT154, 
    LC_LOW_BIT_POS_PROBE_OUT153, LC_LOW_BIT_POS_PROBE_OUT152, 
    LC_LOW_BIT_POS_PROBE_OUT151, LC_LOW_BIT_POS_PROBE_OUT150, 
    LC_LOW_BIT_POS_PROBE_OUT149, LC_LOW_BIT_POS_PROBE_OUT148, 
    LC_LOW_BIT_POS_PROBE_OUT147, LC_LOW_BIT_POS_PROBE_OUT146, 
    LC_LOW_BIT_POS_PROBE_OUT145, LC_LOW_BIT_POS_PROBE_OUT144, 
    LC_LOW_BIT_POS_PROBE_OUT143, LC_LOW_BIT_POS_PROBE_OUT142, 
    LC_LOW_BIT_POS_PROBE_OUT141, LC_LOW_BIT_POS_PROBE_OUT140, 
    LC_LOW_BIT_POS_PROBE_OUT139, LC_LOW_BIT_POS_PROBE_OUT138, 
    LC_LOW_BIT_POS_PROBE_OUT137, LC_LOW_BIT_POS_PROBE_OUT136, 
    LC_LOW_BIT_POS_PROBE_OUT135, LC_LOW_BIT_POS_PROBE_OUT134, 
    LC_LOW_BIT_POS_PROBE_OUT133, LC_LOW_BIT_POS_PROBE_OUT132, 
    LC_LOW_BIT_POS_PROBE_OUT131, LC_LOW_BIT_POS_PROBE_OUT130, 
    LC_LOW_BIT_POS_PROBE_OUT129, LC_LOW_BIT_POS_PROBE_OUT128, 
    LC_LOW_BIT_POS_PROBE_OUT127, LC_LOW_BIT_POS_PROBE_OUT126, 
    LC_LOW_BIT_POS_PROBE_OUT125, LC_LOW_BIT_POS_PROBE_OUT124, 
    LC_LOW_BIT_POS_PROBE_OUT123, LC_LOW_BIT_POS_PROBE_OUT122, 
    LC_LOW_BIT_POS_PROBE_OUT121, LC_LOW_BIT_POS_PROBE_OUT120, 
    LC_LOW_BIT_POS_PROBE_OUT119, LC_LOW_BIT_POS_PROBE_OUT118, 
    LC_LOW_BIT_POS_PROBE_OUT117, LC_LOW_BIT_POS_PROBE_OUT116, 
    LC_LOW_BIT_POS_PROBE_OUT115, LC_LOW_BIT_POS_PROBE_OUT114, 
    LC_LOW_BIT_POS_PROBE_OUT113, LC_LOW_BIT_POS_PROBE_OUT112, 
    LC_LOW_BIT_POS_PROBE_OUT111, LC_LOW_BIT_POS_PROBE_OUT110, 
    LC_LOW_BIT_POS_PROBE_OUT109, LC_LOW_BIT_POS_PROBE_OUT108, 
    LC_LOW_BIT_POS_PROBE_OUT107, LC_LOW_BIT_POS_PROBE_OUT106, 
    LC_LOW_BIT_POS_PROBE_OUT105, LC_LOW_BIT_POS_PROBE_OUT104, 
    LC_LOW_BIT_POS_PROBE_OUT103, LC_LOW_BIT_POS_PROBE_OUT102, 
    LC_LOW_BIT_POS_PROBE_OUT101, LC_LOW_BIT_POS_PROBE_OUT100, 
    LC_LOW_BIT_POS_PROBE_OUT99 , LC_LOW_BIT_POS_PROBE_OUT98 , 
    LC_LOW_BIT_POS_PROBE_OUT97 , LC_LOW_BIT_POS_PROBE_OUT96 , 
    LC_LOW_BIT_POS_PROBE_OUT95 , LC_LOW_BIT_POS_PROBE_OUT94 , 
    LC_LOW_BIT_POS_PROBE_OUT93 , LC_LOW_BIT_POS_PROBE_OUT92 , 
    LC_LOW_BIT_POS_PROBE_OUT91 , LC_LOW_BIT_POS_PROBE_OUT90 , 
    LC_LOW_BIT_POS_PROBE_OUT89 , LC_LOW_BIT_POS_PROBE_OUT88 , 
    LC_LOW_BIT_POS_PROBE_OUT87 , LC_LOW_BIT_POS_PROBE_OUT86 , 
    LC_LOW_BIT_POS_PROBE_OUT85 , LC_LOW_BIT_POS_PROBE_OUT84 , 
    LC_LOW_BIT_POS_PROBE_OUT83 , LC_LOW_BIT_POS_PROBE_OUT82 , 
    LC_LOW_BIT_POS_PROBE_OUT81 , LC_LOW_BIT_POS_PROBE_OUT80 , 
    LC_LOW_BIT_POS_PROBE_OUT79 , LC_LOW_BIT_POS_PROBE_OUT78 , 
    LC_LOW_BIT_POS_PROBE_OUT77 , LC_LOW_BIT_POS_PROBE_OUT76 , 
    LC_LOW_BIT_POS_PROBE_OUT75 , LC_LOW_BIT_POS_PROBE_OUT74 , 
    LC_LOW_BIT_POS_PROBE_OUT73 , LC_LOW_BIT_POS_PROBE_OUT72 , 
    LC_LOW_BIT_POS_PROBE_OUT71 , LC_LOW_BIT_POS_PROBE_OUT70 , 
    LC_LOW_BIT_POS_PROBE_OUT69 , LC_LOW_BIT_POS_PROBE_OUT68 , 
    LC_LOW_BIT_POS_PROBE_OUT67 , LC_LOW_BIT_POS_PROBE_OUT66 , 
    LC_LOW_BIT_POS_PROBE_OUT65 , LC_LOW_BIT_POS_PROBE_OUT64 , 
    LC_LOW_BIT_POS_PROBE_OUT63 , LC_LOW_BIT_POS_PROBE_OUT62 , 
    LC_LOW_BIT_POS_PROBE_OUT61 , LC_LOW_BIT_POS_PROBE_OUT60 , 
    LC_LOW_BIT_POS_PROBE_OUT59 , LC_LOW_BIT_POS_PROBE_OUT58 , 
    LC_LOW_BIT_POS_PROBE_OUT57 , LC_LOW_BIT_POS_PROBE_OUT56 , 
    LC_LOW_BIT_POS_PROBE_OUT55 , LC_LOW_BIT_POS_PROBE_OUT54 , 
    LC_LOW_BIT_POS_PROBE_OUT53 , LC_LOW_BIT_POS_PROBE_OUT52 , 
    LC_LOW_BIT_POS_PROBE_OUT51 , LC_LOW_BIT_POS_PROBE_OUT50 , 
    LC_LOW_BIT_POS_PROBE_OUT49 , LC_LOW_BIT_POS_PROBE_OUT48 , 
    LC_LOW_BIT_POS_PROBE_OUT47 , LC_LOW_BIT_POS_PROBE_OUT46 , 
    LC_LOW_BIT_POS_PROBE_OUT45 , LC_LOW_BIT_POS_PROBE_OUT44 , 
    LC_LOW_BIT_POS_PROBE_OUT43 , LC_LOW_BIT_POS_PROBE_OUT42 , 
    LC_LOW_BIT_POS_PROBE_OUT41 , LC_LOW_BIT_POS_PROBE_OUT40 , 
    LC_LOW_BIT_POS_PROBE_OUT39 , LC_LOW_BIT_POS_PROBE_OUT38 , 
    LC_LOW_BIT_POS_PROBE_OUT37 , LC_LOW_BIT_POS_PROBE_OUT36 , 
    LC_LOW_BIT_POS_PROBE_OUT35 , LC_LOW_BIT_POS_PROBE_OUT34 , 
    LC_LOW_BIT_POS_PROBE_OUT33 , LC_LOW_BIT_POS_PROBE_OUT32 , 
    LC_LOW_BIT_POS_PROBE_OUT31 , LC_LOW_BIT_POS_PROBE_OUT30 , 
    LC_LOW_BIT_POS_PROBE_OUT29 , LC_LOW_BIT_POS_PROBE_OUT28 , 
    LC_LOW_BIT_POS_PROBE_OUT27 , LC_LOW_BIT_POS_PROBE_OUT26 , 
    LC_LOW_BIT_POS_PROBE_OUT25 , LC_LOW_BIT_POS_PROBE_OUT24 , 
    LC_LOW_BIT_POS_PROBE_OUT23 , LC_LOW_BIT_POS_PROBE_OUT22 , 
    LC_LOW_BIT_POS_PROBE_OUT21 , LC_LOW_BIT_POS_PROBE_OUT20 , 
    LC_LOW_BIT_POS_PROBE_OUT19 , LC_LOW_BIT_POS_PROBE_OUT18 , 
    LC_LOW_BIT_POS_PROBE_OUT17 , LC_LOW_BIT_POS_PROBE_OUT16 , 
    LC_LOW_BIT_POS_PROBE_OUT15 , LC_LOW_BIT_POS_PROBE_OUT14 , 
    LC_LOW_BIT_POS_PROBE_OUT13 , LC_LOW_BIT_POS_PROBE_OUT12 , 
    LC_LOW_BIT_POS_PROBE_OUT11 , LC_LOW_BIT_POS_PROBE_OUT10 , 
    LC_LOW_BIT_POS_PROBE_OUT9  , LC_LOW_BIT_POS_PROBE_OUT8  , 
    LC_LOW_BIT_POS_PROBE_OUT7  , LC_LOW_BIT_POS_PROBE_OUT6  , 
    LC_LOW_BIT_POS_PROBE_OUT5  , LC_LOW_BIT_POS_PROBE_OUT4  , 
    LC_LOW_BIT_POS_PROBE_OUT3  , LC_LOW_BIT_POS_PROBE_OUT2  , 
    LC_LOW_BIT_POS_PROBE_OUT1  , LC_LOW_BIT_POS_PROBE_OUT0
  };
  
  localparam [(C_MAX_NUM_PROBE-C_NUM_PROBE_OUT)+LC_TOTAL_PROBE_OUT_WIDTH-1:0] 
    LC_PROBE_OUT_INIT_VAL_STRING = {
      C_PROBE_OUT255_INIT_VAL, C_PROBE_OUT254_INIT_VAL, C_PROBE_OUT253_INIT_VAL,
      C_PROBE_OUT252_INIT_VAL, C_PROBE_OUT251_INIT_VAL, C_PROBE_OUT250_INIT_VAL,
      C_PROBE_OUT249_INIT_VAL, C_PROBE_OUT248_INIT_VAL, C_PROBE_OUT247_INIT_VAL,
      C_PROBE_OUT246_INIT_VAL, C_PROBE_OUT245_INIT_VAL, C_PROBE_OUT244_INIT_VAL,
      C_PROBE_OUT243_INIT_VAL, C_PROBE_OUT242_INIT_VAL, C_PROBE_OUT241_INIT_VAL,
      C_PROBE_OUT240_INIT_VAL, C_PROBE_OUT239_INIT_VAL, C_PROBE_OUT238_INIT_VAL,
      C_PROBE_OUT237_INIT_VAL, C_PROBE_OUT236_INIT_VAL, C_PROBE_OUT235_INIT_VAL,
      C_PROBE_OUT234_INIT_VAL, C_PROBE_OUT233_INIT_VAL, C_PROBE_OUT232_INIT_VAL,
      C_PROBE_OUT231_INIT_VAL, C_PROBE_OUT230_INIT_VAL, C_PROBE_OUT229_INIT_VAL,
      C_PROBE_OUT228_INIT_VAL, C_PROBE_OUT227_INIT_VAL, C_PROBE_OUT226_INIT_VAL,
      C_PROBE_OUT225_INIT_VAL, C_PROBE_OUT224_INIT_VAL, C_PROBE_OUT223_INIT_VAL,
      C_PROBE_OUT222_INIT_VAL, C_PROBE_OUT221_INIT_VAL, C_PROBE_OUT220_INIT_VAL,
      C_PROBE_OUT219_INIT_VAL, C_PROBE_OUT218_INIT_VAL, C_PROBE_OUT217_INIT_VAL,
      C_PROBE_OUT216_INIT_VAL, C_PROBE_OUT215_INIT_VAL, C_PROBE_OUT214_INIT_VAL,
      C_PROBE_OUT213_INIT_VAL, C_PROBE_OUT212_INIT_VAL, C_PROBE_OUT211_INIT_VAL,
      C_PROBE_OUT210_INIT_VAL, C_PROBE_OUT209_INIT_VAL, C_PROBE_OUT208_INIT_VAL,
      C_PROBE_OUT207_INIT_VAL, C_PROBE_OUT206_INIT_VAL, C_PROBE_OUT205_INIT_VAL,
      C_PROBE_OUT204_INIT_VAL, C_PROBE_OUT203_INIT_VAL, C_PROBE_OUT202_INIT_VAL,
      C_PROBE_OUT201_INIT_VAL, C_PROBE_OUT200_INIT_VAL, C_PROBE_OUT199_INIT_VAL,
      C_PROBE_OUT198_INIT_VAL, C_PROBE_OUT197_INIT_VAL, C_PROBE_OUT196_INIT_VAL,
      C_PROBE_OUT195_INIT_VAL, C_PROBE_OUT194_INIT_VAL, C_PROBE_OUT193_INIT_VAL,
      C_PROBE_OUT192_INIT_VAL, C_PROBE_OUT191_INIT_VAL, C_PROBE_OUT190_INIT_VAL,
      C_PROBE_OUT189_INIT_VAL, C_PROBE_OUT188_INIT_VAL, C_PROBE_OUT187_INIT_VAL,
      C_PROBE_OUT186_INIT_VAL, C_PROBE_OUT185_INIT_VAL, C_PROBE_OUT184_INIT_VAL,
      C_PROBE_OUT183_INIT_VAL, C_PROBE_OUT182_INIT_VAL, C_PROBE_OUT181_INIT_VAL,
      C_PROBE_OUT180_INIT_VAL, C_PROBE_OUT179_INIT_VAL, C_PROBE_OUT178_INIT_VAL,
      C_PROBE_OUT177_INIT_VAL, C_PROBE_OUT176_INIT_VAL, C_PROBE_OUT175_INIT_VAL,
      C_PROBE_OUT174_INIT_VAL, C_PROBE_OUT173_INIT_VAL, C_PROBE_OUT172_INIT_VAL,
      C_PROBE_OUT171_INIT_VAL, C_PROBE_OUT170_INIT_VAL, C_PROBE_OUT169_INIT_VAL,
      C_PROBE_OUT168_INIT_VAL, C_PROBE_OUT167_INIT_VAL, C_PROBE_OUT166_INIT_VAL,
      C_PROBE_OUT165_INIT_VAL, C_PROBE_OUT164_INIT_VAL, C_PROBE_OUT163_INIT_VAL,
      C_PROBE_OUT162_INIT_VAL, C_PROBE_OUT161_INIT_VAL, C_PROBE_OUT160_INIT_VAL,
      C_PROBE_OUT159_INIT_VAL, C_PROBE_OUT158_INIT_VAL, C_PROBE_OUT157_INIT_VAL,
      C_PROBE_OUT156_INIT_VAL, C_PROBE_OUT155_INIT_VAL, C_PROBE_OUT154_INIT_VAL,
      C_PROBE_OUT153_INIT_VAL, C_PROBE_OUT152_INIT_VAL, C_PROBE_OUT151_INIT_VAL,
      C_PROBE_OUT150_INIT_VAL, C_PROBE_OUT149_INIT_VAL, C_PROBE_OUT148_INIT_VAL,
      C_PROBE_OUT147_INIT_VAL, C_PROBE_OUT146_INIT_VAL, C_PROBE_OUT145_INIT_VAL,
      C_PROBE_OUT144_INIT_VAL, C_PROBE_OUT143_INIT_VAL, C_PROBE_OUT142_INIT_VAL,
      C_PROBE_OUT141_INIT_VAL, C_PROBE_OUT140_INIT_VAL, C_PROBE_OUT139_INIT_VAL,
      C_PROBE_OUT138_INIT_VAL, C_PROBE_OUT137_INIT_VAL, C_PROBE_OUT136_INIT_VAL,
      C_PROBE_OUT135_INIT_VAL, C_PROBE_OUT134_INIT_VAL, C_PROBE_OUT133_INIT_VAL,
      C_PROBE_OUT132_INIT_VAL, C_PROBE_OUT131_INIT_VAL, C_PROBE_OUT130_INIT_VAL,
      C_PROBE_OUT129_INIT_VAL, C_PROBE_OUT128_INIT_VAL, C_PROBE_OUT127_INIT_VAL,
      C_PROBE_OUT126_INIT_VAL, C_PROBE_OUT125_INIT_VAL, C_PROBE_OUT124_INIT_VAL,
      C_PROBE_OUT123_INIT_VAL, C_PROBE_OUT122_INIT_VAL, C_PROBE_OUT121_INIT_VAL,
      C_PROBE_OUT120_INIT_VAL, C_PROBE_OUT119_INIT_VAL, C_PROBE_OUT118_INIT_VAL,
      C_PROBE_OUT117_INIT_VAL, C_PROBE_OUT116_INIT_VAL, C_PROBE_OUT115_INIT_VAL,
      C_PROBE_OUT114_INIT_VAL, C_PROBE_OUT113_INIT_VAL, C_PROBE_OUT112_INIT_VAL,
      C_PROBE_OUT111_INIT_VAL, C_PROBE_OUT110_INIT_VAL, C_PROBE_OUT109_INIT_VAL,
      C_PROBE_OUT108_INIT_VAL, C_PROBE_OUT107_INIT_VAL, C_PROBE_OUT106_INIT_VAL,
      C_PROBE_OUT105_INIT_VAL, C_PROBE_OUT104_INIT_VAL, C_PROBE_OUT103_INIT_VAL,
      C_PROBE_OUT102_INIT_VAL, C_PROBE_OUT101_INIT_VAL, C_PROBE_OUT100_INIT_VAL,
      C_PROBE_OUT99_INIT_VAL , C_PROBE_OUT98_INIT_VAL , C_PROBE_OUT97_INIT_VAL ,
      C_PROBE_OUT96_INIT_VAL , C_PROBE_OUT95_INIT_VAL , C_PROBE_OUT94_INIT_VAL ,
      C_PROBE_OUT93_INIT_VAL , C_PROBE_OUT92_INIT_VAL , C_PROBE_OUT91_INIT_VAL ,
      C_PROBE_OUT90_INIT_VAL , C_PROBE_OUT89_INIT_VAL , C_PROBE_OUT88_INIT_VAL ,
      C_PROBE_OUT87_INIT_VAL , C_PROBE_OUT86_INIT_VAL , C_PROBE_OUT85_INIT_VAL ,
      C_PROBE_OUT84_INIT_VAL , C_PROBE_OUT83_INIT_VAL , C_PROBE_OUT82_INIT_VAL ,
      C_PROBE_OUT81_INIT_VAL , C_PROBE_OUT80_INIT_VAL , C_PROBE_OUT79_INIT_VAL ,
      C_PROBE_OUT78_INIT_VAL , C_PROBE_OUT77_INIT_VAL , C_PROBE_OUT76_INIT_VAL ,
      C_PROBE_OUT75_INIT_VAL , C_PROBE_OUT74_INIT_VAL , C_PROBE_OUT73_INIT_VAL ,
      C_PROBE_OUT72_INIT_VAL , C_PROBE_OUT71_INIT_VAL , C_PROBE_OUT70_INIT_VAL ,
      C_PROBE_OUT69_INIT_VAL , C_PROBE_OUT68_INIT_VAL , C_PROBE_OUT67_INIT_VAL ,
      C_PROBE_OUT66_INIT_VAL , C_PROBE_OUT65_INIT_VAL , C_PROBE_OUT64_INIT_VAL ,
      C_PROBE_OUT63_INIT_VAL , C_PROBE_OUT62_INIT_VAL , C_PROBE_OUT61_INIT_VAL ,
      C_PROBE_OUT60_INIT_VAL , C_PROBE_OUT59_INIT_VAL , C_PROBE_OUT58_INIT_VAL ,
      C_PROBE_OUT57_INIT_VAL , C_PROBE_OUT56_INIT_VAL , C_PROBE_OUT55_INIT_VAL ,
      C_PROBE_OUT54_INIT_VAL , C_PROBE_OUT53_INIT_VAL , C_PROBE_OUT52_INIT_VAL ,
      C_PROBE_OUT51_INIT_VAL , C_PROBE_OUT50_INIT_VAL , C_PROBE_OUT49_INIT_VAL ,
      C_PROBE_OUT48_INIT_VAL , C_PROBE_OUT47_INIT_VAL , C_PROBE_OUT46_INIT_VAL ,
      C_PROBE_OUT45_INIT_VAL , C_PROBE_OUT44_INIT_VAL , C_PROBE_OUT43_INIT_VAL ,
      C_PROBE_OUT42_INIT_VAL , C_PROBE_OUT41_INIT_VAL , C_PROBE_OUT40_INIT_VAL ,
      C_PROBE_OUT39_INIT_VAL , C_PROBE_OUT38_INIT_VAL , C_PROBE_OUT37_INIT_VAL ,
      C_PROBE_OUT36_INIT_VAL , C_PROBE_OUT35_INIT_VAL , C_PROBE_OUT34_INIT_VAL ,
      C_PROBE_OUT33_INIT_VAL , C_PROBE_OUT32_INIT_VAL , C_PROBE_OUT31_INIT_VAL ,
      C_PROBE_OUT30_INIT_VAL , C_PROBE_OUT29_INIT_VAL , C_PROBE_OUT28_INIT_VAL ,
      C_PROBE_OUT27_INIT_VAL , C_PROBE_OUT26_INIT_VAL , C_PROBE_OUT25_INIT_VAL ,
      C_PROBE_OUT24_INIT_VAL , C_PROBE_OUT23_INIT_VAL , C_PROBE_OUT22_INIT_VAL ,
      C_PROBE_OUT21_INIT_VAL , C_PROBE_OUT20_INIT_VAL , C_PROBE_OUT19_INIT_VAL ,
      C_PROBE_OUT18_INIT_VAL , C_PROBE_OUT17_INIT_VAL , C_PROBE_OUT16_INIT_VAL ,
      C_PROBE_OUT15_INIT_VAL , C_PROBE_OUT14_INIT_VAL , C_PROBE_OUT13_INIT_VAL ,
      C_PROBE_OUT12_INIT_VAL , C_PROBE_OUT11_INIT_VAL , C_PROBE_OUT10_INIT_VAL ,
      C_PROBE_OUT9_INIT_VAL  , C_PROBE_OUT8_INIT_VAL  , C_PROBE_OUT7_INIT_VAL  ,
      C_PROBE_OUT6_INIT_VAL  , C_PROBE_OUT5_INIT_VAL  , C_PROBE_OUT4_INIT_VAL  ,
      C_PROBE_OUT3_INIT_VAL  , C_PROBE_OUT2_INIT_VAL  , C_PROBE_OUT1_INIT_VAL  ,
      C_PROBE_OUT0_INIT_VAL
    };

