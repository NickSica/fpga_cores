 reg [C_PROBE0_WIDTH-1:0]  mem_shift_probe0;
 reg [C_PROBE1_WIDTH-1:0]  mem_shift_probe1;
 reg [C_PROBE2_WIDTH-1:0]  mem_shift_probe2;
 reg [C_PROBE3_WIDTH-1:0]  mem_shift_probe3;
 reg [C_PROBE4_WIDTH-1:0]  mem_shift_probe4;
 reg [C_PROBE5_WIDTH-1:0]  mem_shift_probe5;
 reg [C_PROBE6_WIDTH-1:0]  mem_shift_probe6;
 reg [C_PROBE7_WIDTH-1:0]  mem_shift_probe7;
 reg [C_PROBE8_WIDTH-1:0]  mem_shift_probe8;
 reg [C_PROBE9_WIDTH-1:0]  mem_shift_probe9;
 reg [C_PROBE10_WIDTH-1:0] mem_shift_probe10  ;
 reg [C_PROBE11_WIDTH-1:0] mem_shift_probe11  ;
 reg [C_PROBE12_WIDTH-1:0] mem_shift_probe12  ;
 reg [C_PROBE13_WIDTH-1:0] mem_shift_probe13  ;
 reg [C_PROBE14_WIDTH-1:0] mem_shift_probe14  ;
 reg [C_PROBE15_WIDTH-1:0] mem_shift_probe15  ;
 reg [C_PROBE16_WIDTH-1:0] mem_shift_probe16  ;
 reg [C_PROBE17_WIDTH-1:0] mem_shift_probe17  ;
 reg [C_PROBE18_WIDTH-1:0] mem_shift_probe18  ;
 reg [C_PROBE19_WIDTH-1:0] mem_shift_probe19  ;
 reg [C_PROBE20_WIDTH-1:0] mem_shift_probe20  ;
 reg [C_PROBE21_WIDTH-1:0] mem_shift_probe21  ;
 reg [C_PROBE22_WIDTH-1:0] mem_shift_probe22  ;
 reg [C_PROBE23_WIDTH-1:0] mem_shift_probe23  ;
 reg [C_PROBE24_WIDTH-1:0] mem_shift_probe24  ;
 reg [C_PROBE25_WIDTH-1:0] mem_shift_probe25  ;
 reg [C_PROBE26_WIDTH-1:0] mem_shift_probe26  ;
 reg [C_PROBE27_WIDTH-1:0] mem_shift_probe27  ;
 reg [C_PROBE28_WIDTH-1:0] mem_shift_probe28  ;
 reg [C_PROBE29_WIDTH-1:0] mem_shift_probe29  ;
 reg [C_PROBE30_WIDTH-1:0] mem_shift_probe30  ;
 reg [C_PROBE31_WIDTH-1:0] mem_shift_probe31  ;
 reg [C_PROBE32_WIDTH-1:0] mem_shift_probe32  ;
 reg [C_PROBE33_WIDTH-1:0] mem_shift_probe33  ;
 reg [C_PROBE34_WIDTH-1:0] mem_shift_probe34  ;
 reg [C_PROBE35_WIDTH-1:0] mem_shift_probe35  ;
 reg [C_PROBE36_WIDTH-1:0] mem_shift_probe36  ;
 reg [C_PROBE37_WIDTH-1:0] mem_shift_probe37  ;
 reg [C_PROBE38_WIDTH-1:0] mem_shift_probe38  ;
 reg [C_PROBE39_WIDTH-1:0] mem_shift_probe39  ;
 reg [C_PROBE40_WIDTH-1:0] mem_shift_probe40  ;
 reg [C_PROBE41_WIDTH-1:0] mem_shift_probe41  ;
 reg [C_PROBE42_WIDTH-1:0] mem_shift_probe42  ;
 reg [C_PROBE43_WIDTH-1:0] mem_shift_probe43  ;
 reg [C_PROBE44_WIDTH-1:0] mem_shift_probe44  ;
 reg [C_PROBE45_WIDTH-1:0] mem_shift_probe45  ;
 reg [C_PROBE46_WIDTH-1:0] mem_shift_probe46  ;
 reg [C_PROBE47_WIDTH-1:0] mem_shift_probe47  ;
 reg [C_PROBE48_WIDTH-1:0] mem_shift_probe48  ;
 reg [C_PROBE49_WIDTH-1:0] mem_shift_probe49  ;
 reg [C_PROBE50_WIDTH-1:0] mem_shift_probe50  ;
 reg [C_PROBE51_WIDTH-1:0] mem_shift_probe51  ;
 reg [C_PROBE52_WIDTH-1:0] mem_shift_probe52  ;
 reg [C_PROBE53_WIDTH-1:0] mem_shift_probe53  ;
 reg [C_PROBE54_WIDTH-1:0] mem_shift_probe54  ;
 reg [C_PROBE55_WIDTH-1:0] mem_shift_probe55  ;
 reg [C_PROBE56_WIDTH-1:0] mem_shift_probe56  ;
 reg [C_PROBE57_WIDTH-1:0] mem_shift_probe57  ;
 reg [C_PROBE58_WIDTH-1:0] mem_shift_probe58  ;
 reg [C_PROBE59_WIDTH-1:0] mem_shift_probe59  ;
 reg [C_PROBE60_WIDTH-1:0] mem_shift_probe60  ;
 reg [C_PROBE61_WIDTH-1:0] mem_shift_probe61  ;
 reg [C_PROBE62_WIDTH-1:0] mem_shift_probe62  ;
 reg [C_PROBE63_WIDTH-1:0] mem_shift_probe63  ;
 reg [C_PROBE64_WIDTH-1:0] mem_shift_probe64  ;
 reg [C_PROBE65_WIDTH-1:0] mem_shift_probe65  ;
 reg [C_PROBE66_WIDTH-1:0] mem_shift_probe66  ;
 reg [C_PROBE67_WIDTH-1:0] mem_shift_probe67  ;
 reg [C_PROBE68_WIDTH-1:0] mem_shift_probe68  ;
 reg [C_PROBE69_WIDTH-1:0] mem_shift_probe69  ;
 reg [C_PROBE70_WIDTH-1:0] mem_shift_probe70  ;
 reg [C_PROBE71_WIDTH-1:0] mem_shift_probe71  ;
 reg [C_PROBE72_WIDTH-1:0] mem_shift_probe72  ;
 reg [C_PROBE73_WIDTH-1:0] mem_shift_probe73  ;
 reg [C_PROBE74_WIDTH-1:0] mem_shift_probe74  ;
 reg [C_PROBE75_WIDTH-1:0] mem_shift_probe75  ;
 reg [C_PROBE76_WIDTH-1:0] mem_shift_probe76  ;
 reg [C_PROBE77_WIDTH-1:0] mem_shift_probe77  ;
 reg [C_PROBE78_WIDTH-1:0] mem_shift_probe78  ;
 reg [C_PROBE79_WIDTH-1:0] mem_shift_probe79  ;
 reg [C_PROBE80_WIDTH-1:0] mem_shift_probe80  ;
 reg [C_PROBE81_WIDTH-1:0] mem_shift_probe81  ;
 reg [C_PROBE82_WIDTH-1:0] mem_shift_probe82  ;
 reg [C_PROBE83_WIDTH-1:0] mem_shift_probe83  ;
 reg [C_PROBE84_WIDTH-1:0] mem_shift_probe84  ;
 reg [C_PROBE85_WIDTH-1:0] mem_shift_probe85  ;
 reg [C_PROBE86_WIDTH-1:0] mem_shift_probe86  ;
 reg [C_PROBE87_WIDTH-1:0] mem_shift_probe87  ;
 reg [C_PROBE88_WIDTH-1:0] mem_shift_probe88  ;
 reg [C_PROBE89_WIDTH-1:0] mem_shift_probe89  ;
 reg [C_PROBE90_WIDTH-1:0] mem_shift_probe90  ;
 reg [C_PROBE91_WIDTH-1:0] mem_shift_probe91  ;
 reg [C_PROBE92_WIDTH-1:0] mem_shift_probe92  ;
 reg [C_PROBE93_WIDTH-1:0] mem_shift_probe93  ;
 reg [C_PROBE94_WIDTH-1:0] mem_shift_probe94  ;
 reg [C_PROBE95_WIDTH-1:0] mem_shift_probe95  ;
 reg [C_PROBE96_WIDTH-1:0] mem_shift_probe96  ;
 reg [C_PROBE97_WIDTH-1:0] mem_shift_probe97  ;
 reg [C_PROBE98_WIDTH-1:0] mem_shift_probe98  ;
 reg [C_PROBE99_WIDTH-1:0] mem_shift_probe99  ;
 reg [C_PROBE100_WIDTH-1:0]mem_shift_probe100  ;
 reg [C_PROBE101_WIDTH-1:0]mem_shift_probe101  ;
 reg [C_PROBE102_WIDTH-1:0]mem_shift_probe102  ;
 reg [C_PROBE103_WIDTH-1:0]mem_shift_probe103  ;
 reg [C_PROBE104_WIDTH-1:0]mem_shift_probe104  ;
 reg [C_PROBE105_WIDTH-1:0]mem_shift_probe105  ;
 reg [C_PROBE106_WIDTH-1:0]mem_shift_probe106  ;
 reg [C_PROBE107_WIDTH-1:0]mem_shift_probe107  ;
 reg [C_PROBE108_WIDTH-1:0]mem_shift_probe108  ;
 reg [C_PROBE109_WIDTH-1:0]mem_shift_probe109  ;
 reg [C_PROBE110_WIDTH-1:0]mem_shift_probe110  ;
 reg [C_PROBE111_WIDTH-1:0]mem_shift_probe111  ;
 reg [C_PROBE112_WIDTH-1:0]mem_shift_probe112  ;
 reg [C_PROBE113_WIDTH-1:0]mem_shift_probe113  ;
 reg [C_PROBE114_WIDTH-1:0]mem_shift_probe114  ;
 reg [C_PROBE115_WIDTH-1:0]mem_shift_probe115  ;
 reg [C_PROBE116_WIDTH-1:0]mem_shift_probe116  ;
 reg [C_PROBE117_WIDTH-1:0]mem_shift_probe117  ;
 reg [C_PROBE118_WIDTH-1:0]mem_shift_probe118  ;
 reg [C_PROBE119_WIDTH-1:0]mem_shift_probe119  ;
 reg [C_PROBE120_WIDTH-1:0]mem_shift_probe120  ;
 reg [C_PROBE121_WIDTH-1:0]mem_shift_probe121  ;
 reg [C_PROBE122_WIDTH-1:0]mem_shift_probe122  ;
 reg [C_PROBE123_WIDTH-1:0]mem_shift_probe123  ;
 reg [C_PROBE124_WIDTH-1:0]mem_shift_probe124  ;
 reg [C_PROBE125_WIDTH-1:0]mem_shift_probe125  ;
 reg [C_PROBE126_WIDTH-1:0]mem_shift_probe126  ;
 reg [C_PROBE127_WIDTH-1:0]mem_shift_probe127  ;
 reg [C_PROBE128_WIDTH-1:0]mem_shift_probe128  ;
 reg [C_PROBE129_WIDTH-1:0]mem_shift_probe129  ;
 reg [C_PROBE130_WIDTH-1:0]mem_shift_probe130  ;
 reg [C_PROBE131_WIDTH-1:0]mem_shift_probe131  ;
 reg [C_PROBE132_WIDTH-1:0]mem_shift_probe132  ;
 reg [C_PROBE133_WIDTH-1:0]mem_shift_probe133  ;
 reg [C_PROBE134_WIDTH-1:0]mem_shift_probe134  ;
 reg [C_PROBE135_WIDTH-1:0]mem_shift_probe135  ;
 reg [C_PROBE136_WIDTH-1:0]mem_shift_probe136  ;
 reg [C_PROBE137_WIDTH-1:0]mem_shift_probe137  ;
 reg [C_PROBE138_WIDTH-1:0]mem_shift_probe138  ;
 reg [C_PROBE139_WIDTH-1:0]mem_shift_probe139  ;
 reg [C_PROBE140_WIDTH-1:0]mem_shift_probe140  ;
 reg [C_PROBE141_WIDTH-1:0]mem_shift_probe141  ;
 reg [C_PROBE142_WIDTH-1:0]mem_shift_probe142  ;
 reg [C_PROBE143_WIDTH-1:0]mem_shift_probe143  ;
 reg [C_PROBE144_WIDTH-1:0]mem_shift_probe144  ;
 reg [C_PROBE145_WIDTH-1:0]mem_shift_probe145  ;
 reg [C_PROBE146_WIDTH-1:0]mem_shift_probe146  ;
 reg [C_PROBE147_WIDTH-1:0]mem_shift_probe147  ;
 reg [C_PROBE148_WIDTH-1:0]mem_shift_probe148  ;
 reg [C_PROBE149_WIDTH-1:0]mem_shift_probe149  ;
 reg [C_PROBE150_WIDTH-1:0]mem_shift_probe150  ;
 reg [C_PROBE151_WIDTH-1:0]mem_shift_probe151  ;
 reg [C_PROBE152_WIDTH-1:0]mem_shift_probe152  ;
 reg [C_PROBE153_WIDTH-1:0]mem_shift_probe153  ;
 reg [C_PROBE154_WIDTH-1:0]mem_shift_probe154  ;
 reg [C_PROBE155_WIDTH-1:0]mem_shift_probe155  ;
 reg [C_PROBE156_WIDTH-1:0]mem_shift_probe156  ;
 reg [C_PROBE157_WIDTH-1:0]mem_shift_probe157  ;
 reg [C_PROBE158_WIDTH-1:0]mem_shift_probe158  ;
 reg [C_PROBE159_WIDTH-1:0]mem_shift_probe159  ;
 reg [C_PROBE160_WIDTH-1:0]mem_shift_probe160  ;
 reg [C_PROBE161_WIDTH-1:0]mem_shift_probe161  ;
 reg [C_PROBE162_WIDTH-1:0]mem_shift_probe162  ;
 reg [C_PROBE163_WIDTH-1:0]mem_shift_probe163  ;
 reg [C_PROBE164_WIDTH-1:0]mem_shift_probe164  ;
 reg [C_PROBE165_WIDTH-1:0]mem_shift_probe165  ;
 reg [C_PROBE166_WIDTH-1:0]mem_shift_probe166  ;
 reg [C_PROBE167_WIDTH-1:0]mem_shift_probe167  ;
 reg [C_PROBE168_WIDTH-1:0]mem_shift_probe168  ;
 reg [C_PROBE169_WIDTH-1:0]mem_shift_probe169  ;
 reg [C_PROBE170_WIDTH-1:0]mem_shift_probe170  ;
 reg [C_PROBE171_WIDTH-1:0]mem_shift_probe171  ;
 reg [C_PROBE172_WIDTH-1:0]mem_shift_probe172  ;
 reg [C_PROBE173_WIDTH-1:0]mem_shift_probe173  ;
 reg [C_PROBE174_WIDTH-1:0]mem_shift_probe174  ;
 reg [C_PROBE175_WIDTH-1:0]mem_shift_probe175  ;
 reg [C_PROBE176_WIDTH-1:0]mem_shift_probe176  ;
 reg [C_PROBE177_WIDTH-1:0]mem_shift_probe177  ;
 reg [C_PROBE178_WIDTH-1:0]mem_shift_probe178  ;
 reg [C_PROBE179_WIDTH-1:0]mem_shift_probe179  ;
 reg [C_PROBE180_WIDTH-1:0]mem_shift_probe180  ;
 reg [C_PROBE181_WIDTH-1:0]mem_shift_probe181  ;
 reg [C_PROBE182_WIDTH-1:0]mem_shift_probe182  ;
 reg [C_PROBE183_WIDTH-1:0]mem_shift_probe183  ;
 reg [C_PROBE184_WIDTH-1:0]mem_shift_probe184  ;
 reg [C_PROBE185_WIDTH-1:0]mem_shift_probe185  ;
 reg [C_PROBE186_WIDTH-1:0]mem_shift_probe186  ;
 reg [C_PROBE187_WIDTH-1:0]mem_shift_probe187  ;
 reg [C_PROBE188_WIDTH-1:0]mem_shift_probe188  ;
 reg [C_PROBE189_WIDTH-1:0]mem_shift_probe189  ;
 reg [C_PROBE190_WIDTH-1:0]mem_shift_probe190  ;
 reg [C_PROBE191_WIDTH-1:0]mem_shift_probe191  ;
 reg [C_PROBE192_WIDTH-1:0]mem_shift_probe192  ;
 reg [C_PROBE193_WIDTH-1:0]mem_shift_probe193  ;
 reg [C_PROBE194_WIDTH-1:0]mem_shift_probe194  ;
 reg [C_PROBE195_WIDTH-1:0]mem_shift_probe195  ;
 reg [C_PROBE196_WIDTH-1:0]mem_shift_probe196  ;
 reg [C_PROBE197_WIDTH-1:0]mem_shift_probe197  ;
 reg [C_PROBE198_WIDTH-1:0]mem_shift_probe198  ;
 reg [C_PROBE199_WIDTH-1:0]mem_shift_probe199  ;
 reg [C_PROBE200_WIDTH-1:0]mem_shift_probe200  ;
 reg [C_PROBE201_WIDTH-1:0]mem_shift_probe201  ;
 reg [C_PROBE202_WIDTH-1:0]mem_shift_probe202  ;
 reg [C_PROBE203_WIDTH-1:0]mem_shift_probe203  ;
 reg [C_PROBE204_WIDTH-1:0]mem_shift_probe204  ;
 reg [C_PROBE205_WIDTH-1:0]mem_shift_probe205  ;
 reg [C_PROBE206_WIDTH-1:0]mem_shift_probe206  ;
 reg [C_PROBE207_WIDTH-1:0]mem_shift_probe207  ;
 reg [C_PROBE208_WIDTH-1:0]mem_shift_probe208  ;
 reg [C_PROBE209_WIDTH-1:0]mem_shift_probe209  ;
 reg [C_PROBE210_WIDTH-1:0]mem_shift_probe210  ;
 reg [C_PROBE211_WIDTH-1:0]mem_shift_probe211  ;
 reg [C_PROBE212_WIDTH-1:0]mem_shift_probe212  ;
 reg [C_PROBE213_WIDTH-1:0]mem_shift_probe213  ;
 reg [C_PROBE214_WIDTH-1:0]mem_shift_probe214  ;
 reg [C_PROBE215_WIDTH-1:0]mem_shift_probe215  ;
 reg [C_PROBE216_WIDTH-1:0]mem_shift_probe216  ;
 reg [C_PROBE217_WIDTH-1:0]mem_shift_probe217  ;
 reg [C_PROBE218_WIDTH-1:0]mem_shift_probe218  ;
 reg [C_PROBE219_WIDTH-1:0]mem_shift_probe219  ;
 reg [C_PROBE220_WIDTH-1:0]mem_shift_probe220  ;
 reg [C_PROBE221_WIDTH-1:0]mem_shift_probe221  ;
 reg [C_PROBE222_WIDTH-1:0]mem_shift_probe222  ;
 reg [C_PROBE223_WIDTH-1:0]mem_shift_probe223  ;
 reg [C_PROBE224_WIDTH-1:0]mem_shift_probe224  ;
 reg [C_PROBE225_WIDTH-1:0]mem_shift_probe225  ;
 reg [C_PROBE226_WIDTH-1:0]mem_shift_probe226  ;
 reg [C_PROBE227_WIDTH-1:0]mem_shift_probe227  ;
 reg [C_PROBE228_WIDTH-1:0]mem_shift_probe228  ;
 reg [C_PROBE229_WIDTH-1:0]mem_shift_probe229  ;
 reg [C_PROBE230_WIDTH-1:0]mem_shift_probe230  ;
 reg [C_PROBE231_WIDTH-1:0]mem_shift_probe231  ;
 reg [C_PROBE232_WIDTH-1:0]mem_shift_probe232  ;
 reg [C_PROBE233_WIDTH-1:0]mem_shift_probe233  ;
 reg [C_PROBE234_WIDTH-1:0]mem_shift_probe234  ;
 reg [C_PROBE235_WIDTH-1:0]mem_shift_probe235  ;
 reg [C_PROBE236_WIDTH-1:0]mem_shift_probe236  ;
 reg [C_PROBE237_WIDTH-1:0]mem_shift_probe237  ;
 reg [C_PROBE238_WIDTH-1:0]mem_shift_probe238  ;
 reg [C_PROBE239_WIDTH-1:0]mem_shift_probe239  ;
 reg [C_PROBE240_WIDTH-1:0]mem_shift_probe240  ;
 reg [C_PROBE241_WIDTH-1:0]mem_shift_probe241  ;
 reg [C_PROBE242_WIDTH-1:0]mem_shift_probe242  ;
 reg [C_PROBE243_WIDTH-1:0]mem_shift_probe243  ;
 reg [C_PROBE244_WIDTH-1:0]mem_shift_probe244  ;
 reg [C_PROBE245_WIDTH-1:0]mem_shift_probe245  ;
 reg [C_PROBE246_WIDTH-1:0]mem_shift_probe246  ;
 reg [C_PROBE247_WIDTH-1:0]mem_shift_probe247  ;
 reg [C_PROBE248_WIDTH-1:0]mem_shift_probe248  ;
 reg [C_PROBE249_WIDTH-1:0]mem_shift_probe249  ;
 reg [C_PROBE250_WIDTH-1:0]mem_shift_probe250  ;
 reg [C_PROBE251_WIDTH-1:0]mem_shift_probe251  ;
 reg [C_PROBE252_WIDTH-1:0]mem_shift_probe252  ;
 reg [C_PROBE253_WIDTH-1:0]mem_shift_probe253  ;
 reg [C_PROBE254_WIDTH-1:0]mem_shift_probe254  ;
 reg [C_PROBE255_WIDTH-1:0]mem_shift_probe255  ;
 reg [C_PROBE256_WIDTH-1:0]mem_shift_probe256  ;
 reg [C_PROBE257_WIDTH-1:0]mem_shift_probe257  ;
 reg [C_PROBE258_WIDTH-1:0]mem_shift_probe258  ;
 reg [C_PROBE259_WIDTH-1:0]mem_shift_probe259  ;
 reg [C_PROBE260_WIDTH-1:0]mem_shift_probe260  ;
 reg [C_PROBE261_WIDTH-1:0]mem_shift_probe261  ;
 reg [C_PROBE262_WIDTH-1:0]mem_shift_probe262  ;
 reg [C_PROBE263_WIDTH-1:0]mem_shift_probe263  ;
 reg [C_PROBE264_WIDTH-1:0]mem_shift_probe264  ;
 reg [C_PROBE265_WIDTH-1:0]mem_shift_probe265  ;
 reg [C_PROBE266_WIDTH-1:0]mem_shift_probe266  ;
 reg [C_PROBE267_WIDTH-1:0]mem_shift_probe267  ;
 reg [C_PROBE268_WIDTH-1:0]mem_shift_probe268  ;
 reg [C_PROBE269_WIDTH-1:0]mem_shift_probe269  ;
 reg [C_PROBE270_WIDTH-1:0]mem_shift_probe270  ;
 reg [C_PROBE271_WIDTH-1:0]mem_shift_probe271  ;
 reg [C_PROBE272_WIDTH-1:0]mem_shift_probe272  ;
 reg [C_PROBE273_WIDTH-1:0]mem_shift_probe273  ;
 reg [C_PROBE274_WIDTH-1:0]mem_shift_probe274  ;
 reg [C_PROBE275_WIDTH-1:0]mem_shift_probe275  ;
 reg [C_PROBE276_WIDTH-1:0]mem_shift_probe276  ;
 reg [C_PROBE277_WIDTH-1:0]mem_shift_probe277  ;
 reg [C_PROBE278_WIDTH-1:0]mem_shift_probe278  ;
 reg [C_PROBE279_WIDTH-1:0]mem_shift_probe279  ;
 reg [C_PROBE280_WIDTH-1:0]mem_shift_probe280  ;
 reg [C_PROBE281_WIDTH-1:0]mem_shift_probe281  ;
 reg [C_PROBE282_WIDTH-1:0]mem_shift_probe282  ;
 reg [C_PROBE283_WIDTH-1:0]mem_shift_probe283  ;
 reg [C_PROBE284_WIDTH-1:0]mem_shift_probe284  ;
 reg [C_PROBE285_WIDTH-1:0]mem_shift_probe285  ;
 reg [C_PROBE286_WIDTH-1:0]mem_shift_probe286  ;
 reg [C_PROBE287_WIDTH-1:0]mem_shift_probe287  ;
 reg [C_PROBE288_WIDTH-1:0]mem_shift_probe288  ;
 reg [C_PROBE289_WIDTH-1:0]mem_shift_probe289  ;
 reg [C_PROBE290_WIDTH-1:0]mem_shift_probe290  ;
 reg [C_PROBE291_WIDTH-1:0]mem_shift_probe291  ;
 reg [C_PROBE292_WIDTH-1:0]mem_shift_probe292  ;
 reg [C_PROBE293_WIDTH-1:0]mem_shift_probe293  ;
 reg [C_PROBE294_WIDTH-1:0]mem_shift_probe294  ;
 reg [C_PROBE295_WIDTH-1:0]mem_shift_probe295  ;
 reg [C_PROBE296_WIDTH-1:0]mem_shift_probe296  ;
 reg [C_PROBE297_WIDTH-1:0]mem_shift_probe297  ;
 reg [C_PROBE298_WIDTH-1:0]mem_shift_probe298  ;
 reg [C_PROBE299_WIDTH-1:0]mem_shift_probe299  ;
 reg [C_PROBE300_WIDTH-1:0]mem_shift_probe300  ;
 reg [C_PROBE301_WIDTH-1:0]mem_shift_probe301  ;
 reg [C_PROBE302_WIDTH-1:0]mem_shift_probe302  ;
 reg [C_PROBE303_WIDTH-1:0]mem_shift_probe303  ;
 reg [C_PROBE304_WIDTH-1:0]mem_shift_probe304  ;
 reg [C_PROBE305_WIDTH-1:0]mem_shift_probe305  ;
 reg [C_PROBE306_WIDTH-1:0]mem_shift_probe306  ;
 reg [C_PROBE307_WIDTH-1:0]mem_shift_probe307  ;
 reg [C_PROBE308_WIDTH-1:0]mem_shift_probe308  ;
 reg [C_PROBE309_WIDTH-1:0]mem_shift_probe309  ;
 reg [C_PROBE310_WIDTH-1:0]mem_shift_probe310  ;
 reg [C_PROBE311_WIDTH-1:0]mem_shift_probe311  ;
 reg [C_PROBE312_WIDTH-1:0]mem_shift_probe312  ;
 reg [C_PROBE313_WIDTH-1:0]mem_shift_probe313  ;
 reg [C_PROBE314_WIDTH-1:0]mem_shift_probe314  ;
 reg [C_PROBE315_WIDTH-1:0]mem_shift_probe315  ;
 reg [C_PROBE316_WIDTH-1:0]mem_shift_probe316  ;
 reg [C_PROBE317_WIDTH-1:0]mem_shift_probe317  ;
 reg [C_PROBE318_WIDTH-1:0]mem_shift_probe318  ;
 reg [C_PROBE319_WIDTH-1:0]mem_shift_probe319  ;
 reg [C_PROBE320_WIDTH-1:0]mem_shift_probe320  ;
 reg [C_PROBE321_WIDTH-1:0]mem_shift_probe321  ;
 reg [C_PROBE322_WIDTH-1:0]mem_shift_probe322  ;
 reg [C_PROBE323_WIDTH-1:0]mem_shift_probe323  ;
 reg [C_PROBE324_WIDTH-1:0]mem_shift_probe324  ;
 reg [C_PROBE325_WIDTH-1:0]mem_shift_probe325  ;
 reg [C_PROBE326_WIDTH-1:0]mem_shift_probe326  ;
 reg [C_PROBE327_WIDTH-1:0]mem_shift_probe327  ;
 reg [C_PROBE328_WIDTH-1:0]mem_shift_probe328  ;
 reg [C_PROBE329_WIDTH-1:0]mem_shift_probe329  ;
 reg [C_PROBE330_WIDTH-1:0]mem_shift_probe330  ;
 reg [C_PROBE331_WIDTH-1:0]mem_shift_probe331  ;
 reg [C_PROBE332_WIDTH-1:0]mem_shift_probe332  ;
 reg [C_PROBE333_WIDTH-1:0]mem_shift_probe333  ;
 reg [C_PROBE334_WIDTH-1:0]mem_shift_probe334  ;
 reg [C_PROBE335_WIDTH-1:0]mem_shift_probe335  ;
 reg [C_PROBE336_WIDTH-1:0]mem_shift_probe336  ;
 reg [C_PROBE337_WIDTH-1:0]mem_shift_probe337  ;
 reg [C_PROBE338_WIDTH-1:0]mem_shift_probe338  ;
 reg [C_PROBE339_WIDTH-1:0]mem_shift_probe339  ;
 reg [C_PROBE340_WIDTH-1:0]mem_shift_probe340  ;
 reg [C_PROBE341_WIDTH-1:0]mem_shift_probe341  ;
 reg [C_PROBE342_WIDTH-1:0]mem_shift_probe342  ;
 reg [C_PROBE343_WIDTH-1:0]mem_shift_probe343  ;
 reg [C_PROBE344_WIDTH-1:0]mem_shift_probe344  ;
 reg [C_PROBE345_WIDTH-1:0]mem_shift_probe345  ;
 reg [C_PROBE346_WIDTH-1:0]mem_shift_probe346  ;
 reg [C_PROBE347_WIDTH-1:0]mem_shift_probe347  ;
 reg [C_PROBE348_WIDTH-1:0]mem_shift_probe348  ;
 reg [C_PROBE349_WIDTH-1:0]mem_shift_probe349  ;
 reg [C_PROBE350_WIDTH-1:0]mem_shift_probe350  ;
 reg [C_PROBE351_WIDTH-1:0]mem_shift_probe351  ;
 reg [C_PROBE352_WIDTH-1:0]mem_shift_probe352  ;
 reg [C_PROBE353_WIDTH-1:0]mem_shift_probe353  ;
 reg [C_PROBE354_WIDTH-1:0]mem_shift_probe354  ;
 reg [C_PROBE355_WIDTH-1:0]mem_shift_probe355  ;
 reg [C_PROBE356_WIDTH-1:0]mem_shift_probe356  ;
 reg [C_PROBE357_WIDTH-1:0]mem_shift_probe357  ;
 reg [C_PROBE358_WIDTH-1:0]mem_shift_probe358  ;
 reg [C_PROBE359_WIDTH-1:0]mem_shift_probe359  ;
 reg [C_PROBE360_WIDTH-1:0]mem_shift_probe360  ;
 reg [C_PROBE361_WIDTH-1:0]mem_shift_probe361  ;
 reg [C_PROBE362_WIDTH-1:0]mem_shift_probe362  ;
 reg [C_PROBE363_WIDTH-1:0]mem_shift_probe363  ;
 reg [C_PROBE364_WIDTH-1:0]mem_shift_probe364  ;
 reg [C_PROBE365_WIDTH-1:0]mem_shift_probe365  ;
 reg [C_PROBE366_WIDTH-1:0]mem_shift_probe366  ;
 reg [C_PROBE367_WIDTH-1:0]mem_shift_probe367  ;
 reg [C_PROBE368_WIDTH-1:0]mem_shift_probe368  ;
 reg [C_PROBE369_WIDTH-1:0]mem_shift_probe369  ;
 reg [C_PROBE370_WIDTH-1:0]mem_shift_probe370  ;
 reg [C_PROBE371_WIDTH-1:0]mem_shift_probe371  ;
 reg [C_PROBE372_WIDTH-1:0]mem_shift_probe372  ;
 reg [C_PROBE373_WIDTH-1:0]mem_shift_probe373  ;
 reg [C_PROBE374_WIDTH-1:0]mem_shift_probe374  ;
 reg [C_PROBE375_WIDTH-1:0]mem_shift_probe375  ;
 reg [C_PROBE376_WIDTH-1:0]mem_shift_probe376  ;
 reg [C_PROBE377_WIDTH-1:0]mem_shift_probe377  ;
 reg [C_PROBE378_WIDTH-1:0]mem_shift_probe378  ;
 reg [C_PROBE379_WIDTH-1:0]mem_shift_probe379  ;
 reg [C_PROBE380_WIDTH-1:0]mem_shift_probe380  ;
 reg [C_PROBE381_WIDTH-1:0]mem_shift_probe381  ;
 reg [C_PROBE382_WIDTH-1:0]mem_shift_probe382  ;
 reg [C_PROBE383_WIDTH-1:0]mem_shift_probe383  ;
 reg [C_PROBE384_WIDTH-1:0]mem_shift_probe384  ;
 reg [C_PROBE385_WIDTH-1:0]mem_shift_probe385  ;
 reg [C_PROBE386_WIDTH-1:0]mem_shift_probe386  ;
 reg [C_PROBE387_WIDTH-1:0]mem_shift_probe387  ;
 reg [C_PROBE388_WIDTH-1:0]mem_shift_probe388  ;
 reg [C_PROBE389_WIDTH-1:0]mem_shift_probe389  ;
 reg [C_PROBE390_WIDTH-1:0]mem_shift_probe390  ;
 reg [C_PROBE391_WIDTH-1:0]mem_shift_probe391  ;
 reg [C_PROBE392_WIDTH-1:0]mem_shift_probe392  ;
 reg [C_PROBE393_WIDTH-1:0]mem_shift_probe393  ;
 reg [C_PROBE394_WIDTH-1:0]mem_shift_probe394  ;
 reg [C_PROBE395_WIDTH-1:0]mem_shift_probe395  ;
 reg [C_PROBE396_WIDTH-1:0]mem_shift_probe396  ;
 reg [C_PROBE397_WIDTH-1:0]mem_shift_probe397  ;
 reg [C_PROBE398_WIDTH-1:0]mem_shift_probe398  ;
 reg [C_PROBE399_WIDTH-1:0]mem_shift_probe399  ;
 reg [C_PROBE400_WIDTH-1:0]mem_shift_probe400  ;
 reg [C_PROBE401_WIDTH-1:0]mem_shift_probe401  ;
 reg [C_PROBE402_WIDTH-1:0]mem_shift_probe402  ;
 reg [C_PROBE403_WIDTH-1:0]mem_shift_probe403  ;
 reg [C_PROBE404_WIDTH-1:0]mem_shift_probe404  ;
 reg [C_PROBE405_WIDTH-1:0]mem_shift_probe405  ;
 reg [C_PROBE406_WIDTH-1:0]mem_shift_probe406  ;
 reg [C_PROBE407_WIDTH-1:0]mem_shift_probe407  ;
 reg [C_PROBE408_WIDTH-1:0]mem_shift_probe408  ;
 reg [C_PROBE409_WIDTH-1:0]mem_shift_probe409  ;
 reg [C_PROBE410_WIDTH-1:0]mem_shift_probe410  ;
 reg [C_PROBE411_WIDTH-1:0]mem_shift_probe411  ;
 reg [C_PROBE412_WIDTH-1:0]mem_shift_probe412  ;
 reg [C_PROBE413_WIDTH-1:0]mem_shift_probe413  ;
 reg [C_PROBE414_WIDTH-1:0]mem_shift_probe414  ;
 reg [C_PROBE415_WIDTH-1:0]mem_shift_probe415  ;
 reg [C_PROBE416_WIDTH-1:0]mem_shift_probe416  ;
 reg [C_PROBE417_WIDTH-1:0]mem_shift_probe417  ;
 reg [C_PROBE418_WIDTH-1:0]mem_shift_probe418  ;
 reg [C_PROBE419_WIDTH-1:0]mem_shift_probe419  ;
 reg [C_PROBE420_WIDTH-1:0]mem_shift_probe420  ;
 reg [C_PROBE421_WIDTH-1:0]mem_shift_probe421  ;
 reg [C_PROBE422_WIDTH-1:0]mem_shift_probe422  ;
 reg [C_PROBE423_WIDTH-1:0]mem_shift_probe423  ;
 reg [C_PROBE424_WIDTH-1:0]mem_shift_probe424  ;
 reg [C_PROBE425_WIDTH-1:0]mem_shift_probe425  ;
 reg [C_PROBE426_WIDTH-1:0]mem_shift_probe426  ;
 reg [C_PROBE427_WIDTH-1:0]mem_shift_probe427  ;
 reg [C_PROBE428_WIDTH-1:0]mem_shift_probe428  ;
 reg [C_PROBE429_WIDTH-1:0]mem_shift_probe429  ;
 reg [C_PROBE430_WIDTH-1:0]mem_shift_probe430  ;
 reg [C_PROBE431_WIDTH-1:0]mem_shift_probe431  ;
 reg [C_PROBE432_WIDTH-1:0]mem_shift_probe432  ;
 reg [C_PROBE433_WIDTH-1:0]mem_shift_probe433  ;
 reg [C_PROBE434_WIDTH-1:0]mem_shift_probe434  ;
 reg [C_PROBE435_WIDTH-1:0]mem_shift_probe435  ;
 reg [C_PROBE436_WIDTH-1:0]mem_shift_probe436  ;
 reg [C_PROBE437_WIDTH-1:0]mem_shift_probe437  ;
 reg [C_PROBE438_WIDTH-1:0]mem_shift_probe438  ;
 reg [C_PROBE439_WIDTH-1:0]mem_shift_probe439  ;
 reg [C_PROBE440_WIDTH-1:0]mem_shift_probe440  ;
 reg [C_PROBE441_WIDTH-1:0]mem_shift_probe441  ;
 reg [C_PROBE442_WIDTH-1:0]mem_shift_probe442  ;
 reg [C_PROBE443_WIDTH-1:0]mem_shift_probe443  ;
 reg [C_PROBE444_WIDTH-1:0]mem_shift_probe444  ;
 reg [C_PROBE445_WIDTH-1:0]mem_shift_probe445  ;
 reg [C_PROBE446_WIDTH-1:0]mem_shift_probe446  ;
 reg [C_PROBE447_WIDTH-1:0]mem_shift_probe447  ;
 reg [C_PROBE448_WIDTH-1:0]mem_shift_probe448  ;
 reg [C_PROBE449_WIDTH-1:0]mem_shift_probe449  ;
 reg [C_PROBE450_WIDTH-1:0]mem_shift_probe450  ;
 reg [C_PROBE451_WIDTH-1:0]mem_shift_probe451  ;
 reg [C_PROBE452_WIDTH-1:0]mem_shift_probe452  ;
 reg [C_PROBE453_WIDTH-1:0]mem_shift_probe453  ;
 reg [C_PROBE454_WIDTH-1:0]mem_shift_probe454  ;
 reg [C_PROBE455_WIDTH-1:0]mem_shift_probe455  ;
 reg [C_PROBE456_WIDTH-1:0]mem_shift_probe456  ;
 reg [C_PROBE457_WIDTH-1:0]mem_shift_probe457  ;
 reg [C_PROBE458_WIDTH-1:0]mem_shift_probe458  ;
 reg [C_PROBE459_WIDTH-1:0]mem_shift_probe459  ;
 reg [C_PROBE460_WIDTH-1:0]mem_shift_probe460  ;
 reg [C_PROBE461_WIDTH-1:0]mem_shift_probe461  ;
 reg [C_PROBE462_WIDTH-1:0]mem_shift_probe462  ;
 reg [C_PROBE463_WIDTH-1:0]mem_shift_probe463  ;
 reg [C_PROBE464_WIDTH-1:0]mem_shift_probe464  ;
 reg [C_PROBE465_WIDTH-1:0]mem_shift_probe465  ;
 reg [C_PROBE466_WIDTH-1:0]mem_shift_probe466  ;
 reg [C_PROBE467_WIDTH-1:0]mem_shift_probe467  ;
 reg [C_PROBE468_WIDTH-1:0]mem_shift_probe468  ;
 reg [C_PROBE469_WIDTH-1:0]mem_shift_probe469  ;
 reg [C_PROBE470_WIDTH-1:0]mem_shift_probe470  ;
 reg [C_PROBE471_WIDTH-1:0]mem_shift_probe471  ;
 reg [C_PROBE472_WIDTH-1:0]mem_shift_probe472  ;
 reg [C_PROBE473_WIDTH-1:0]mem_shift_probe473  ;
 reg [C_PROBE474_WIDTH-1:0]mem_shift_probe474  ;
 reg [C_PROBE475_WIDTH-1:0]mem_shift_probe475  ;
 reg [C_PROBE476_WIDTH-1:0]mem_shift_probe476  ;
 reg [C_PROBE477_WIDTH-1:0]mem_shift_probe477  ;
 reg [C_PROBE478_WIDTH-1:0]mem_shift_probe478  ;
 reg [C_PROBE479_WIDTH-1:0]mem_shift_probe479  ;
 reg [C_PROBE480_WIDTH-1:0]mem_shift_probe480  ;
 reg [C_PROBE481_WIDTH-1:0]mem_shift_probe481  ;
 reg [C_PROBE482_WIDTH-1:0]mem_shift_probe482  ;
 reg [C_PROBE483_WIDTH-1:0]mem_shift_probe483  ;
 reg [C_PROBE484_WIDTH-1:0]mem_shift_probe484  ;
 reg [C_PROBE485_WIDTH-1:0]mem_shift_probe485  ;
 reg [C_PROBE486_WIDTH-1:0]mem_shift_probe486  ;
 reg [C_PROBE487_WIDTH-1:0]mem_shift_probe487  ;
 reg [C_PROBE488_WIDTH-1:0]mem_shift_probe488  ;
 reg [C_PROBE489_WIDTH-1:0]mem_shift_probe489  ;
 reg [C_PROBE490_WIDTH-1:0]mem_shift_probe490  ;
 reg [C_PROBE491_WIDTH-1:0]mem_shift_probe491  ;
 reg [C_PROBE492_WIDTH-1:0]mem_shift_probe492  ;
 reg [C_PROBE493_WIDTH-1:0]mem_shift_probe493  ;
 reg [C_PROBE494_WIDTH-1:0]mem_shift_probe494  ;
 reg [C_PROBE495_WIDTH-1:0]mem_shift_probe495  ;
 reg [C_PROBE496_WIDTH-1:0]mem_shift_probe496  ;
 reg [C_PROBE497_WIDTH-1:0]mem_shift_probe497  ;
 reg [C_PROBE498_WIDTH-1:0]mem_shift_probe498  ;
 reg [C_PROBE499_WIDTH-1:0]mem_shift_probe499  ;
 reg [C_PROBE500_WIDTH-1:0]mem_shift_probe500  ;
 reg [C_PROBE501_WIDTH-1:0]mem_shift_probe501  ;
 reg [C_PROBE502_WIDTH-1:0]mem_shift_probe502  ;
 reg [C_PROBE503_WIDTH-1:0]mem_shift_probe503  ;
 reg [C_PROBE504_WIDTH-1:0]mem_shift_probe504  ;
 reg [C_PROBE505_WIDTH-1:0]mem_shift_probe505  ;
 reg [C_PROBE506_WIDTH-1:0]mem_shift_probe506  ;
 reg [C_PROBE507_WIDTH-1:0]mem_shift_probe507  ;
 reg [C_PROBE508_WIDTH-1:0]mem_shift_probe508  ;
 reg [C_PROBE509_WIDTH-1:0]mem_shift_probe509  ;
 reg [C_PROBE510_WIDTH-1:0]mem_shift_probe510  ;
 reg [C_PROBE511_WIDTH-1:0]mem_shift_probe511  ;

 reg [C_PROBE0_WIDTH-1:0]  shift_probe0;
 reg [C_PROBE1_WIDTH-1:0]  shift_probe1;
 reg [C_PROBE2_WIDTH-1:0]  shift_probe2;
 reg [C_PROBE3_WIDTH-1:0]  shift_probe3;
 reg [C_PROBE4_WIDTH-1:0]  shift_probe4;
 reg [C_PROBE5_WIDTH-1:0]  shift_probe5;
 reg [C_PROBE6_WIDTH-1:0]  shift_probe6;
 reg [C_PROBE7_WIDTH-1:0]  shift_probe7;
 reg [C_PROBE8_WIDTH-1:0]  shift_probe8;
 reg [C_PROBE9_WIDTH-1:0]  shift_probe9;
 reg [C_PROBE10_WIDTH-1:0] shift_probe10  ;
 reg [C_PROBE11_WIDTH-1:0] shift_probe11  ;
 reg [C_PROBE12_WIDTH-1:0] shift_probe12  ;
 reg [C_PROBE13_WIDTH-1:0] shift_probe13  ;
 reg [C_PROBE14_WIDTH-1:0] shift_probe14  ;
 reg [C_PROBE15_WIDTH-1:0] shift_probe15  ;
 reg [C_PROBE16_WIDTH-1:0] shift_probe16  ;
 reg [C_PROBE17_WIDTH-1:0] shift_probe17  ;
 reg [C_PROBE18_WIDTH-1:0] shift_probe18  ;
 reg [C_PROBE19_WIDTH-1:0] shift_probe19  ;
 reg [C_PROBE20_WIDTH-1:0] shift_probe20  ;
 reg [C_PROBE21_WIDTH-1:0] shift_probe21  ;
 reg [C_PROBE22_WIDTH-1:0] shift_probe22  ;
 reg [C_PROBE23_WIDTH-1:0] shift_probe23  ;
 reg [C_PROBE24_WIDTH-1:0] shift_probe24  ;
 reg [C_PROBE25_WIDTH-1:0] shift_probe25  ;
 reg [C_PROBE26_WIDTH-1:0] shift_probe26  ;
 reg [C_PROBE27_WIDTH-1:0] shift_probe27  ;
 reg [C_PROBE28_WIDTH-1:0] shift_probe28  ;
 reg [C_PROBE29_WIDTH-1:0] shift_probe29  ;
 reg [C_PROBE30_WIDTH-1:0] shift_probe30  ;
 reg [C_PROBE31_WIDTH-1:0] shift_probe31  ;
 reg [C_PROBE32_WIDTH-1:0] shift_probe32  ;
 reg [C_PROBE33_WIDTH-1:0] shift_probe33  ;
 reg [C_PROBE34_WIDTH-1:0] shift_probe34  ;
 reg [C_PROBE35_WIDTH-1:0] shift_probe35  ;
 reg [C_PROBE36_WIDTH-1:0] shift_probe36  ;
 reg [C_PROBE37_WIDTH-1:0] shift_probe37  ;
 reg [C_PROBE38_WIDTH-1:0] shift_probe38  ;
 reg [C_PROBE39_WIDTH-1:0] shift_probe39  ;
 reg [C_PROBE40_WIDTH-1:0] shift_probe40  ;
 reg [C_PROBE41_WIDTH-1:0] shift_probe41  ;
 reg [C_PROBE42_WIDTH-1:0] shift_probe42  ;
 reg [C_PROBE43_WIDTH-1:0] shift_probe43  ;
 reg [C_PROBE44_WIDTH-1:0] shift_probe44  ;
 reg [C_PROBE45_WIDTH-1:0] shift_probe45  ;
 reg [C_PROBE46_WIDTH-1:0] shift_probe46  ;
 reg [C_PROBE47_WIDTH-1:0] shift_probe47  ;
 reg [C_PROBE48_WIDTH-1:0] shift_probe48  ;
 reg [C_PROBE49_WIDTH-1:0] shift_probe49  ;
 reg [C_PROBE50_WIDTH-1:0] shift_probe50  ;
 reg [C_PROBE51_WIDTH-1:0] shift_probe51  ;
 reg [C_PROBE52_WIDTH-1:0] shift_probe52  ;
 reg [C_PROBE53_WIDTH-1:0] shift_probe53  ;
 reg [C_PROBE54_WIDTH-1:0] shift_probe54  ;
 reg [C_PROBE55_WIDTH-1:0] shift_probe55  ;
 reg [C_PROBE56_WIDTH-1:0] shift_probe56  ;
 reg [C_PROBE57_WIDTH-1:0] shift_probe57  ;
 reg [C_PROBE58_WIDTH-1:0] shift_probe58  ;
 reg [C_PROBE59_WIDTH-1:0] shift_probe59  ;
 reg [C_PROBE60_WIDTH-1:0] shift_probe60  ;
 reg [C_PROBE61_WIDTH-1:0] shift_probe61  ;
 reg [C_PROBE62_WIDTH-1:0] shift_probe62  ;
 reg [C_PROBE63_WIDTH-1:0] shift_probe63  ;
 reg [C_PROBE64_WIDTH-1:0] shift_probe64  ;
 reg [C_PROBE65_WIDTH-1:0] shift_probe65  ;
 reg [C_PROBE66_WIDTH-1:0] shift_probe66  ;
 reg [C_PROBE67_WIDTH-1:0] shift_probe67  ;
 reg [C_PROBE68_WIDTH-1:0] shift_probe68  ;
 reg [C_PROBE69_WIDTH-1:0] shift_probe69  ;
 reg [C_PROBE70_WIDTH-1:0] shift_probe70  ;
 reg [C_PROBE71_WIDTH-1:0] shift_probe71  ;
 reg [C_PROBE72_WIDTH-1:0] shift_probe72  ;
 reg [C_PROBE73_WIDTH-1:0] shift_probe73  ;
 reg [C_PROBE74_WIDTH-1:0] shift_probe74  ;
 reg [C_PROBE75_WIDTH-1:0] shift_probe75  ;
 reg [C_PROBE76_WIDTH-1:0] shift_probe76  ;
 reg [C_PROBE77_WIDTH-1:0] shift_probe77  ;
 reg [C_PROBE78_WIDTH-1:0] shift_probe78  ;
 reg [C_PROBE79_WIDTH-1:0] shift_probe79  ;
 reg [C_PROBE80_WIDTH-1:0] shift_probe80  ;
 reg [C_PROBE81_WIDTH-1:0] shift_probe81  ;
 reg [C_PROBE82_WIDTH-1:0] shift_probe82  ;
 reg [C_PROBE83_WIDTH-1:0] shift_probe83  ;
 reg [C_PROBE84_WIDTH-1:0] shift_probe84  ;
 reg [C_PROBE85_WIDTH-1:0] shift_probe85  ;
 reg [C_PROBE86_WIDTH-1:0] shift_probe86  ;
 reg [C_PROBE87_WIDTH-1:0] shift_probe87  ;
 reg [C_PROBE88_WIDTH-1:0] shift_probe88  ;
 reg [C_PROBE89_WIDTH-1:0] shift_probe89  ;
 reg [C_PROBE90_WIDTH-1:0] shift_probe90  ;
 reg [C_PROBE91_WIDTH-1:0] shift_probe91  ;
 reg [C_PROBE92_WIDTH-1:0] shift_probe92  ;
 reg [C_PROBE93_WIDTH-1:0] shift_probe93  ;
 reg [C_PROBE94_WIDTH-1:0] shift_probe94  ;
 reg [C_PROBE95_WIDTH-1:0] shift_probe95  ;
 reg [C_PROBE96_WIDTH-1:0] shift_probe96  ;
 reg [C_PROBE97_WIDTH-1:0] shift_probe97  ;
 reg [C_PROBE98_WIDTH-1:0] shift_probe98  ;
 reg [C_PROBE99_WIDTH-1:0] shift_probe99  ;
 reg [C_PROBE100_WIDTH-1:0]shift_probe100  ;
 reg [C_PROBE101_WIDTH-1:0]shift_probe101  ;
 reg [C_PROBE102_WIDTH-1:0]shift_probe102  ;
 reg [C_PROBE103_WIDTH-1:0]shift_probe103  ;
 reg [C_PROBE104_WIDTH-1:0]shift_probe104  ;
 reg [C_PROBE105_WIDTH-1:0]shift_probe105  ;
 reg [C_PROBE106_WIDTH-1:0]shift_probe106  ;
 reg [C_PROBE107_WIDTH-1:0]shift_probe107  ;
 reg [C_PROBE108_WIDTH-1:0]shift_probe108  ;
 reg [C_PROBE109_WIDTH-1:0]shift_probe109  ;
 reg [C_PROBE110_WIDTH-1:0]shift_probe110  ;
 reg [C_PROBE111_WIDTH-1:0]shift_probe111  ;
 reg [C_PROBE112_WIDTH-1:0]shift_probe112  ;
 reg [C_PROBE113_WIDTH-1:0]shift_probe113  ;
 reg [C_PROBE114_WIDTH-1:0]shift_probe114  ;
 reg [C_PROBE115_WIDTH-1:0]shift_probe115  ;
 reg [C_PROBE116_WIDTH-1:0]shift_probe116  ;
 reg [C_PROBE117_WIDTH-1:0]shift_probe117  ;
 reg [C_PROBE118_WIDTH-1:0]shift_probe118  ;
 reg [C_PROBE119_WIDTH-1:0]shift_probe119  ;
 reg [C_PROBE120_WIDTH-1:0]shift_probe120  ;
 reg [C_PROBE121_WIDTH-1:0]shift_probe121  ;
 reg [C_PROBE122_WIDTH-1:0]shift_probe122  ;
 reg [C_PROBE123_WIDTH-1:0]shift_probe123  ;
 reg [C_PROBE124_WIDTH-1:0]shift_probe124  ;
 reg [C_PROBE125_WIDTH-1:0]shift_probe125  ;
 reg [C_PROBE126_WIDTH-1:0]shift_probe126  ;
 reg [C_PROBE127_WIDTH-1:0]shift_probe127  ;
 reg [C_PROBE128_WIDTH-1:0]shift_probe128  ;
 reg [C_PROBE129_WIDTH-1:0]shift_probe129  ;
 reg [C_PROBE130_WIDTH-1:0]shift_probe130  ;
 reg [C_PROBE131_WIDTH-1:0]shift_probe131  ;
 reg [C_PROBE132_WIDTH-1:0]shift_probe132  ;
 reg [C_PROBE133_WIDTH-1:0]shift_probe133  ;
 reg [C_PROBE134_WIDTH-1:0]shift_probe134  ;
 reg [C_PROBE135_WIDTH-1:0]shift_probe135  ;
 reg [C_PROBE136_WIDTH-1:0]shift_probe136  ;
 reg [C_PROBE137_WIDTH-1:0]shift_probe137  ;
 reg [C_PROBE138_WIDTH-1:0]shift_probe138  ;
 reg [C_PROBE139_WIDTH-1:0]shift_probe139  ;
 reg [C_PROBE140_WIDTH-1:0]shift_probe140  ;
 reg [C_PROBE141_WIDTH-1:0]shift_probe141  ;
 reg [C_PROBE142_WIDTH-1:0]shift_probe142  ;
 reg [C_PROBE143_WIDTH-1:0]shift_probe143  ;
 reg [C_PROBE144_WIDTH-1:0]shift_probe144  ;
 reg [C_PROBE145_WIDTH-1:0]shift_probe145  ;
 reg [C_PROBE146_WIDTH-1:0]shift_probe146  ;
 reg [C_PROBE147_WIDTH-1:0]shift_probe147  ;
 reg [C_PROBE148_WIDTH-1:0]shift_probe148  ;
 reg [C_PROBE149_WIDTH-1:0]shift_probe149  ;
 reg [C_PROBE150_WIDTH-1:0]shift_probe150  ;
 reg [C_PROBE151_WIDTH-1:0]shift_probe151  ;
 reg [C_PROBE152_WIDTH-1:0]shift_probe152  ;
 reg [C_PROBE153_WIDTH-1:0]shift_probe153  ;
 reg [C_PROBE154_WIDTH-1:0]shift_probe154  ;
 reg [C_PROBE155_WIDTH-1:0]shift_probe155  ;
 reg [C_PROBE156_WIDTH-1:0]shift_probe156  ;
 reg [C_PROBE157_WIDTH-1:0]shift_probe157  ;
 reg [C_PROBE158_WIDTH-1:0]shift_probe158  ;
 reg [C_PROBE159_WIDTH-1:0]shift_probe159  ;
 reg [C_PROBE160_WIDTH-1:0]shift_probe160  ;
 reg [C_PROBE161_WIDTH-1:0]shift_probe161  ;
 reg [C_PROBE162_WIDTH-1:0]shift_probe162  ;
 reg [C_PROBE163_WIDTH-1:0]shift_probe163  ;
 reg [C_PROBE164_WIDTH-1:0]shift_probe164  ;
 reg [C_PROBE165_WIDTH-1:0]shift_probe165  ;
 reg [C_PROBE166_WIDTH-1:0]shift_probe166  ;
 reg [C_PROBE167_WIDTH-1:0]shift_probe167  ;
 reg [C_PROBE168_WIDTH-1:0]shift_probe168  ;
 reg [C_PROBE169_WIDTH-1:0]shift_probe169  ;
 reg [C_PROBE170_WIDTH-1:0]shift_probe170  ;
 reg [C_PROBE171_WIDTH-1:0]shift_probe171  ;
 reg [C_PROBE172_WIDTH-1:0]shift_probe172  ;
 reg [C_PROBE173_WIDTH-1:0]shift_probe173  ;
 reg [C_PROBE174_WIDTH-1:0]shift_probe174  ;
 reg [C_PROBE175_WIDTH-1:0]shift_probe175  ;
 reg [C_PROBE176_WIDTH-1:0]shift_probe176  ;
 reg [C_PROBE177_WIDTH-1:0]shift_probe177  ;
 reg [C_PROBE178_WIDTH-1:0]shift_probe178  ;
 reg [C_PROBE179_WIDTH-1:0]shift_probe179  ;
 reg [C_PROBE180_WIDTH-1:0]shift_probe180  ;
 reg [C_PROBE181_WIDTH-1:0]shift_probe181  ;
 reg [C_PROBE182_WIDTH-1:0]shift_probe182  ;
 reg [C_PROBE183_WIDTH-1:0]shift_probe183  ;
 reg [C_PROBE184_WIDTH-1:0]shift_probe184  ;
 reg [C_PROBE185_WIDTH-1:0]shift_probe185  ;
 reg [C_PROBE186_WIDTH-1:0]shift_probe186  ;
 reg [C_PROBE187_WIDTH-1:0]shift_probe187  ;
 reg [C_PROBE188_WIDTH-1:0]shift_probe188  ;
 reg [C_PROBE189_WIDTH-1:0]shift_probe189  ;
 reg [C_PROBE190_WIDTH-1:0]shift_probe190  ;
 reg [C_PROBE191_WIDTH-1:0]shift_probe191  ;
 reg [C_PROBE192_WIDTH-1:0]shift_probe192  ;
 reg [C_PROBE193_WIDTH-1:0]shift_probe193  ;
 reg [C_PROBE194_WIDTH-1:0]shift_probe194  ;
 reg [C_PROBE195_WIDTH-1:0]shift_probe195  ;
 reg [C_PROBE196_WIDTH-1:0]shift_probe196  ;
 reg [C_PROBE197_WIDTH-1:0]shift_probe197  ;
 reg [C_PROBE198_WIDTH-1:0]shift_probe198  ;
 reg [C_PROBE199_WIDTH-1:0]shift_probe199  ;
 reg [C_PROBE200_WIDTH-1:0]shift_probe200  ;
 reg [C_PROBE201_WIDTH-1:0]shift_probe201  ;
 reg [C_PROBE202_WIDTH-1:0]shift_probe202  ;
 reg [C_PROBE203_WIDTH-1:0]shift_probe203  ;
 reg [C_PROBE204_WIDTH-1:0]shift_probe204  ;
 reg [C_PROBE205_WIDTH-1:0]shift_probe205  ;
 reg [C_PROBE206_WIDTH-1:0]shift_probe206  ;
 reg [C_PROBE207_WIDTH-1:0]shift_probe207  ;
 reg [C_PROBE208_WIDTH-1:0]shift_probe208  ;
 reg [C_PROBE209_WIDTH-1:0]shift_probe209  ;
 reg [C_PROBE210_WIDTH-1:0]shift_probe210  ;
 reg [C_PROBE211_WIDTH-1:0]shift_probe211  ;
 reg [C_PROBE212_WIDTH-1:0]shift_probe212  ;
 reg [C_PROBE213_WIDTH-1:0]shift_probe213  ;
 reg [C_PROBE214_WIDTH-1:0]shift_probe214  ;
 reg [C_PROBE215_WIDTH-1:0]shift_probe215  ;
 reg [C_PROBE216_WIDTH-1:0]shift_probe216  ;
 reg [C_PROBE217_WIDTH-1:0]shift_probe217  ;
 reg [C_PROBE218_WIDTH-1:0]shift_probe218  ;
 reg [C_PROBE219_WIDTH-1:0]shift_probe219  ;
 reg [C_PROBE220_WIDTH-1:0]shift_probe220  ;
 reg [C_PROBE221_WIDTH-1:0]shift_probe221  ;
 reg [C_PROBE222_WIDTH-1:0]shift_probe222  ;
 reg [C_PROBE223_WIDTH-1:0]shift_probe223  ;
 reg [C_PROBE224_WIDTH-1:0]shift_probe224  ;
 reg [C_PROBE225_WIDTH-1:0]shift_probe225  ;
 reg [C_PROBE226_WIDTH-1:0]shift_probe226  ;
 reg [C_PROBE227_WIDTH-1:0]shift_probe227  ;
 reg [C_PROBE228_WIDTH-1:0]shift_probe228  ;
 reg [C_PROBE229_WIDTH-1:0]shift_probe229  ;
 reg [C_PROBE230_WIDTH-1:0]shift_probe230  ;
 reg [C_PROBE231_WIDTH-1:0]shift_probe231  ;
 reg [C_PROBE232_WIDTH-1:0]shift_probe232  ;
 reg [C_PROBE233_WIDTH-1:0]shift_probe233  ;
 reg [C_PROBE234_WIDTH-1:0]shift_probe234  ;
 reg [C_PROBE235_WIDTH-1:0]shift_probe235  ;
 reg [C_PROBE236_WIDTH-1:0]shift_probe236  ;
 reg [C_PROBE237_WIDTH-1:0]shift_probe237  ;
 reg [C_PROBE238_WIDTH-1:0]shift_probe238  ;
 reg [C_PROBE239_WIDTH-1:0]shift_probe239  ;
 reg [C_PROBE240_WIDTH-1:0]shift_probe240  ;
 reg [C_PROBE241_WIDTH-1:0]shift_probe241  ;
 reg [C_PROBE242_WIDTH-1:0]shift_probe242  ;
 reg [C_PROBE243_WIDTH-1:0]shift_probe243  ;
 reg [C_PROBE244_WIDTH-1:0]shift_probe244  ;
 reg [C_PROBE245_WIDTH-1:0]shift_probe245  ;
 reg [C_PROBE246_WIDTH-1:0]shift_probe246  ;
 reg [C_PROBE247_WIDTH-1:0]shift_probe247  ;
 reg [C_PROBE248_WIDTH-1:0]shift_probe248  ;
 reg [C_PROBE249_WIDTH-1:0]shift_probe249  ;
 reg [C_PROBE250_WIDTH-1:0]shift_probe250  ;
 reg [C_PROBE251_WIDTH-1:0]shift_probe251  ;
 reg [C_PROBE252_WIDTH-1:0]shift_probe252  ;
 reg [C_PROBE253_WIDTH-1:0]shift_probe253  ;
 reg [C_PROBE254_WIDTH-1:0]shift_probe254  ;
 reg [C_PROBE255_WIDTH-1:0]shift_probe255  ;
 reg [C_PROBE256_WIDTH-1:0]shift_probe256  ;
 reg [C_PROBE257_WIDTH-1:0]shift_probe257  ;
 reg [C_PROBE258_WIDTH-1:0]shift_probe258  ;
 reg [C_PROBE259_WIDTH-1:0]shift_probe259  ;
 reg [C_PROBE260_WIDTH-1:0]shift_probe260  ;
 reg [C_PROBE261_WIDTH-1:0]shift_probe261  ;
 reg [C_PROBE262_WIDTH-1:0]shift_probe262  ;
 reg [C_PROBE263_WIDTH-1:0]shift_probe263  ;
 reg [C_PROBE264_WIDTH-1:0]shift_probe264  ;
 reg [C_PROBE265_WIDTH-1:0]shift_probe265  ;
 reg [C_PROBE266_WIDTH-1:0]shift_probe266  ;
 reg [C_PROBE267_WIDTH-1:0]shift_probe267  ;
 reg [C_PROBE268_WIDTH-1:0]shift_probe268  ;
 reg [C_PROBE269_WIDTH-1:0]shift_probe269  ;
 reg [C_PROBE270_WIDTH-1:0]shift_probe270  ;
 reg [C_PROBE271_WIDTH-1:0]shift_probe271  ;
 reg [C_PROBE272_WIDTH-1:0]shift_probe272  ;
 reg [C_PROBE273_WIDTH-1:0]shift_probe273  ;
 reg [C_PROBE274_WIDTH-1:0]shift_probe274  ;
 reg [C_PROBE275_WIDTH-1:0]shift_probe275  ;
 reg [C_PROBE276_WIDTH-1:0]shift_probe276  ;
 reg [C_PROBE277_WIDTH-1:0]shift_probe277  ;
 reg [C_PROBE278_WIDTH-1:0]shift_probe278  ;
 reg [C_PROBE279_WIDTH-1:0]shift_probe279  ;
 reg [C_PROBE280_WIDTH-1:0]shift_probe280  ;
 reg [C_PROBE281_WIDTH-1:0]shift_probe281  ;
 reg [C_PROBE282_WIDTH-1:0]shift_probe282  ;
 reg [C_PROBE283_WIDTH-1:0]shift_probe283  ;
 reg [C_PROBE284_WIDTH-1:0]shift_probe284  ;
 reg [C_PROBE285_WIDTH-1:0]shift_probe285  ;
 reg [C_PROBE286_WIDTH-1:0]shift_probe286  ;
 reg [C_PROBE287_WIDTH-1:0]shift_probe287  ;
 reg [C_PROBE288_WIDTH-1:0]shift_probe288  ;
 reg [C_PROBE289_WIDTH-1:0]shift_probe289  ;
 reg [C_PROBE290_WIDTH-1:0]shift_probe290  ;
 reg [C_PROBE291_WIDTH-1:0]shift_probe291  ;
 reg [C_PROBE292_WIDTH-1:0]shift_probe292  ;
 reg [C_PROBE293_WIDTH-1:0]shift_probe293  ;
 reg [C_PROBE294_WIDTH-1:0]shift_probe294  ;
 reg [C_PROBE295_WIDTH-1:0]shift_probe295  ;
 reg [C_PROBE296_WIDTH-1:0]shift_probe296  ;
 reg [C_PROBE297_WIDTH-1:0]shift_probe297  ;
 reg [C_PROBE298_WIDTH-1:0]shift_probe298  ;
 reg [C_PROBE299_WIDTH-1:0]shift_probe299  ;
 reg [C_PROBE300_WIDTH-1:0]shift_probe300  ;
 reg [C_PROBE301_WIDTH-1:0]shift_probe301  ;
 reg [C_PROBE302_WIDTH-1:0]shift_probe302  ;
 reg [C_PROBE303_WIDTH-1:0]shift_probe303  ;
 reg [C_PROBE304_WIDTH-1:0]shift_probe304  ;
 reg [C_PROBE305_WIDTH-1:0]shift_probe305  ;
 reg [C_PROBE306_WIDTH-1:0]shift_probe306  ;
 reg [C_PROBE307_WIDTH-1:0]shift_probe307  ;
 reg [C_PROBE308_WIDTH-1:0]shift_probe308  ;
 reg [C_PROBE309_WIDTH-1:0]shift_probe309  ;
 reg [C_PROBE310_WIDTH-1:0]shift_probe310  ;
 reg [C_PROBE311_WIDTH-1:0]shift_probe311  ;
 reg [C_PROBE312_WIDTH-1:0]shift_probe312  ;
 reg [C_PROBE313_WIDTH-1:0]shift_probe313  ;
 reg [C_PROBE314_WIDTH-1:0]shift_probe314  ;
 reg [C_PROBE315_WIDTH-1:0]shift_probe315  ;
 reg [C_PROBE316_WIDTH-1:0]shift_probe316  ;
 reg [C_PROBE317_WIDTH-1:0]shift_probe317  ;
 reg [C_PROBE318_WIDTH-1:0]shift_probe318  ;
 reg [C_PROBE319_WIDTH-1:0]shift_probe319  ;
 reg [C_PROBE320_WIDTH-1:0]shift_probe320  ;
 reg [C_PROBE321_WIDTH-1:0]shift_probe321  ;
 reg [C_PROBE322_WIDTH-1:0]shift_probe322  ;
 reg [C_PROBE323_WIDTH-1:0]shift_probe323  ;
 reg [C_PROBE324_WIDTH-1:0]shift_probe324  ;
 reg [C_PROBE325_WIDTH-1:0]shift_probe325  ;
 reg [C_PROBE326_WIDTH-1:0]shift_probe326  ;
 reg [C_PROBE327_WIDTH-1:0]shift_probe327  ;
 reg [C_PROBE328_WIDTH-1:0]shift_probe328  ;
 reg [C_PROBE329_WIDTH-1:0]shift_probe329  ;
 reg [C_PROBE330_WIDTH-1:0]shift_probe330  ;
 reg [C_PROBE331_WIDTH-1:0]shift_probe331  ;
 reg [C_PROBE332_WIDTH-1:0]shift_probe332  ;
 reg [C_PROBE333_WIDTH-1:0]shift_probe333  ;
 reg [C_PROBE334_WIDTH-1:0]shift_probe334  ;
 reg [C_PROBE335_WIDTH-1:0]shift_probe335  ;
 reg [C_PROBE336_WIDTH-1:0]shift_probe336  ;
 reg [C_PROBE337_WIDTH-1:0]shift_probe337  ;
 reg [C_PROBE338_WIDTH-1:0]shift_probe338  ;
 reg [C_PROBE339_WIDTH-1:0]shift_probe339  ;
 reg [C_PROBE340_WIDTH-1:0]shift_probe340  ;
 reg [C_PROBE341_WIDTH-1:0]shift_probe341  ;
 reg [C_PROBE342_WIDTH-1:0]shift_probe342  ;
 reg [C_PROBE343_WIDTH-1:0]shift_probe343  ;
 reg [C_PROBE344_WIDTH-1:0]shift_probe344  ;
 reg [C_PROBE345_WIDTH-1:0]shift_probe345  ;
 reg [C_PROBE346_WIDTH-1:0]shift_probe346  ;
 reg [C_PROBE347_WIDTH-1:0]shift_probe347  ;
 reg [C_PROBE348_WIDTH-1:0]shift_probe348  ;
 reg [C_PROBE349_WIDTH-1:0]shift_probe349  ;
 reg [C_PROBE350_WIDTH-1:0]shift_probe350  ;
 reg [C_PROBE351_WIDTH-1:0]shift_probe351  ;
 reg [C_PROBE352_WIDTH-1:0]shift_probe352  ;
 reg [C_PROBE353_WIDTH-1:0]shift_probe353  ;
 reg [C_PROBE354_WIDTH-1:0]shift_probe354  ;
 reg [C_PROBE355_WIDTH-1:0]shift_probe355  ;
 reg [C_PROBE356_WIDTH-1:0]shift_probe356  ;
 reg [C_PROBE357_WIDTH-1:0]shift_probe357  ;
 reg [C_PROBE358_WIDTH-1:0]shift_probe358  ;
 reg [C_PROBE359_WIDTH-1:0]shift_probe359  ;
 reg [C_PROBE360_WIDTH-1:0]shift_probe360  ;
 reg [C_PROBE361_WIDTH-1:0]shift_probe361  ;
 reg [C_PROBE362_WIDTH-1:0]shift_probe362  ;
 reg [C_PROBE363_WIDTH-1:0]shift_probe363  ;
 reg [C_PROBE364_WIDTH-1:0]shift_probe364  ;
 reg [C_PROBE365_WIDTH-1:0]shift_probe365  ;
 reg [C_PROBE366_WIDTH-1:0]shift_probe366  ;
 reg [C_PROBE367_WIDTH-1:0]shift_probe367  ;
 reg [C_PROBE368_WIDTH-1:0]shift_probe368  ;
 reg [C_PROBE369_WIDTH-1:0]shift_probe369  ;
 reg [C_PROBE370_WIDTH-1:0]shift_probe370  ;
 reg [C_PROBE371_WIDTH-1:0]shift_probe371  ;
 reg [C_PROBE372_WIDTH-1:0]shift_probe372  ;
 reg [C_PROBE373_WIDTH-1:0]shift_probe373  ;
 reg [C_PROBE374_WIDTH-1:0]shift_probe374  ;
 reg [C_PROBE375_WIDTH-1:0]shift_probe375  ;
 reg [C_PROBE376_WIDTH-1:0]shift_probe376  ;
 reg [C_PROBE377_WIDTH-1:0]shift_probe377  ;
 reg [C_PROBE378_WIDTH-1:0]shift_probe378  ;
 reg [C_PROBE379_WIDTH-1:0]shift_probe379  ;
 reg [C_PROBE380_WIDTH-1:0]shift_probe380  ;
 reg [C_PROBE381_WIDTH-1:0]shift_probe381  ;
 reg [C_PROBE382_WIDTH-1:0]shift_probe382  ;
 reg [C_PROBE383_WIDTH-1:0]shift_probe383  ;
 reg [C_PROBE384_WIDTH-1:0]shift_probe384  ;
 reg [C_PROBE385_WIDTH-1:0]shift_probe385  ;
 reg [C_PROBE386_WIDTH-1:0]shift_probe386  ;
 reg [C_PROBE387_WIDTH-1:0]shift_probe387  ;
 reg [C_PROBE388_WIDTH-1:0]shift_probe388  ;
 reg [C_PROBE389_WIDTH-1:0]shift_probe389  ;
 reg [C_PROBE390_WIDTH-1:0]shift_probe390  ;
 reg [C_PROBE391_WIDTH-1:0]shift_probe391  ;
 reg [C_PROBE392_WIDTH-1:0]shift_probe392  ;
 reg [C_PROBE393_WIDTH-1:0]shift_probe393  ;
 reg [C_PROBE394_WIDTH-1:0]shift_probe394  ;
 reg [C_PROBE395_WIDTH-1:0]shift_probe395  ;
 reg [C_PROBE396_WIDTH-1:0]shift_probe396  ;
 reg [C_PROBE397_WIDTH-1:0]shift_probe397  ;
 reg [C_PROBE398_WIDTH-1:0]shift_probe398  ;
 reg [C_PROBE399_WIDTH-1:0]shift_probe399  ;
 reg [C_PROBE400_WIDTH-1:0]shift_probe400  ;
 reg [C_PROBE401_WIDTH-1:0]shift_probe401  ;
 reg [C_PROBE402_WIDTH-1:0]shift_probe402  ;
 reg [C_PROBE403_WIDTH-1:0]shift_probe403  ;
 reg [C_PROBE404_WIDTH-1:0]shift_probe404  ;
 reg [C_PROBE405_WIDTH-1:0]shift_probe405  ;
 reg [C_PROBE406_WIDTH-1:0]shift_probe406  ;
 reg [C_PROBE407_WIDTH-1:0]shift_probe407  ;
 reg [C_PROBE408_WIDTH-1:0]shift_probe408  ;
 reg [C_PROBE409_WIDTH-1:0]shift_probe409  ;
 reg [C_PROBE410_WIDTH-1:0]shift_probe410  ;
 reg [C_PROBE411_WIDTH-1:0]shift_probe411  ;
 reg [C_PROBE412_WIDTH-1:0]shift_probe412  ;
 reg [C_PROBE413_WIDTH-1:0]shift_probe413  ;
 reg [C_PROBE414_WIDTH-1:0]shift_probe414  ;
 reg [C_PROBE415_WIDTH-1:0]shift_probe415  ;
 reg [C_PROBE416_WIDTH-1:0]shift_probe416  ;
 reg [C_PROBE417_WIDTH-1:0]shift_probe417  ;
 reg [C_PROBE418_WIDTH-1:0]shift_probe418  ;
 reg [C_PROBE419_WIDTH-1:0]shift_probe419  ;
 reg [C_PROBE420_WIDTH-1:0]shift_probe420  ;
 reg [C_PROBE421_WIDTH-1:0]shift_probe421  ;
 reg [C_PROBE422_WIDTH-1:0]shift_probe422  ;
 reg [C_PROBE423_WIDTH-1:0]shift_probe423  ;
 reg [C_PROBE424_WIDTH-1:0]shift_probe424  ;
 reg [C_PROBE425_WIDTH-1:0]shift_probe425  ;
 reg [C_PROBE426_WIDTH-1:0]shift_probe426  ;
 reg [C_PROBE427_WIDTH-1:0]shift_probe427  ;
 reg [C_PROBE428_WIDTH-1:0]shift_probe428  ;
 reg [C_PROBE429_WIDTH-1:0]shift_probe429  ;
 reg [C_PROBE430_WIDTH-1:0]shift_probe430  ;
 reg [C_PROBE431_WIDTH-1:0]shift_probe431  ;
 reg [C_PROBE432_WIDTH-1:0]shift_probe432  ;
 reg [C_PROBE433_WIDTH-1:0]shift_probe433  ;
 reg [C_PROBE434_WIDTH-1:0]shift_probe434  ;
 reg [C_PROBE435_WIDTH-1:0]shift_probe435  ;
 reg [C_PROBE436_WIDTH-1:0]shift_probe436  ;
 reg [C_PROBE437_WIDTH-1:0]shift_probe437  ;
 reg [C_PROBE438_WIDTH-1:0]shift_probe438  ;
 reg [C_PROBE439_WIDTH-1:0]shift_probe439  ;
 reg [C_PROBE440_WIDTH-1:0]shift_probe440  ;
 reg [C_PROBE441_WIDTH-1:0]shift_probe441  ;
 reg [C_PROBE442_WIDTH-1:0]shift_probe442  ;
 reg [C_PROBE443_WIDTH-1:0]shift_probe443  ;
 reg [C_PROBE444_WIDTH-1:0]shift_probe444  ;
 reg [C_PROBE445_WIDTH-1:0]shift_probe445  ;
 reg [C_PROBE446_WIDTH-1:0]shift_probe446  ;
 reg [C_PROBE447_WIDTH-1:0]shift_probe447  ;
 reg [C_PROBE448_WIDTH-1:0]shift_probe448  ;
 reg [C_PROBE449_WIDTH-1:0]shift_probe449  ;
 reg [C_PROBE450_WIDTH-1:0]shift_probe450  ;
 reg [C_PROBE451_WIDTH-1:0]shift_probe451  ;
 reg [C_PROBE452_WIDTH-1:0]shift_probe452  ;
 reg [C_PROBE453_WIDTH-1:0]shift_probe453  ;
 reg [C_PROBE454_WIDTH-1:0]shift_probe454  ;
 reg [C_PROBE455_WIDTH-1:0]shift_probe455  ;
 reg [C_PROBE456_WIDTH-1:0]shift_probe456  ;
 reg [C_PROBE457_WIDTH-1:0]shift_probe457  ;
 reg [C_PROBE458_WIDTH-1:0]shift_probe458  ;
 reg [C_PROBE459_WIDTH-1:0]shift_probe459  ;
 reg [C_PROBE460_WIDTH-1:0]shift_probe460  ;
 reg [C_PROBE461_WIDTH-1:0]shift_probe461  ;
 reg [C_PROBE462_WIDTH-1:0]shift_probe462  ;
 reg [C_PROBE463_WIDTH-1:0]shift_probe463  ;
 reg [C_PROBE464_WIDTH-1:0]shift_probe464  ;
 reg [C_PROBE465_WIDTH-1:0]shift_probe465  ;
 reg [C_PROBE466_WIDTH-1:0]shift_probe466  ;
 reg [C_PROBE467_WIDTH-1:0]shift_probe467  ;
 reg [C_PROBE468_WIDTH-1:0]shift_probe468  ;
 reg [C_PROBE469_WIDTH-1:0]shift_probe469  ;
 reg [C_PROBE470_WIDTH-1:0]shift_probe470  ;
 reg [C_PROBE471_WIDTH-1:0]shift_probe471  ;
 reg [C_PROBE472_WIDTH-1:0]shift_probe472  ;
 reg [C_PROBE473_WIDTH-1:0]shift_probe473  ;
 reg [C_PROBE474_WIDTH-1:0]shift_probe474  ;
 reg [C_PROBE475_WIDTH-1:0]shift_probe475  ;
 reg [C_PROBE476_WIDTH-1:0]shift_probe476  ;
 reg [C_PROBE477_WIDTH-1:0]shift_probe477  ;
 reg [C_PROBE478_WIDTH-1:0]shift_probe478  ;
 reg [C_PROBE479_WIDTH-1:0]shift_probe479  ;
 reg [C_PROBE480_WIDTH-1:0]shift_probe480  ;
 reg [C_PROBE481_WIDTH-1:0]shift_probe481  ;
 reg [C_PROBE482_WIDTH-1:0]shift_probe482  ;
 reg [C_PROBE483_WIDTH-1:0]shift_probe483  ;
 reg [C_PROBE484_WIDTH-1:0]shift_probe484  ;
 reg [C_PROBE485_WIDTH-1:0]shift_probe485  ;
 reg [C_PROBE486_WIDTH-1:0]shift_probe486  ;
 reg [C_PROBE487_WIDTH-1:0]shift_probe487  ;
 reg [C_PROBE488_WIDTH-1:0]shift_probe488  ;
 reg [C_PROBE489_WIDTH-1:0]shift_probe489  ;
 reg [C_PROBE490_WIDTH-1:0]shift_probe490  ;
 reg [C_PROBE491_WIDTH-1:0]shift_probe491  ;
 reg [C_PROBE492_WIDTH-1:0]shift_probe492  ;
 reg [C_PROBE493_WIDTH-1:0]shift_probe493  ;
 reg [C_PROBE494_WIDTH-1:0]shift_probe494  ;
 reg [C_PROBE495_WIDTH-1:0]shift_probe495  ;
 reg [C_PROBE496_WIDTH-1:0]shift_probe496  ;
 reg [C_PROBE497_WIDTH-1:0]shift_probe497  ;
 reg [C_PROBE498_WIDTH-1:0]shift_probe498  ;
 reg [C_PROBE499_WIDTH-1:0]shift_probe499  ;
 reg [C_PROBE500_WIDTH-1:0]shift_probe500  ;
 reg [C_PROBE501_WIDTH-1:0]shift_probe501  ;
 reg [C_PROBE502_WIDTH-1:0]shift_probe502  ;
 reg [C_PROBE503_WIDTH-1:0]shift_probe503  ;
 reg [C_PROBE504_WIDTH-1:0]shift_probe504  ;
 reg [C_PROBE505_WIDTH-1:0]shift_probe505  ;
 reg [C_PROBE506_WIDTH-1:0]shift_probe506  ;
 reg [C_PROBE507_WIDTH-1:0]shift_probe507  ;
 reg [C_PROBE508_WIDTH-1:0]shift_probe508  ;
 reg [C_PROBE509_WIDTH-1:0]shift_probe509  ;
 reg [C_PROBE510_WIDTH-1:0]shift_probe510  ;
 reg [C_PROBE511_WIDTH-1:0]shift_probe511  ;

generate
  if (C_NUM_PROBES > 0) begin : FF_MEM_PROBE0
    always @ (posedge clk)
    begin
      shift_probe0 <= probe0;
      mem_shift_probe0 <= shift_probe0;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 1) begin : FF_MEM_PROBE1
    always @ (posedge clk)
    begin
      shift_probe1 <= probe1;
      mem_shift_probe1 <= shift_probe1;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 2) begin : FF_MEM_PROBE2
    always @ (posedge clk)
    begin
      shift_probe2 <= probe2;
      mem_shift_probe2 <= shift_probe2;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 3) begin : FF_MEM_PROBE3
    always @ (posedge clk)
    begin
      shift_probe3 <= probe3;
      mem_shift_probe3 <= shift_probe3;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 4) begin : FF_MEM_PROBE4
    always @ (posedge clk)
    begin
      shift_probe4 <= probe4;
      mem_shift_probe4 <= shift_probe4;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 5) begin : FF_MEM_PROBE5
    always @ (posedge clk)
    begin
      shift_probe5 <= probe5;
      mem_shift_probe5 <= shift_probe5;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 6) begin : FF_MEM_PROBE6
    always @ (posedge clk)
    begin
      shift_probe6 <= probe6;
      mem_shift_probe6 <= shift_probe6;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 7) begin : FF_MEM_PROBE7
    always @ (posedge clk)
    begin
      shift_probe7 <= probe7;
      mem_shift_probe7 <= shift_probe7;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 8) begin : FF_MEM_PROBE8
    always @ (posedge clk)
    begin
      shift_probe8 <= probe8;
      mem_shift_probe8 <= shift_probe8;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 9) begin : FF_MEM_PROBE9
    always @ (posedge clk)
    begin
      shift_probe9 <= probe9;
      mem_shift_probe9 <= shift_probe9;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 10) begin : FF_MEM_PROBE10
    always @ (posedge clk)
    begin
      shift_probe10 <= probe10;
      mem_shift_probe10 <= shift_probe10;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 11) begin : FF_MEM_PROBE11
    always @ (posedge clk)
    begin
      shift_probe11 <= probe11;
      mem_shift_probe11 <= shift_probe11;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 12) begin : FF_MEM_PROBE12
    always @ (posedge clk)
    begin
      shift_probe12 <= probe12;
      mem_shift_probe12 <= shift_probe12;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 13) begin : FF_MEM_PROBE13
    always @ (posedge clk)
    begin
      shift_probe13 <= probe13;
      mem_shift_probe13 <= shift_probe13;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 14) begin : FF_MEM_PROBE14
    always @ (posedge clk)
    begin
      shift_probe14 <= probe14;
      mem_shift_probe14 <= shift_probe14;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 15) begin : FF_MEM_PROBE15
    always @ (posedge clk)
    begin
      shift_probe15 <= probe15;
      mem_shift_probe15 <= shift_probe15;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 16) begin : FF_MEM_PROBE16
    always @ (posedge clk)
    begin
      shift_probe16 <= probe16;
      mem_shift_probe16 <= shift_probe16;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 17) begin : FF_MEM_PROBE17
    always @ (posedge clk)
    begin
      shift_probe17 <= probe17;
      mem_shift_probe17 <= shift_probe17;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 18) begin : FF_MEM_PROBE18
    always @ (posedge clk)
    begin
      shift_probe18 <= probe18;
      mem_shift_probe18 <= shift_probe18;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 19) begin : FF_MEM_PROBE19
    always @ (posedge clk)
    begin
      shift_probe19 <= probe19;
      mem_shift_probe19 <= shift_probe19;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 20) begin : FF_MEM_PROBE20
    always @ (posedge clk)
    begin
      shift_probe20 <= probe20;
      mem_shift_probe20 <= shift_probe20;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 21) begin : FF_MEM_PROBE21
    always @ (posedge clk)
    begin
      shift_probe21 <= probe21;
      mem_shift_probe21 <= shift_probe21;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 22) begin : FF_MEM_PROBE22
    always @ (posedge clk)
    begin
      shift_probe22 <= probe22;
      mem_shift_probe22 <= shift_probe22;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 23) begin : FF_MEM_PROBE23
    always @ (posedge clk)
    begin
      shift_probe23 <= probe23;
      mem_shift_probe23 <= shift_probe23;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 24) begin : FF_MEM_PROBE24
    always @ (posedge clk)
    begin
      shift_probe24 <= probe24;
      mem_shift_probe24 <= shift_probe24;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 25) begin : FF_MEM_PROBE25
    always @ (posedge clk)
    begin
      shift_probe25 <= probe25;
      mem_shift_probe25 <= shift_probe25;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 26) begin : FF_MEM_PROBE26
    always @ (posedge clk)
    begin
      shift_probe26 <= probe26;
      mem_shift_probe26 <= shift_probe26;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 27) begin : FF_MEM_PROBE27
    always @ (posedge clk)
    begin
      shift_probe27 <= probe27;
      mem_shift_probe27 <= shift_probe27;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 28) begin : FF_MEM_PROBE28
    always @ (posedge clk)
    begin
      shift_probe28 <= probe28;
      mem_shift_probe28 <= shift_probe28;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 29) begin : FF_MEM_PROBE29
    always @ (posedge clk)
    begin
      shift_probe29 <= probe29;
      mem_shift_probe29 <= shift_probe29;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 30) begin : FF_MEM_PROBE30
    always @ (posedge clk)
    begin
      shift_probe30 <= probe30;
      mem_shift_probe30 <= shift_probe30;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 31) begin : FF_MEM_PROBE31
    always @ (posedge clk)
    begin
      shift_probe31 <= probe31;
      mem_shift_probe31 <= shift_probe31;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 32) begin : FF_MEM_PROBE32
    always @ (posedge clk)
    begin
      shift_probe32 <= probe32;
      mem_shift_probe32 <= shift_probe32;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 33) begin : FF_MEM_PROBE33
    always @ (posedge clk)
    begin
      shift_probe33 <= probe33;
      mem_shift_probe33 <= shift_probe33;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 34) begin : FF_MEM_PROBE34
    always @ (posedge clk)
    begin
      shift_probe34 <= probe34;
      mem_shift_probe34 <= shift_probe34;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 35) begin : FF_MEM_PROBE35
    always @ (posedge clk)
    begin
      shift_probe35 <= probe35;
      mem_shift_probe35 <= shift_probe35;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 36) begin : FF_MEM_PROBE36
    always @ (posedge clk)
    begin
      shift_probe36 <= probe36;
      mem_shift_probe36 <= shift_probe36;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 37) begin : FF_MEM_PROBE37
    always @ (posedge clk)
    begin
      shift_probe37 <= probe37;
      mem_shift_probe37 <= shift_probe37;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 38) begin : FF_MEM_PROBE38
    always @ (posedge clk)
    begin
      shift_probe38 <= probe38;
      mem_shift_probe38 <= shift_probe38;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 39) begin : FF_MEM_PROBE39
    always @ (posedge clk)
    begin
      shift_probe39 <= probe39;
      mem_shift_probe39 <= shift_probe39;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 40) begin : FF_MEM_PROBE40
    always @ (posedge clk)
    begin
      shift_probe40 <= probe40;
      mem_shift_probe40 <= shift_probe40;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 41) begin : FF_MEM_PROBE41
    always @ (posedge clk)
    begin
      shift_probe41 <= probe41;
      mem_shift_probe41 <= shift_probe41;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 42) begin : FF_MEM_PROBE42
    always @ (posedge clk)
    begin
      shift_probe42 <= probe42;
      mem_shift_probe42 <= shift_probe42;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 43) begin : FF_MEM_PROBE43
    always @ (posedge clk)
    begin
      shift_probe43 <= probe43;
      mem_shift_probe43 <= shift_probe43;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 44) begin : FF_MEM_PROBE44
    always @ (posedge clk)
    begin
      shift_probe44 <= probe44;
      mem_shift_probe44 <= shift_probe44;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 45) begin : FF_MEM_PROBE45
    always @ (posedge clk)
    begin
      shift_probe45 <= probe45;
      mem_shift_probe45 <= shift_probe45;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 46) begin : FF_MEM_PROBE46
    always @ (posedge clk)
    begin
      shift_probe46 <= probe46;
      mem_shift_probe46 <= shift_probe46;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 47) begin : FF_MEM_PROBE47
    always @ (posedge clk)
    begin
      shift_probe47 <= probe47;
      mem_shift_probe47 <= shift_probe47;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 48) begin : FF_MEM_PROBE48
    always @ (posedge clk)
    begin
      shift_probe48 <= probe48;
      mem_shift_probe48 <= shift_probe48;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 49) begin : FF_MEM_PROBE49
    always @ (posedge clk)
    begin
      shift_probe49 <= probe49;
      mem_shift_probe49 <= shift_probe49;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 50) begin : FF_MEM_PROBE50
    always @ (posedge clk)
    begin
      shift_probe50 <= probe50;
      mem_shift_probe50 <= shift_probe50;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 51) begin : FF_MEM_PROBE51
    always @ (posedge clk)
    begin
      shift_probe51 <= probe51;
      mem_shift_probe51 <= shift_probe51;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 52) begin : FF_MEM_PROBE52
    always @ (posedge clk)
    begin
      shift_probe52 <= probe52;
      mem_shift_probe52 <= shift_probe52;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 53) begin : FF_MEM_PROBE53
    always @ (posedge clk)
    begin
      shift_probe53 <= probe53;
      mem_shift_probe53 <= shift_probe53;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 54) begin : FF_MEM_PROBE54
    always @ (posedge clk)
    begin
      shift_probe54 <= probe54;
      mem_shift_probe54 <= shift_probe54;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 55) begin : FF_MEM_PROBE55
    always @ (posedge clk)
    begin
      shift_probe55 <= probe55;
      mem_shift_probe55 <= shift_probe55;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 56) begin : FF_MEM_PROBE56
    always @ (posedge clk)
    begin
      shift_probe56 <= probe56;
      mem_shift_probe56 <= shift_probe56;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 57) begin : FF_MEM_PROBE57
    always @ (posedge clk)
    begin
      shift_probe57 <= probe57;
      mem_shift_probe57 <= shift_probe57;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 58) begin : FF_MEM_PROBE58
    always @ (posedge clk)
    begin
      shift_probe58 <= probe58;
      mem_shift_probe58 <= shift_probe58;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 59) begin : FF_MEM_PROBE59
    always @ (posedge clk)
    begin
      shift_probe59 <= probe59;
      mem_shift_probe59 <= shift_probe59;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 60) begin : FF_MEM_PROBE60
    always @ (posedge clk)
    begin
      shift_probe60 <= probe60;
      mem_shift_probe60 <= shift_probe60;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 61) begin : FF_MEM_PROBE61
    always @ (posedge clk)
    begin
      shift_probe61 <= probe61;
      mem_shift_probe61 <= shift_probe61;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 62) begin : FF_MEM_PROBE62
    always @ (posedge clk)
    begin
      shift_probe62 <= probe62;
      mem_shift_probe62 <= shift_probe62;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 63) begin : FF_MEM_PROBE63
    always @ (posedge clk)
    begin
      shift_probe63 <= probe63;
      mem_shift_probe63 <= shift_probe63;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 64) begin : FF_MEM_PROBE64
    always @ (posedge clk)
    begin
      shift_probe64 <= probe64;
      mem_shift_probe64 <= shift_probe64;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 65) begin : FF_MEM_PROBE65
    always @ (posedge clk)
    begin
      shift_probe65 <= probe65;
      mem_shift_probe65 <= shift_probe65;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 66) begin : FF_MEM_PROBE66
    always @ (posedge clk)
    begin
      shift_probe66 <= probe66;
      mem_shift_probe66 <= shift_probe66;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 67) begin : FF_MEM_PROBE67
    always @ (posedge clk)
    begin
      shift_probe67 <= probe67;
      mem_shift_probe67 <= shift_probe67;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 68) begin : FF_MEM_PROBE68
    always @ (posedge clk)
    begin
      shift_probe68 <= probe68;
      mem_shift_probe68 <= shift_probe68;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 69) begin : FF_MEM_PROBE69
    always @ (posedge clk)
    begin
      shift_probe69 <= probe69;
      mem_shift_probe69 <= shift_probe69;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 70) begin : FF_MEM_PROBE70
    always @ (posedge clk)
    begin
      shift_probe70 <= probe70;
      mem_shift_probe70 <= shift_probe70;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 71) begin : FF_MEM_PROBE71
    always @ (posedge clk)
    begin
      shift_probe71 <= probe71;
      mem_shift_probe71 <= shift_probe71;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 72) begin : FF_MEM_PROBE72
    always @ (posedge clk)
    begin
      shift_probe72 <= probe72;
      mem_shift_probe72 <= shift_probe72;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 73) begin : FF_MEM_PROBE73
    always @ (posedge clk)
    begin
      shift_probe73 <= probe73;
      mem_shift_probe73 <= shift_probe73;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 74) begin : FF_MEM_PROBE74
    always @ (posedge clk)
    begin
      shift_probe74 <= probe74;
      mem_shift_probe74 <= shift_probe74;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 75) begin : FF_MEM_PROBE75
    always @ (posedge clk)
    begin
      shift_probe75 <= probe75;
      mem_shift_probe75 <= shift_probe75;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 76) begin : FF_MEM_PROBE76
    always @ (posedge clk)
    begin
      shift_probe76 <= probe76;
      mem_shift_probe76 <= shift_probe76;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 77) begin : FF_MEM_PROBE77
    always @ (posedge clk)
    begin
      shift_probe77 <= probe77;
      mem_shift_probe77 <= shift_probe77;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 78) begin : FF_MEM_PROBE78
    always @ (posedge clk)
    begin
      shift_probe78 <= probe78;
      mem_shift_probe78 <= shift_probe78;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 79) begin : FF_MEM_PROBE79
    always @ (posedge clk)
    begin
      shift_probe79 <= probe79;
      mem_shift_probe79 <= shift_probe79;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 80) begin : FF_MEM_PROBE80
    always @ (posedge clk)
    begin
      shift_probe80 <= probe80;
      mem_shift_probe80 <= shift_probe80;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 81) begin : FF_MEM_PROBE81
    always @ (posedge clk)
    begin
      shift_probe81 <= probe81;
      mem_shift_probe81 <= shift_probe81;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 82) begin : FF_MEM_PROBE82
    always @ (posedge clk)
    begin
      shift_probe82 <= probe82;
      mem_shift_probe82 <= shift_probe82;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 83) begin : FF_MEM_PROBE83
    always @ (posedge clk)
    begin
      shift_probe83 <= probe83;
      mem_shift_probe83 <= shift_probe83;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 84) begin : FF_MEM_PROBE84
    always @ (posedge clk)
    begin
      shift_probe84 <= probe84;
      mem_shift_probe84 <= shift_probe84;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 85) begin : FF_MEM_PROBE85
    always @ (posedge clk)
    begin
      shift_probe85 <= probe85;
      mem_shift_probe85 <= shift_probe85;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 86) begin : FF_MEM_PROBE86
    always @ (posedge clk)
    begin
      shift_probe86 <= probe86;
      mem_shift_probe86 <= shift_probe86;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 87) begin : FF_MEM_PROBE87
    always @ (posedge clk)
    begin
      shift_probe87 <= probe87;
      mem_shift_probe87 <= shift_probe87;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 88) begin : FF_MEM_PROBE88
    always @ (posedge clk)
    begin
      shift_probe88 <= probe88;
      mem_shift_probe88 <= shift_probe88;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 89) begin : FF_MEM_PROBE89
    always @ (posedge clk)
    begin
      shift_probe89 <= probe89;
      mem_shift_probe89 <= shift_probe89;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 90) begin : FF_MEM_PROBE90
    always @ (posedge clk)
    begin
      shift_probe90 <= probe90;
      mem_shift_probe90 <= shift_probe90;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 91) begin : FF_MEM_PROBE91
    always @ (posedge clk)
    begin
      shift_probe91 <= probe91;
      mem_shift_probe91 <= shift_probe91;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 92) begin : FF_MEM_PROBE92
    always @ (posedge clk)
    begin
      shift_probe92 <= probe92;
      mem_shift_probe92 <= shift_probe92;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 93) begin : FF_MEM_PROBE93
    always @ (posedge clk)
    begin
      shift_probe93 <= probe93;
      mem_shift_probe93 <= shift_probe93;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 94) begin : FF_MEM_PROBE94
    always @ (posedge clk)
    begin
      shift_probe94 <= probe94;
      mem_shift_probe94 <= shift_probe94;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 95) begin : FF_MEM_PROBE95
    always @ (posedge clk)
    begin
      shift_probe95 <= probe95;
      mem_shift_probe95 <= shift_probe95;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 96) begin : FF_MEM_PROBE96
    always @ (posedge clk)
    begin
      shift_probe96 <= probe96;
      mem_shift_probe96 <= shift_probe96;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 97) begin : FF_MEM_PROBE97
    always @ (posedge clk)
    begin
      shift_probe97 <= probe97;
      mem_shift_probe97 <= shift_probe97;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 98) begin : FF_MEM_PROBE98
    always @ (posedge clk)
    begin
      shift_probe98 <= probe98;
      mem_shift_probe98 <= shift_probe98;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 99) begin : FF_MEM_PROBE99
    always @ (posedge clk)
    begin
      shift_probe99 <= probe99;
      mem_shift_probe99 <= shift_probe99;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 100) begin : FF_MEM_PROBE100
    always @ (posedge clk)
    begin
      shift_probe100 <= probe100;
      mem_shift_probe100 <= shift_probe100;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 101) begin : FF_MEM_PROBE101
    always @ (posedge clk)
    begin
      shift_probe101 <= probe101;
      mem_shift_probe101 <= shift_probe101;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 102) begin : FF_MEM_PROBE102
    always @ (posedge clk)
    begin
      shift_probe102 <= probe102;
      mem_shift_probe102 <= shift_probe102;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 103) begin : FF_MEM_PROBE103
    always @ (posedge clk)
    begin
      shift_probe103 <= probe103;
      mem_shift_probe103 <= shift_probe103;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 104) begin : FF_MEM_PROBE104
    always @ (posedge clk)
    begin
      shift_probe104 <= probe104;
      mem_shift_probe104 <= shift_probe104;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 105) begin : FF_MEM_PROBE105
    always @ (posedge clk)
    begin
      shift_probe105 <= probe105;
      mem_shift_probe105 <= shift_probe105;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 106) begin : FF_MEM_PROBE106
    always @ (posedge clk)
    begin
      shift_probe106 <= probe106;
      mem_shift_probe106 <= shift_probe106;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 107) begin : FF_MEM_PROBE107
    always @ (posedge clk)
    begin
      shift_probe107 <= probe107;
      mem_shift_probe107 <= shift_probe107;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 108) begin : FF_MEM_PROBE108
    always @ (posedge clk)
    begin
      shift_probe108 <= probe108;
      mem_shift_probe108 <= shift_probe108;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 109) begin : FF_MEM_PROBE109
    always @ (posedge clk)
    begin
      shift_probe109 <= probe109;
      mem_shift_probe109 <= shift_probe109;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 110) begin : FF_MEM_PROBE110
    always @ (posedge clk)
    begin
      shift_probe110 <= probe110;
      mem_shift_probe110 <= shift_probe110;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 111) begin : FF_MEM_PROBE111
    always @ (posedge clk)
    begin
      shift_probe111 <= probe111;
      mem_shift_probe111 <= shift_probe111;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 112) begin : FF_MEM_PROBE112
    always @ (posedge clk)
    begin
      shift_probe112 <= probe112;
      mem_shift_probe112 <= shift_probe112;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 113) begin : FF_MEM_PROBE113
    always @ (posedge clk)
    begin
      shift_probe113 <= probe113;
      mem_shift_probe113 <= shift_probe113;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 114) begin : FF_MEM_PROBE114
    always @ (posedge clk)
    begin
      shift_probe114 <= probe114;
      mem_shift_probe114 <= shift_probe114;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 115) begin : FF_MEM_PROBE115
    always @ (posedge clk)
    begin
      shift_probe115 <= probe115;
      mem_shift_probe115 <= shift_probe115;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 116) begin : FF_MEM_PROBE116
    always @ (posedge clk)
    begin
      shift_probe116 <= probe116;
      mem_shift_probe116 <= shift_probe116;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 117) begin : FF_MEM_PROBE117
    always @ (posedge clk)
    begin
      shift_probe117 <= probe117;
      mem_shift_probe117 <= shift_probe117;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 118) begin : FF_MEM_PROBE118
    always @ (posedge clk)
    begin
      shift_probe118 <= probe118;
      mem_shift_probe118 <= shift_probe118;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 119) begin : FF_MEM_PROBE119
    always @ (posedge clk)
    begin
      shift_probe119 <= probe119;
      mem_shift_probe119 <= shift_probe119;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 120) begin : FF_MEM_PROBE120
    always @ (posedge clk)
    begin
      shift_probe120 <= probe120;
      mem_shift_probe120 <= shift_probe120;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 121) begin : FF_MEM_PROBE121
    always @ (posedge clk)
    begin
      shift_probe121 <= probe121;
      mem_shift_probe121 <= shift_probe121;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 122) begin : FF_MEM_PROBE122
    always @ (posedge clk)
    begin
      shift_probe122 <= probe122;
      mem_shift_probe122 <= shift_probe122;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 123) begin : FF_MEM_PROBE123
    always @ (posedge clk)
    begin
      shift_probe123 <= probe123;
      mem_shift_probe123 <= shift_probe123;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 124) begin : FF_MEM_PROBE124
    always @ (posedge clk)
    begin
      shift_probe124 <= probe124;
      mem_shift_probe124 <= shift_probe124;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 125) begin : FF_MEM_PROBE125
    always @ (posedge clk)
    begin
      shift_probe125 <= probe125;
      mem_shift_probe125 <= shift_probe125;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 126) begin : FF_MEM_PROBE126
    always @ (posedge clk)
    begin
      shift_probe126 <= probe126;
      mem_shift_probe126 <= shift_probe126;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 127) begin : FF_MEM_PROBE127
    always @ (posedge clk)
    begin
      shift_probe127 <= probe127;
      mem_shift_probe127 <= shift_probe127;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 128) begin : FF_MEM_PROBE128
    always @ (posedge clk)
    begin
      shift_probe128 <= probe128;
      mem_shift_probe128 <= shift_probe128;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 129) begin : FF_MEM_PROBE129
    always @ (posedge clk)
    begin
      shift_probe129 <= probe129;
      mem_shift_probe129 <= shift_probe129;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 130) begin : FF_MEM_PROBE130
    always @ (posedge clk)
    begin
      shift_probe130 <= probe130;
      mem_shift_probe130 <= shift_probe130;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 131) begin : FF_MEM_PROBE131
    always @ (posedge clk)
    begin
      shift_probe131 <= probe131;
      mem_shift_probe131 <= shift_probe131;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 132) begin : FF_MEM_PROBE132
    always @ (posedge clk)
    begin
      shift_probe132 <= probe132;
      mem_shift_probe132 <= shift_probe132;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 133) begin : FF_MEM_PROBE133
    always @ (posedge clk)
    begin
      shift_probe133 <= probe133;
      mem_shift_probe133 <= shift_probe133;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 134) begin : FF_MEM_PROBE134
    always @ (posedge clk)
    begin
      shift_probe134 <= probe134;
      mem_shift_probe134 <= shift_probe134;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 135) begin : FF_MEM_PROBE135
    always @ (posedge clk)
    begin
      shift_probe135 <= probe135;
      mem_shift_probe135 <= shift_probe135;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 136) begin : FF_MEM_PROBE136
    always @ (posedge clk)
    begin
      shift_probe136 <= probe136;
      mem_shift_probe136 <= shift_probe136;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 137) begin : FF_MEM_PROBE137
    always @ (posedge clk)
    begin
      shift_probe137 <= probe137;
      mem_shift_probe137 <= shift_probe137;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 138) begin : FF_MEM_PROBE138
    always @ (posedge clk)
    begin
      shift_probe138 <= probe138;
      mem_shift_probe138 <= shift_probe138;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 139) begin : FF_MEM_PROBE139
    always @ (posedge clk)
    begin
      shift_probe139 <= probe139;
      mem_shift_probe139 <= shift_probe139;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 140) begin : FF_MEM_PROBE140
    always @ (posedge clk)
    begin
      shift_probe140 <= probe140;
      mem_shift_probe140 <= shift_probe140;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 141) begin : FF_MEM_PROBE141
    always @ (posedge clk)
    begin
      shift_probe141 <= probe141;
      mem_shift_probe141 <= shift_probe141;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 142) begin : FF_MEM_PROBE142
    always @ (posedge clk)
    begin
      shift_probe142 <= probe142;
      mem_shift_probe142 <= shift_probe142;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 143) begin : FF_MEM_PROBE143
    always @ (posedge clk)
    begin
      shift_probe143 <= probe143;
      mem_shift_probe143 <= shift_probe143;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 144) begin : FF_MEM_PROBE144
    always @ (posedge clk)
    begin
      shift_probe144 <= probe144;
      mem_shift_probe144 <= shift_probe144;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 145) begin : FF_MEM_PROBE145
    always @ (posedge clk)
    begin
      shift_probe145 <= probe145;
      mem_shift_probe145 <= shift_probe145;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 146) begin : FF_MEM_PROBE146
    always @ (posedge clk)
    begin
      shift_probe146 <= probe146;
      mem_shift_probe146 <= shift_probe146;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 147) begin : FF_MEM_PROBE147
    always @ (posedge clk)
    begin
      shift_probe147 <= probe147;
      mem_shift_probe147 <= shift_probe147;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 148) begin : FF_MEM_PROBE148
    always @ (posedge clk)
    begin
      shift_probe148 <= probe148;
      mem_shift_probe148 <= shift_probe148;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 149) begin : FF_MEM_PROBE149
    always @ (posedge clk)
    begin
      shift_probe149 <= probe149;
      mem_shift_probe149 <= shift_probe149;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 150) begin : FF_MEM_PROBE150
    always @ (posedge clk)
    begin
      shift_probe150 <= probe150;
      mem_shift_probe150 <= shift_probe150;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 151) begin : FF_MEM_PROBE151
    always @ (posedge clk)
    begin
      shift_probe151 <= probe151;
      mem_shift_probe151 <= shift_probe151;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 152) begin : FF_MEM_PROBE152
    always @ (posedge clk)
    begin
      shift_probe152 <= probe152;
      mem_shift_probe152 <= shift_probe152;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 153) begin : FF_MEM_PROBE153
    always @ (posedge clk)
    begin
      shift_probe153 <= probe153;
      mem_shift_probe153 <= shift_probe153;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 154) begin : FF_MEM_PROBE154
    always @ (posedge clk)
    begin
      shift_probe154 <= probe154;
      mem_shift_probe154 <= shift_probe154;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 155) begin : FF_MEM_PROBE155
    always @ (posedge clk)
    begin
      shift_probe155 <= probe155;
      mem_shift_probe155 <= shift_probe155;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 156) begin : FF_MEM_PROBE156
    always @ (posedge clk)
    begin
      shift_probe156 <= probe156;
      mem_shift_probe156 <= shift_probe156;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 157) begin : FF_MEM_PROBE157
    always @ (posedge clk)
    begin
      shift_probe157 <= probe157;
      mem_shift_probe157 <= shift_probe157;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 158) begin : FF_MEM_PROBE158
    always @ (posedge clk)
    begin
      shift_probe158 <= probe158;
      mem_shift_probe158 <= shift_probe158;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 159) begin : FF_MEM_PROBE159
    always @ (posedge clk)
    begin
      shift_probe159 <= probe159;
      mem_shift_probe159 <= shift_probe159;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 160) begin : FF_MEM_PROBE160
    always @ (posedge clk)
    begin
      shift_probe160 <= probe160;
      mem_shift_probe160 <= shift_probe160;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 161) begin : FF_MEM_PROBE161
    always @ (posedge clk)
    begin
      shift_probe161 <= probe161;
      mem_shift_probe161 <= shift_probe161;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 162) begin : FF_MEM_PROBE162
    always @ (posedge clk)
    begin
      shift_probe162 <= probe162;
      mem_shift_probe162 <= shift_probe162;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 163) begin : FF_MEM_PROBE163
    always @ (posedge clk)
    begin
      shift_probe163 <= probe163;
      mem_shift_probe163 <= shift_probe163;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 164) begin : FF_MEM_PROBE164
    always @ (posedge clk)
    begin
      shift_probe164 <= probe164;
      mem_shift_probe164 <= shift_probe164;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 165) begin : FF_MEM_PROBE165
    always @ (posedge clk)
    begin
      shift_probe165 <= probe165;
      mem_shift_probe165 <= shift_probe165;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 166) begin : FF_MEM_PROBE166
    always @ (posedge clk)
    begin
      shift_probe166 <= probe166;
      mem_shift_probe166 <= shift_probe166;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 167) begin : FF_MEM_PROBE167
    always @ (posedge clk)
    begin
      shift_probe167 <= probe167;
      mem_shift_probe167 <= shift_probe167;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 168) begin : FF_MEM_PROBE168
    always @ (posedge clk)
    begin
      shift_probe168 <= probe168;
      mem_shift_probe168 <= shift_probe168;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 169) begin : FF_MEM_PROBE169
    always @ (posedge clk)
    begin
      shift_probe169 <= probe169;
      mem_shift_probe169 <= shift_probe169;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 170) begin : FF_MEM_PROBE170
    always @ (posedge clk)
    begin
      shift_probe170 <= probe170;
      mem_shift_probe170 <= shift_probe170;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 171) begin : FF_MEM_PROBE171
    always @ (posedge clk)
    begin
      shift_probe171 <= probe171;
      mem_shift_probe171 <= shift_probe171;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 172) begin : FF_MEM_PROBE172
    always @ (posedge clk)
    begin
      shift_probe172 <= probe172;
      mem_shift_probe172 <= shift_probe172;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 173) begin : FF_MEM_PROBE173
    always @ (posedge clk)
    begin
      shift_probe173 <= probe173;
      mem_shift_probe173 <= shift_probe173;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 174) begin : FF_MEM_PROBE174
    always @ (posedge clk)
    begin
      shift_probe174 <= probe174;
      mem_shift_probe174 <= shift_probe174;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 175) begin : FF_MEM_PROBE175
    always @ (posedge clk)
    begin
      shift_probe175 <= probe175;
      mem_shift_probe175 <= shift_probe175;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 176) begin : FF_MEM_PROBE176
    always @ (posedge clk)
    begin
      shift_probe176 <= probe176;
      mem_shift_probe176 <= shift_probe176;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 177) begin : FF_MEM_PROBE177
    always @ (posedge clk)
    begin
      shift_probe177 <= probe177;
      mem_shift_probe177 <= shift_probe177;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 178) begin : FF_MEM_PROBE178
    always @ (posedge clk)
    begin
      shift_probe178 <= probe178;
      mem_shift_probe178 <= shift_probe178;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 179) begin : FF_MEM_PROBE179
    always @ (posedge clk)
    begin
      shift_probe179 <= probe179;
      mem_shift_probe179 <= shift_probe179;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 180) begin : FF_MEM_PROBE180
    always @ (posedge clk)
    begin
      shift_probe180 <= probe180;
      mem_shift_probe180 <= shift_probe180;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 181) begin : FF_MEM_PROBE181
    always @ (posedge clk)
    begin
      shift_probe181 <= probe181;
      mem_shift_probe181 <= shift_probe181;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 182) begin : FF_MEM_PROBE182
    always @ (posedge clk)
    begin
      shift_probe182 <= probe182;
      mem_shift_probe182 <= shift_probe182;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 183) begin : FF_MEM_PROBE183
    always @ (posedge clk)
    begin
      shift_probe183 <= probe183;
      mem_shift_probe183 <= shift_probe183;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 184) begin : FF_MEM_PROBE184
    always @ (posedge clk)
    begin
      shift_probe184 <= probe184;
      mem_shift_probe184 <= shift_probe184;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 185) begin : FF_MEM_PROBE185
    always @ (posedge clk)
    begin
      shift_probe185 <= probe185;
      mem_shift_probe185 <= shift_probe185;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 186) begin : FF_MEM_PROBE186
    always @ (posedge clk)
    begin
      shift_probe186 <= probe186;
      mem_shift_probe186 <= shift_probe186;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 187) begin : FF_MEM_PROBE187
    always @ (posedge clk)
    begin
      shift_probe187 <= probe187;
      mem_shift_probe187 <= shift_probe187;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 188) begin : FF_MEM_PROBE188
    always @ (posedge clk)
    begin
      shift_probe188 <= probe188;
      mem_shift_probe188 <= shift_probe188;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 189) begin : FF_MEM_PROBE189
    always @ (posedge clk)
    begin
      shift_probe189 <= probe189;
      mem_shift_probe189 <= shift_probe189;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 190) begin : FF_MEM_PROBE190
    always @ (posedge clk)
    begin
      shift_probe190 <= probe190;
      mem_shift_probe190 <= shift_probe190;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 191) begin : FF_MEM_PROBE191
    always @ (posedge clk)
    begin
      shift_probe191 <= probe191;
      mem_shift_probe191 <= shift_probe191;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 192) begin : FF_MEM_PROBE192
    always @ (posedge clk)
    begin
      shift_probe192 <= probe192;
      mem_shift_probe192 <= shift_probe192;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 193) begin : FF_MEM_PROBE193
    always @ (posedge clk)
    begin
      shift_probe193 <= probe193;
      mem_shift_probe193 <= shift_probe193;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 194) begin : FF_MEM_PROBE194
    always @ (posedge clk)
    begin
      shift_probe194 <= probe194;
      mem_shift_probe194 <= shift_probe194;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 195) begin : FF_MEM_PROBE195
    always @ (posedge clk)
    begin
      shift_probe195 <= probe195;
      mem_shift_probe195 <= shift_probe195;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 196) begin : FF_MEM_PROBE196
    always @ (posedge clk)
    begin
      shift_probe196 <= probe196;
      mem_shift_probe196 <= shift_probe196;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 197) begin : FF_MEM_PROBE197
    always @ (posedge clk)
    begin
      shift_probe197 <= probe197;
      mem_shift_probe197 <= shift_probe197;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 198) begin : FF_MEM_PROBE198
    always @ (posedge clk)
    begin
      shift_probe198 <= probe198;
      mem_shift_probe198 <= shift_probe198;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 199) begin : FF_MEM_PROBE199
    always @ (posedge clk)
    begin
      shift_probe199 <= probe199;
      mem_shift_probe199 <= shift_probe199;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 200) begin : FF_MEM_PROBE200
    always @ (posedge clk)
    begin
      shift_probe200 <= probe200;
      mem_shift_probe200 <= shift_probe200;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 201) begin : FF_MEM_PROBE201
    always @ (posedge clk)
    begin
      shift_probe201 <= probe201;
      mem_shift_probe201 <= shift_probe201;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 202) begin : FF_MEM_PROBE202
    always @ (posedge clk)
    begin
      shift_probe202 <= probe202;
      mem_shift_probe202 <= shift_probe202;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 203) begin : FF_MEM_PROBE203
    always @ (posedge clk)
    begin
      shift_probe203 <= probe203;
      mem_shift_probe203 <= shift_probe203;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 204) begin : FF_MEM_PROBE204
    always @ (posedge clk)
    begin
      shift_probe204 <= probe204;
      mem_shift_probe204 <= shift_probe204;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 205) begin : FF_MEM_PROBE205
    always @ (posedge clk)
    begin
      shift_probe205 <= probe205;
      mem_shift_probe205 <= shift_probe205;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 206) begin : FF_MEM_PROBE206
    always @ (posedge clk)
    begin
      shift_probe206 <= probe206;
      mem_shift_probe206 <= shift_probe206;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 207) begin : FF_MEM_PROBE207
    always @ (posedge clk)
    begin
      shift_probe207 <= probe207;
      mem_shift_probe207 <= shift_probe207;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 208) begin : FF_MEM_PROBE208
    always @ (posedge clk)
    begin
      shift_probe208 <= probe208;
      mem_shift_probe208 <= shift_probe208;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 209) begin : FF_MEM_PROBE209
    always @ (posedge clk)
    begin
      shift_probe209 <= probe209;
      mem_shift_probe209 <= shift_probe209;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 210) begin : FF_MEM_PROBE210
    always @ (posedge clk)
    begin
      shift_probe210 <= probe210;
      mem_shift_probe210 <= shift_probe210;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 211) begin : FF_MEM_PROBE211
    always @ (posedge clk)
    begin
      shift_probe211 <= probe211;
      mem_shift_probe211 <= shift_probe211;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 212) begin : FF_MEM_PROBE212
    always @ (posedge clk)
    begin
      shift_probe212 <= probe212;
      mem_shift_probe212 <= shift_probe212;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 213) begin : FF_MEM_PROBE213
    always @ (posedge clk)
    begin
      shift_probe213 <= probe213;
      mem_shift_probe213 <= shift_probe213;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 214) begin : FF_MEM_PROBE214
    always @ (posedge clk)
    begin
      shift_probe214 <= probe214;
      mem_shift_probe214 <= shift_probe214;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 215) begin : FF_MEM_PROBE215
    always @ (posedge clk)
    begin
      shift_probe215 <= probe215;
      mem_shift_probe215 <= shift_probe215;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 216) begin : FF_MEM_PROBE216
    always @ (posedge clk)
    begin
      shift_probe216 <= probe216;
      mem_shift_probe216 <= shift_probe216;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 217) begin : FF_MEM_PROBE217
    always @ (posedge clk)
    begin
      shift_probe217 <= probe217;
      mem_shift_probe217 <= shift_probe217;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 218) begin : FF_MEM_PROBE218
    always @ (posedge clk)
    begin
      shift_probe218 <= probe218;
      mem_shift_probe218 <= shift_probe218;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 219) begin : FF_MEM_PROBE219
    always @ (posedge clk)
    begin
      shift_probe219 <= probe219;
      mem_shift_probe219 <= shift_probe219;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 220) begin : FF_MEM_PROBE220
    always @ (posedge clk)
    begin
      shift_probe220 <= probe220;
      mem_shift_probe220 <= shift_probe220;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 221) begin : FF_MEM_PROBE221
    always @ (posedge clk)
    begin
      shift_probe221 <= probe221;
      mem_shift_probe221 <= shift_probe221;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 222) begin : FF_MEM_PROBE222
    always @ (posedge clk)
    begin
      shift_probe222 <= probe222;
      mem_shift_probe222 <= shift_probe222;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 223) begin : FF_MEM_PROBE223
    always @ (posedge clk)
    begin
      shift_probe223 <= probe223;
      mem_shift_probe223 <= shift_probe223;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 224) begin : FF_MEM_PROBE224
    always @ (posedge clk)
    begin
      shift_probe224 <= probe224;
      mem_shift_probe224 <= shift_probe224;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 225) begin : FF_MEM_PROBE225
    always @ (posedge clk)
    begin
      shift_probe225 <= probe225;
      mem_shift_probe225 <= shift_probe225;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 226) begin : FF_MEM_PROBE226
    always @ (posedge clk)
    begin
      shift_probe226 <= probe226;
      mem_shift_probe226 <= shift_probe226;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 227) begin : FF_MEM_PROBE227
    always @ (posedge clk)
    begin
      shift_probe227 <= probe227;
      mem_shift_probe227 <= shift_probe227;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 228) begin : FF_MEM_PROBE228
    always @ (posedge clk)
    begin
      shift_probe228 <= probe228;
      mem_shift_probe228 <= shift_probe228;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 229) begin : FF_MEM_PROBE229
    always @ (posedge clk)
    begin
      shift_probe229 <= probe229;
      mem_shift_probe229 <= shift_probe229;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 230) begin : FF_MEM_PROBE230
    always @ (posedge clk)
    begin
      shift_probe230 <= probe230;
      mem_shift_probe230 <= shift_probe230;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 231) begin : FF_MEM_PROBE231
    always @ (posedge clk)
    begin
      shift_probe231 <= probe231;
      mem_shift_probe231 <= shift_probe231;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 232) begin : FF_MEM_PROBE232
    always @ (posedge clk)
    begin
      shift_probe232 <= probe232;
      mem_shift_probe232 <= shift_probe232;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 233) begin : FF_MEM_PROBE233
    always @ (posedge clk)
    begin
      shift_probe233 <= probe233;
      mem_shift_probe233 <= shift_probe233;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 234) begin : FF_MEM_PROBE234
    always @ (posedge clk)
    begin
      shift_probe234 <= probe234;
      mem_shift_probe234 <= shift_probe234;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 235) begin : FF_MEM_PROBE235
    always @ (posedge clk)
    begin
      shift_probe235 <= probe235;
      mem_shift_probe235 <= shift_probe235;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 236) begin : FF_MEM_PROBE236
    always @ (posedge clk)
    begin
      shift_probe236 <= probe236;
      mem_shift_probe236 <= shift_probe236;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 237) begin : FF_MEM_PROBE237
    always @ (posedge clk)
    begin
      shift_probe237 <= probe237;
      mem_shift_probe237 <= shift_probe237;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 238) begin : FF_MEM_PROBE238
    always @ (posedge clk)
    begin
      shift_probe238 <= probe238;
      mem_shift_probe238 <= shift_probe238;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 239) begin : FF_MEM_PROBE239
    always @ (posedge clk)
    begin
      shift_probe239 <= probe239;
      mem_shift_probe239 <= shift_probe239;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 240) begin : FF_MEM_PROBE240
    always @ (posedge clk)
    begin
      shift_probe240 <= probe240;
      mem_shift_probe240 <= shift_probe240;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 241) begin : FF_MEM_PROBE241
    always @ (posedge clk)
    begin
      shift_probe241 <= probe241;
      mem_shift_probe241 <= shift_probe241;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 242) begin : FF_MEM_PROBE242
    always @ (posedge clk)
    begin
      shift_probe242 <= probe242;
      mem_shift_probe242 <= shift_probe242;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 243) begin : FF_MEM_PROBE243
    always @ (posedge clk)
    begin
      shift_probe243 <= probe243;
      mem_shift_probe243 <= shift_probe243;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 244) begin : FF_MEM_PROBE244
    always @ (posedge clk)
    begin
      shift_probe244 <= probe244;
      mem_shift_probe244 <= shift_probe244;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 245) begin : FF_MEM_PROBE245
    always @ (posedge clk)
    begin
      shift_probe245 <= probe245;
      mem_shift_probe245 <= shift_probe245;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 246) begin : FF_MEM_PROBE246
    always @ (posedge clk)
    begin
      shift_probe246 <= probe246;
      mem_shift_probe246 <= shift_probe246;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 247) begin : FF_MEM_PROBE247
    always @ (posedge clk)
    begin
      shift_probe247 <= probe247;
      mem_shift_probe247 <= shift_probe247;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 248) begin : FF_MEM_PROBE248
    always @ (posedge clk)
    begin
      shift_probe248 <= probe248;
      mem_shift_probe248 <= shift_probe248;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 249) begin : FF_MEM_PROBE249
    always @ (posedge clk)
    begin
      shift_probe249 <= probe249;
      mem_shift_probe249 <= shift_probe249;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 250) begin : FF_MEM_PROBE250
    always @ (posedge clk)
    begin
      shift_probe250 <= probe250;
      mem_shift_probe250 <= shift_probe250;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 251) begin : FF_MEM_PROBE251
    always @ (posedge clk)
    begin
      shift_probe251 <= probe251;
      mem_shift_probe251 <= shift_probe251;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 252) begin : FF_MEM_PROBE252
    always @ (posedge clk)
    begin
      shift_probe252 <= probe252;
      mem_shift_probe252 <= shift_probe252;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 253) begin : FF_MEM_PROBE253
    always @ (posedge clk)
    begin
      shift_probe253 <= probe253;
      mem_shift_probe253 <= shift_probe253;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 254) begin : FF_MEM_PROBE254
    always @ (posedge clk)
    begin
      shift_probe254 <= probe254;
      mem_shift_probe254 <= shift_probe254;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 255) begin : FF_MEM_PROBE255
    always @ (posedge clk)
    begin
      shift_probe255 <= probe255;
      mem_shift_probe255 <= shift_probe255;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 256) begin : FF_MEM_PROBE256
    always @ (posedge clk)
    begin
      shift_probe256 <= probe256;
      mem_shift_probe256 <= shift_probe256;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 257) begin : FF_MEM_PROBE257
    always @ (posedge clk)
    begin
      shift_probe257 <= probe257;
      mem_shift_probe257 <= shift_probe257;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 258) begin : FF_MEM_PROBE258
    always @ (posedge clk)
    begin
      shift_probe258 <= probe258;
      mem_shift_probe258 <= shift_probe258;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 259) begin : FF_MEM_PROBE259
    always @ (posedge clk)
    begin
      shift_probe259 <= probe259;
      mem_shift_probe259 <= shift_probe259;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 260) begin : FF_MEM_PROBE260
    always @ (posedge clk)
    begin
      shift_probe260 <= probe260;
      mem_shift_probe260 <= shift_probe260;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 261) begin : FF_MEM_PROBE261
    always @ (posedge clk)
    begin
      shift_probe261 <= probe261;
      mem_shift_probe261 <= shift_probe261;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 262) begin : FF_MEM_PROBE262
    always @ (posedge clk)
    begin
      shift_probe262 <= probe262;
      mem_shift_probe262 <= shift_probe262;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 263) begin : FF_MEM_PROBE263
    always @ (posedge clk)
    begin
      shift_probe263 <= probe263;
      mem_shift_probe263 <= shift_probe263;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 264) begin : FF_MEM_PROBE264
    always @ (posedge clk)
    begin
      shift_probe264 <= probe264;
      mem_shift_probe264 <= shift_probe264;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 265) begin : FF_MEM_PROBE265
    always @ (posedge clk)
    begin
      shift_probe265 <= probe265;
      mem_shift_probe265 <= shift_probe265;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 266) begin : FF_MEM_PROBE266
    always @ (posedge clk)
    begin
      shift_probe266 <= probe266;
      mem_shift_probe266 <= shift_probe266;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 267) begin : FF_MEM_PROBE267
    always @ (posedge clk)
    begin
      shift_probe267 <= probe267;
      mem_shift_probe267 <= shift_probe267;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 268) begin : FF_MEM_PROBE268
    always @ (posedge clk)
    begin
      shift_probe268 <= probe268;
      mem_shift_probe268 <= shift_probe268;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 269) begin : FF_MEM_PROBE269
    always @ (posedge clk)
    begin
      shift_probe269 <= probe269;
      mem_shift_probe269 <= shift_probe269;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 270) begin : FF_MEM_PROBE270
    always @ (posedge clk)
    begin
      shift_probe270 <= probe270;
      mem_shift_probe270 <= shift_probe270;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 271) begin : FF_MEM_PROBE271
    always @ (posedge clk)
    begin
      shift_probe271 <= probe271;
      mem_shift_probe271 <= shift_probe271;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 272) begin : FF_MEM_PROBE272
    always @ (posedge clk)
    begin
      shift_probe272 <= probe272;
      mem_shift_probe272 <= shift_probe272;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 273) begin : FF_MEM_PROBE273
    always @ (posedge clk)
    begin
      shift_probe273 <= probe273;
      mem_shift_probe273 <= shift_probe273;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 274) begin : FF_MEM_PROBE274
    always @ (posedge clk)
    begin
      shift_probe274 <= probe274;
      mem_shift_probe274 <= shift_probe274;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 275) begin : FF_MEM_PROBE275
    always @ (posedge clk)
    begin
      shift_probe275 <= probe275;
      mem_shift_probe275 <= shift_probe275;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 276) begin : FF_MEM_PROBE276
    always @ (posedge clk)
    begin
      shift_probe276 <= probe276;
      mem_shift_probe276 <= shift_probe276;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 277) begin : FF_MEM_PROBE277
    always @ (posedge clk)
    begin
      shift_probe277 <= probe277;
      mem_shift_probe277 <= shift_probe277;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 278) begin : FF_MEM_PROBE278
    always @ (posedge clk)
    begin
      shift_probe278 <= probe278;
      mem_shift_probe278 <= shift_probe278;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 279) begin : FF_MEM_PROBE279
    always @ (posedge clk)
    begin
      shift_probe279 <= probe279;
      mem_shift_probe279 <= shift_probe279;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 280) begin : FF_MEM_PROBE280
    always @ (posedge clk)
    begin
      shift_probe280 <= probe280;
      mem_shift_probe280 <= shift_probe280;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 281) begin : FF_MEM_PROBE281
    always @ (posedge clk)
    begin
      shift_probe281 <= probe281;
      mem_shift_probe281 <= shift_probe281;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 282) begin : FF_MEM_PROBE282
    always @ (posedge clk)
    begin
      shift_probe282 <= probe282;
      mem_shift_probe282 <= shift_probe282;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 283) begin : FF_MEM_PROBE283
    always @ (posedge clk)
    begin
      shift_probe283 <= probe283;
      mem_shift_probe283 <= shift_probe283;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 284) begin : FF_MEM_PROBE284
    always @ (posedge clk)
    begin
      shift_probe284 <= probe284;
      mem_shift_probe284 <= shift_probe284;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 285) begin : FF_MEM_PROBE285
    always @ (posedge clk)
    begin
      shift_probe285 <= probe285;
      mem_shift_probe285 <= shift_probe285;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 286) begin : FF_MEM_PROBE286
    always @ (posedge clk)
    begin
      shift_probe286 <= probe286;
      mem_shift_probe286 <= shift_probe286;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 287) begin : FF_MEM_PROBE287
    always @ (posedge clk)
    begin
      shift_probe287 <= probe287;
      mem_shift_probe287 <= shift_probe287;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 288) begin : FF_MEM_PROBE288
    always @ (posedge clk)
    begin
      shift_probe288 <= probe288;
      mem_shift_probe288 <= shift_probe288;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 289) begin : FF_MEM_PROBE289
    always @ (posedge clk)
    begin
      shift_probe289 <= probe289;
      mem_shift_probe289 <= shift_probe289;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 290) begin : FF_MEM_PROBE290
    always @ (posedge clk)
    begin
      shift_probe290 <= probe290;
      mem_shift_probe290 <= shift_probe290;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 291) begin : FF_MEM_PROBE291
    always @ (posedge clk)
    begin
      shift_probe291 <= probe291;
      mem_shift_probe291 <= shift_probe291;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 292) begin : FF_MEM_PROBE292
    always @ (posedge clk)
    begin
      shift_probe292 <= probe292;
      mem_shift_probe292 <= shift_probe292;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 293) begin : FF_MEM_PROBE293
    always @ (posedge clk)
    begin
      shift_probe293 <= probe293;
      mem_shift_probe293 <= shift_probe293;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 294) begin : FF_MEM_PROBE294
    always @ (posedge clk)
    begin
      shift_probe294 <= probe294;
      mem_shift_probe294 <= shift_probe294;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 295) begin : FF_MEM_PROBE295
    always @ (posedge clk)
    begin
      shift_probe295 <= probe295;
      mem_shift_probe295 <= shift_probe295;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 296) begin : FF_MEM_PROBE296
    always @ (posedge clk)
    begin
      shift_probe296 <= probe296;
      mem_shift_probe296 <= shift_probe296;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 297) begin : FF_MEM_PROBE297
    always @ (posedge clk)
    begin
      shift_probe297 <= probe297;
      mem_shift_probe297 <= shift_probe297;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 298) begin : FF_MEM_PROBE298
    always @ (posedge clk)
    begin
      shift_probe298 <= probe298;
      mem_shift_probe298 <= shift_probe298;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 299) begin : FF_MEM_PROBE299
    always @ (posedge clk)
    begin
      shift_probe299 <= probe299;
      mem_shift_probe299 <= shift_probe299;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 300) begin : FF_MEM_PROBE300
    always @ (posedge clk)
    begin
      shift_probe300 <= probe300;
      mem_shift_probe300 <= shift_probe300;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 301) begin : FF_MEM_PROBE301
    always @ (posedge clk)
    begin
      shift_probe301 <= probe301;
      mem_shift_probe301 <= shift_probe301;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 302) begin : FF_MEM_PROBE302
    always @ (posedge clk)
    begin
      shift_probe302 <= probe302;
      mem_shift_probe302 <= shift_probe302;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 303) begin : FF_MEM_PROBE303
    always @ (posedge clk)
    begin
      shift_probe303 <= probe303;
      mem_shift_probe303 <= shift_probe303;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 304) begin : FF_MEM_PROBE304
    always @ (posedge clk)
    begin
      shift_probe304 <= probe304;
      mem_shift_probe304 <= shift_probe304;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 305) begin : FF_MEM_PROBE305
    always @ (posedge clk)
    begin
      shift_probe305 <= probe305;
      mem_shift_probe305 <= shift_probe305;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 306) begin : FF_MEM_PROBE306
    always @ (posedge clk)
    begin
      shift_probe306 <= probe306;
      mem_shift_probe306 <= shift_probe306;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 307) begin : FF_MEM_PROBE307
    always @ (posedge clk)
    begin
      shift_probe307 <= probe307;
      mem_shift_probe307 <= shift_probe307;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 308) begin : FF_MEM_PROBE308
    always @ (posedge clk)
    begin
      shift_probe308 <= probe308;
      mem_shift_probe308 <= shift_probe308;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 309) begin : FF_MEM_PROBE309
    always @ (posedge clk)
    begin
      shift_probe309 <= probe309;
      mem_shift_probe309 <= shift_probe309;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 310) begin : FF_MEM_PROBE310
    always @ (posedge clk)
    begin
      shift_probe310 <= probe310;
      mem_shift_probe310 <= shift_probe310;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 311) begin : FF_MEM_PROBE311
    always @ (posedge clk)
    begin
      shift_probe311 <= probe311;
      mem_shift_probe311 <= shift_probe311;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 312) begin : FF_MEM_PROBE312
    always @ (posedge clk)
    begin
      shift_probe312 <= probe312;
      mem_shift_probe312 <= shift_probe312;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 313) begin : FF_MEM_PROBE313
    always @ (posedge clk)
    begin
      shift_probe313 <= probe313;
      mem_shift_probe313 <= shift_probe313;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 314) begin : FF_MEM_PROBE314
    always @ (posedge clk)
    begin
      shift_probe314 <= probe314;
      mem_shift_probe314 <= shift_probe314;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 315) begin : FF_MEM_PROBE315
    always @ (posedge clk)
    begin
      shift_probe315 <= probe315;
      mem_shift_probe315 <= shift_probe315;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 316) begin : FF_MEM_PROBE316
    always @ (posedge clk)
    begin
      shift_probe316 <= probe316;
      mem_shift_probe316 <= shift_probe316;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 317) begin : FF_MEM_PROBE317
    always @ (posedge clk)
    begin
      shift_probe317 <= probe317;
      mem_shift_probe317 <= shift_probe317;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 318) begin : FF_MEM_PROBE318
    always @ (posedge clk)
    begin
      shift_probe318 <= probe318;
      mem_shift_probe318 <= shift_probe318;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 319) begin : FF_MEM_PROBE319
    always @ (posedge clk)
    begin
      shift_probe319 <= probe319;
      mem_shift_probe319 <= shift_probe319;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 320) begin : FF_MEM_PROBE320
    always @ (posedge clk)
    begin
      shift_probe320 <= probe320;
      mem_shift_probe320 <= shift_probe320;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 321) begin : FF_MEM_PROBE321
    always @ (posedge clk)
    begin
      shift_probe321 <= probe321;
      mem_shift_probe321 <= shift_probe321;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 322) begin : FF_MEM_PROBE322
    always @ (posedge clk)
    begin
      shift_probe322 <= probe322;
      mem_shift_probe322 <= shift_probe322;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 323) begin : FF_MEM_PROBE323
    always @ (posedge clk)
    begin
      shift_probe323 <= probe323;
      mem_shift_probe323 <= shift_probe323;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 324) begin : FF_MEM_PROBE324
    always @ (posedge clk)
    begin
      shift_probe324 <= probe324;
      mem_shift_probe324 <= shift_probe324;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 325) begin : FF_MEM_PROBE325
    always @ (posedge clk)
    begin
      shift_probe325 <= probe325;
      mem_shift_probe325 <= shift_probe325;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 326) begin : FF_MEM_PROBE326
    always @ (posedge clk)
    begin
      shift_probe326 <= probe326;
      mem_shift_probe326 <= shift_probe326;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 327) begin : FF_MEM_PROBE327
    always @ (posedge clk)
    begin
      shift_probe327 <= probe327;
      mem_shift_probe327 <= shift_probe327;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 328) begin : FF_MEM_PROBE328
    always @ (posedge clk)
    begin
      shift_probe328 <= probe328;
      mem_shift_probe328 <= shift_probe328;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 329) begin : FF_MEM_PROBE329
    always @ (posedge clk)
    begin
      shift_probe329 <= probe329;
      mem_shift_probe329 <= shift_probe329;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 330) begin : FF_MEM_PROBE330
    always @ (posedge clk)
    begin
      shift_probe330 <= probe330;
      mem_shift_probe330 <= shift_probe330;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 331) begin : FF_MEM_PROBE331
    always @ (posedge clk)
    begin
      shift_probe331 <= probe331;
      mem_shift_probe331 <= shift_probe331;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 332) begin : FF_MEM_PROBE332
    always @ (posedge clk)
    begin
      shift_probe332 <= probe332;
      mem_shift_probe332 <= shift_probe332;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 333) begin : FF_MEM_PROBE333
    always @ (posedge clk)
    begin
      shift_probe333 <= probe333;
      mem_shift_probe333 <= shift_probe333;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 334) begin : FF_MEM_PROBE334
    always @ (posedge clk)
    begin
      shift_probe334 <= probe334;
      mem_shift_probe334 <= shift_probe334;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 335) begin : FF_MEM_PROBE335
    always @ (posedge clk)
    begin
      shift_probe335 <= probe335;
      mem_shift_probe335 <= shift_probe335;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 336) begin : FF_MEM_PROBE336
    always @ (posedge clk)
    begin
      shift_probe336 <= probe336;
      mem_shift_probe336 <= shift_probe336;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 337) begin : FF_MEM_PROBE337
    always @ (posedge clk)
    begin
      shift_probe337 <= probe337;
      mem_shift_probe337 <= shift_probe337;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 338) begin : FF_MEM_PROBE338
    always @ (posedge clk)
    begin
      shift_probe338 <= probe338;
      mem_shift_probe338 <= shift_probe338;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 339) begin : FF_MEM_PROBE339
    always @ (posedge clk)
    begin
      shift_probe339 <= probe339;
      mem_shift_probe339 <= shift_probe339;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 340) begin : FF_MEM_PROBE340
    always @ (posedge clk)
    begin
      shift_probe340 <= probe340;
      mem_shift_probe340 <= shift_probe340;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 341) begin : FF_MEM_PROBE341
    always @ (posedge clk)
    begin
      shift_probe341 <= probe341;
      mem_shift_probe341 <= shift_probe341;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 342) begin : FF_MEM_PROBE342
    always @ (posedge clk)
    begin
      shift_probe342 <= probe342;
      mem_shift_probe342 <= shift_probe342;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 343) begin : FF_MEM_PROBE343
    always @ (posedge clk)
    begin
      shift_probe343 <= probe343;
      mem_shift_probe343 <= shift_probe343;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 344) begin : FF_MEM_PROBE344
    always @ (posedge clk)
    begin
      shift_probe344 <= probe344;
      mem_shift_probe344 <= shift_probe344;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 345) begin : FF_MEM_PROBE345
    always @ (posedge clk)
    begin
      shift_probe345 <= probe345;
      mem_shift_probe345 <= shift_probe345;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 346) begin : FF_MEM_PROBE346
    always @ (posedge clk)
    begin
      shift_probe346 <= probe346;
      mem_shift_probe346 <= shift_probe346;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 347) begin : FF_MEM_PROBE347
    always @ (posedge clk)
    begin
      shift_probe347 <= probe347;
      mem_shift_probe347 <= shift_probe347;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 348) begin : FF_MEM_PROBE348
    always @ (posedge clk)
    begin
      shift_probe348 <= probe348;
      mem_shift_probe348 <= shift_probe348;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 349) begin : FF_MEM_PROBE349
    always @ (posedge clk)
    begin
      shift_probe349 <= probe349;
      mem_shift_probe349 <= shift_probe349;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 350) begin : FF_MEM_PROBE350
    always @ (posedge clk)
    begin
      shift_probe350 <= probe350;
      mem_shift_probe350 <= shift_probe350;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 351) begin : FF_MEM_PROBE351
    always @ (posedge clk)
    begin
      shift_probe351 <= probe351;
      mem_shift_probe351 <= shift_probe351;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 352) begin : FF_MEM_PROBE352
    always @ (posedge clk)
    begin
      shift_probe352 <= probe352;
      mem_shift_probe352 <= shift_probe352;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 353) begin : FF_MEM_PROBE353
    always @ (posedge clk)
    begin
      shift_probe353 <= probe353;
      mem_shift_probe353 <= shift_probe353;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 354) begin : FF_MEM_PROBE354
    always @ (posedge clk)
    begin
      shift_probe354 <= probe354;
      mem_shift_probe354 <= shift_probe354;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 355) begin : FF_MEM_PROBE355
    always @ (posedge clk)
    begin
      shift_probe355 <= probe355;
      mem_shift_probe355 <= shift_probe355;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 356) begin : FF_MEM_PROBE356
    always @ (posedge clk)
    begin
      shift_probe356 <= probe356;
      mem_shift_probe356 <= shift_probe356;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 357) begin : FF_MEM_PROBE357
    always @ (posedge clk)
    begin
      shift_probe357 <= probe357;
      mem_shift_probe357 <= shift_probe357;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 358) begin : FF_MEM_PROBE358
    always @ (posedge clk)
    begin
      shift_probe358 <= probe358;
      mem_shift_probe358 <= shift_probe358;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 359) begin : FF_MEM_PROBE359
    always @ (posedge clk)
    begin
      shift_probe359 <= probe359;
      mem_shift_probe359 <= shift_probe359;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 360) begin : FF_MEM_PROBE360
    always @ (posedge clk)
    begin
      shift_probe360 <= probe360;
      mem_shift_probe360 <= shift_probe360;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 361) begin : FF_MEM_PROBE361
    always @ (posedge clk)
    begin
      shift_probe361 <= probe361;
      mem_shift_probe361 <= shift_probe361;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 362) begin : FF_MEM_PROBE362
    always @ (posedge clk)
    begin
      shift_probe362 <= probe362;
      mem_shift_probe362 <= shift_probe362;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 363) begin : FF_MEM_PROBE363
    always @ (posedge clk)
    begin
      shift_probe363 <= probe363;
      mem_shift_probe363 <= shift_probe363;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 364) begin : FF_MEM_PROBE364
    always @ (posedge clk)
    begin
      shift_probe364 <= probe364;
      mem_shift_probe364 <= shift_probe364;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 365) begin : FF_MEM_PROBE365
    always @ (posedge clk)
    begin
      shift_probe365 <= probe365;
      mem_shift_probe365 <= shift_probe365;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 366) begin : FF_MEM_PROBE366
    always @ (posedge clk)
    begin
      shift_probe366 <= probe366;
      mem_shift_probe366 <= shift_probe366;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 367) begin : FF_MEM_PROBE367
    always @ (posedge clk)
    begin
      shift_probe367 <= probe367;
      mem_shift_probe367 <= shift_probe367;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 368) begin : FF_MEM_PROBE368
    always @ (posedge clk)
    begin
      shift_probe368 <= probe368;
      mem_shift_probe368 <= shift_probe368;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 369) begin : FF_MEM_PROBE369
    always @ (posedge clk)
    begin
      shift_probe369 <= probe369;
      mem_shift_probe369 <= shift_probe369;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 370) begin : FF_MEM_PROBE370
    always @ (posedge clk)
    begin
      shift_probe370 <= probe370;
      mem_shift_probe370 <= shift_probe370;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 371) begin : FF_MEM_PROBE371
    always @ (posedge clk)
    begin
      shift_probe371 <= probe371;
      mem_shift_probe371 <= shift_probe371;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 372) begin : FF_MEM_PROBE372
    always @ (posedge clk)
    begin
      shift_probe372 <= probe372;
      mem_shift_probe372 <= shift_probe372;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 373) begin : FF_MEM_PROBE373
    always @ (posedge clk)
    begin
      shift_probe373 <= probe373;
      mem_shift_probe373 <= shift_probe373;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 374) begin : FF_MEM_PROBE374
    always @ (posedge clk)
    begin
      shift_probe374 <= probe374;
      mem_shift_probe374 <= shift_probe374;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 375) begin : FF_MEM_PROBE375
    always @ (posedge clk)
    begin
      shift_probe375 <= probe375;
      mem_shift_probe375 <= shift_probe375;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 376) begin : FF_MEM_PROBE376
    always @ (posedge clk)
    begin
      shift_probe376 <= probe376;
      mem_shift_probe376 <= shift_probe376;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 377) begin : FF_MEM_PROBE377
    always @ (posedge clk)
    begin
      shift_probe377 <= probe377;
      mem_shift_probe377 <= shift_probe377;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 378) begin : FF_MEM_PROBE378
    always @ (posedge clk)
    begin
      shift_probe378 <= probe378;
      mem_shift_probe378 <= shift_probe378;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 379) begin : FF_MEM_PROBE379
    always @ (posedge clk)
    begin
      shift_probe379 <= probe379;
      mem_shift_probe379 <= shift_probe379;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 380) begin : FF_MEM_PROBE380
    always @ (posedge clk)
    begin
      shift_probe380 <= probe380;
      mem_shift_probe380 <= shift_probe380;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 381) begin : FF_MEM_PROBE381
    always @ (posedge clk)
    begin
      shift_probe381 <= probe381;
      mem_shift_probe381 <= shift_probe381;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 382) begin : FF_MEM_PROBE382
    always @ (posedge clk)
    begin
      shift_probe382 <= probe382;
      mem_shift_probe382 <= shift_probe382;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 383) begin : FF_MEM_PROBE383
    always @ (posedge clk)
    begin
      shift_probe383 <= probe383;
      mem_shift_probe383 <= shift_probe383;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 384) begin : FF_MEM_PROBE384
    always @ (posedge clk)
    begin
      shift_probe384 <= probe384;
      mem_shift_probe384 <= shift_probe384;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 385) begin : FF_MEM_PROBE385
    always @ (posedge clk)
    begin
      shift_probe385 <= probe385;
      mem_shift_probe385 <= shift_probe385;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 386) begin : FF_MEM_PROBE386
    always @ (posedge clk)
    begin
      shift_probe386 <= probe386;
      mem_shift_probe386 <= shift_probe386;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 387) begin : FF_MEM_PROBE387
    always @ (posedge clk)
    begin
      shift_probe387 <= probe387;
      mem_shift_probe387 <= shift_probe387;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 388) begin : FF_MEM_PROBE388
    always @ (posedge clk)
    begin
      shift_probe388 <= probe388;
      mem_shift_probe388 <= shift_probe388;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 389) begin : FF_MEM_PROBE389
    always @ (posedge clk)
    begin
      shift_probe389 <= probe389;
      mem_shift_probe389 <= shift_probe389;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 390) begin : FF_MEM_PROBE390
    always @ (posedge clk)
    begin
      shift_probe390 <= probe390;
      mem_shift_probe390 <= shift_probe390;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 391) begin : FF_MEM_PROBE391
    always @ (posedge clk)
    begin
      shift_probe391 <= probe391;
      mem_shift_probe391 <= shift_probe391;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 392) begin : FF_MEM_PROBE392
    always @ (posedge clk)
    begin
      shift_probe392 <= probe392;
      mem_shift_probe392 <= shift_probe392;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 393) begin : FF_MEM_PROBE393
    always @ (posedge clk)
    begin
      shift_probe393 <= probe393;
      mem_shift_probe393 <= shift_probe393;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 394) begin : FF_MEM_PROBE394
    always @ (posedge clk)
    begin
      shift_probe394 <= probe394;
      mem_shift_probe394 <= shift_probe394;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 395) begin : FF_MEM_PROBE395
    always @ (posedge clk)
    begin
      shift_probe395 <= probe395;
      mem_shift_probe395 <= shift_probe395;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 396) begin : FF_MEM_PROBE396
    always @ (posedge clk)
    begin
      shift_probe396 <= probe396;
      mem_shift_probe396 <= shift_probe396;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 397) begin : FF_MEM_PROBE397
    always @ (posedge clk)
    begin
      shift_probe397 <= probe397;
      mem_shift_probe397 <= shift_probe397;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 398) begin : FF_MEM_PROBE398
    always @ (posedge clk)
    begin
      shift_probe398 <= probe398;
      mem_shift_probe398 <= shift_probe398;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 399) begin : FF_MEM_PROBE399
    always @ (posedge clk)
    begin
      shift_probe399 <= probe399;
      mem_shift_probe399 <= shift_probe399;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 400) begin : FF_MEM_PROBE400
    always @ (posedge clk)
    begin
      shift_probe400 <= probe400;
      mem_shift_probe400 <= shift_probe400;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 401) begin : FF_MEM_PROBE401
    always @ (posedge clk)
    begin
      shift_probe401 <= probe401;
      mem_shift_probe401 <= shift_probe401;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 402) begin : FF_MEM_PROBE402
    always @ (posedge clk)
    begin
      shift_probe402 <= probe402;
      mem_shift_probe402 <= shift_probe402;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 403) begin : FF_MEM_PROBE403
    always @ (posedge clk)
    begin
      shift_probe403 <= probe403;
      mem_shift_probe403 <= shift_probe403;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 404) begin : FF_MEM_PROBE404
    always @ (posedge clk)
    begin
      shift_probe404 <= probe404;
      mem_shift_probe404 <= shift_probe404;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 405) begin : FF_MEM_PROBE405
    always @ (posedge clk)
    begin
      shift_probe405 <= probe405;
      mem_shift_probe405 <= shift_probe405;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 406) begin : FF_MEM_PROBE406
    always @ (posedge clk)
    begin
      shift_probe406 <= probe406;
      mem_shift_probe406 <= shift_probe406;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 407) begin : FF_MEM_PROBE407
    always @ (posedge clk)
    begin
      shift_probe407 <= probe407;
      mem_shift_probe407 <= shift_probe407;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 408) begin : FF_MEM_PROBE408
    always @ (posedge clk)
    begin
      shift_probe408 <= probe408;
      mem_shift_probe408 <= shift_probe408;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 409) begin : FF_MEM_PROBE409
    always @ (posedge clk)
    begin
      shift_probe409 <= probe409;
      mem_shift_probe409 <= shift_probe409;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 410) begin : FF_MEM_PROBE410
    always @ (posedge clk)
    begin
      shift_probe410 <= probe410;
      mem_shift_probe410 <= shift_probe410;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 411) begin : FF_MEM_PROBE411
    always @ (posedge clk)
    begin
      shift_probe411 <= probe411;
      mem_shift_probe411 <= shift_probe411;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 412) begin : FF_MEM_PROBE412
    always @ (posedge clk)
    begin
      shift_probe412 <= probe412;
      mem_shift_probe412 <= shift_probe412;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 413) begin : FF_MEM_PROBE413
    always @ (posedge clk)
    begin
      shift_probe413 <= probe413;
      mem_shift_probe413 <= shift_probe413;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 414) begin : FF_MEM_PROBE414
    always @ (posedge clk)
    begin
      shift_probe414 <= probe414;
      mem_shift_probe414 <= shift_probe414;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 415) begin : FF_MEM_PROBE415
    always @ (posedge clk)
    begin
      shift_probe415 <= probe415;
      mem_shift_probe415 <= shift_probe415;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 416) begin : FF_MEM_PROBE416
    always @ (posedge clk)
    begin
      shift_probe416 <= probe416;
      mem_shift_probe416 <= shift_probe416;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 417) begin : FF_MEM_PROBE417
    always @ (posedge clk)
    begin
      shift_probe417 <= probe417;
      mem_shift_probe417 <= shift_probe417;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 418) begin : FF_MEM_PROBE418
    always @ (posedge clk)
    begin
      shift_probe418 <= probe418;
      mem_shift_probe418 <= shift_probe418;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 419) begin : FF_MEM_PROBE419
    always @ (posedge clk)
    begin
      shift_probe419 <= probe419;
      mem_shift_probe419 <= shift_probe419;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 420) begin : FF_MEM_PROBE420
    always @ (posedge clk)
    begin
      shift_probe420 <= probe420;
      mem_shift_probe420 <= shift_probe420;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 421) begin : FF_MEM_PROBE421
    always @ (posedge clk)
    begin
      shift_probe421 <= probe421;
      mem_shift_probe421 <= shift_probe421;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 422) begin : FF_MEM_PROBE422
    always @ (posedge clk)
    begin
      shift_probe422 <= probe422;
      mem_shift_probe422 <= shift_probe422;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 423) begin : FF_MEM_PROBE423
    always @ (posedge clk)
    begin
      shift_probe423 <= probe423;
      mem_shift_probe423 <= shift_probe423;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 424) begin : FF_MEM_PROBE424
    always @ (posedge clk)
    begin
      shift_probe424 <= probe424;
      mem_shift_probe424 <= shift_probe424;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 425) begin : FF_MEM_PROBE425
    always @ (posedge clk)
    begin
      shift_probe425 <= probe425;
      mem_shift_probe425 <= shift_probe425;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 426) begin : FF_MEM_PROBE426
    always @ (posedge clk)
    begin
      shift_probe426 <= probe426;
      mem_shift_probe426 <= shift_probe426;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 427) begin : FF_MEM_PROBE427
    always @ (posedge clk)
    begin
      shift_probe427 <= probe427;
      mem_shift_probe427 <= shift_probe427;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 428) begin : FF_MEM_PROBE428
    always @ (posedge clk)
    begin
      shift_probe428 <= probe428;
      mem_shift_probe428 <= shift_probe428;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 429) begin : FF_MEM_PROBE429
    always @ (posedge clk)
    begin
      shift_probe429 <= probe429;
      mem_shift_probe429 <= shift_probe429;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 430) begin : FF_MEM_PROBE430
    always @ (posedge clk)
    begin
      shift_probe430 <= probe430;
      mem_shift_probe430 <= shift_probe430;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 431) begin : FF_MEM_PROBE431
    always @ (posedge clk)
    begin
      shift_probe431 <= probe431;
      mem_shift_probe431 <= shift_probe431;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 432) begin : FF_MEM_PROBE432
    always @ (posedge clk)
    begin
      shift_probe432 <= probe432;
      mem_shift_probe432 <= shift_probe432;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 433) begin : FF_MEM_PROBE433
    always @ (posedge clk)
    begin
      shift_probe433 <= probe433;
      mem_shift_probe433 <= shift_probe433;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 434) begin : FF_MEM_PROBE434
    always @ (posedge clk)
    begin
      shift_probe434 <= probe434;
      mem_shift_probe434 <= shift_probe434;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 435) begin : FF_MEM_PROBE435
    always @ (posedge clk)
    begin
      shift_probe435 <= probe435;
      mem_shift_probe435 <= shift_probe435;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 436) begin : FF_MEM_PROBE436
    always @ (posedge clk)
    begin
      shift_probe436 <= probe436;
      mem_shift_probe436 <= shift_probe436;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 437) begin : FF_MEM_PROBE437
    always @ (posedge clk)
    begin
      shift_probe437 <= probe437;
      mem_shift_probe437 <= shift_probe437;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 438) begin : FF_MEM_PROBE438
    always @ (posedge clk)
    begin
      shift_probe438 <= probe438;
      mem_shift_probe438 <= shift_probe438;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 439) begin : FF_MEM_PROBE439
    always @ (posedge clk)
    begin
      shift_probe439 <= probe439;
      mem_shift_probe439 <= shift_probe439;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 440) begin : FF_MEM_PROBE440
    always @ (posedge clk)
    begin
      shift_probe440 <= probe440;
      mem_shift_probe440 <= shift_probe440;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 441) begin : FF_MEM_PROBE441
    always @ (posedge clk)
    begin
      shift_probe441 <= probe441;
      mem_shift_probe441 <= shift_probe441;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 442) begin : FF_MEM_PROBE442
    always @ (posedge clk)
    begin
      shift_probe442 <= probe442;
      mem_shift_probe442 <= shift_probe442;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 443) begin : FF_MEM_PROBE443
    always @ (posedge clk)
    begin
      shift_probe443 <= probe443;
      mem_shift_probe443 <= shift_probe443;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 444) begin : FF_MEM_PROBE444
    always @ (posedge clk)
    begin
      shift_probe444 <= probe444;
      mem_shift_probe444 <= shift_probe444;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 445) begin : FF_MEM_PROBE445
    always @ (posedge clk)
    begin
      shift_probe445 <= probe445;
      mem_shift_probe445 <= shift_probe445;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 446) begin : FF_MEM_PROBE446
    always @ (posedge clk)
    begin
      shift_probe446 <= probe446;
      mem_shift_probe446 <= shift_probe446;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 447) begin : FF_MEM_PROBE447
    always @ (posedge clk)
    begin
      shift_probe447 <= probe447;
      mem_shift_probe447 <= shift_probe447;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 448) begin : FF_MEM_PROBE448
    always @ (posedge clk)
    begin
      shift_probe448 <= probe448;
      mem_shift_probe448 <= shift_probe448;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 449) begin : FF_MEM_PROBE449
    always @ (posedge clk)
    begin
      shift_probe449 <= probe449;
      mem_shift_probe449 <= shift_probe449;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 450) begin : FF_MEM_PROBE450
    always @ (posedge clk)
    begin
      shift_probe450 <= probe450;
      mem_shift_probe450 <= shift_probe450;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 451) begin : FF_MEM_PROBE451
    always @ (posedge clk)
    begin
      shift_probe451 <= probe451;
      mem_shift_probe451 <= shift_probe451;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 452) begin : FF_MEM_PROBE452
    always @ (posedge clk)
    begin
      shift_probe452 <= probe452;
      mem_shift_probe452 <= shift_probe452;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 453) begin : FF_MEM_PROBE453
    always @ (posedge clk)
    begin
      shift_probe453 <= probe453;
      mem_shift_probe453 <= shift_probe453;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 454) begin : FF_MEM_PROBE454
    always @ (posedge clk)
    begin
      shift_probe454 <= probe454;
      mem_shift_probe454 <= shift_probe454;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 455) begin : FF_MEM_PROBE455
    always @ (posedge clk)
    begin
      shift_probe455 <= probe455;
      mem_shift_probe455 <= shift_probe455;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 456) begin : FF_MEM_PROBE456
    always @ (posedge clk)
    begin
      shift_probe456 <= probe456;
      mem_shift_probe456 <= shift_probe456;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 457) begin : FF_MEM_PROBE457
    always @ (posedge clk)
    begin
      shift_probe457 <= probe457;
      mem_shift_probe457 <= shift_probe457;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 458) begin : FF_MEM_PROBE458
    always @ (posedge clk)
    begin
      shift_probe458 <= probe458;
      mem_shift_probe458 <= shift_probe458;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 459) begin : FF_MEM_PROBE459
    always @ (posedge clk)
    begin
      shift_probe459 <= probe459;
      mem_shift_probe459 <= shift_probe459;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 460) begin : FF_MEM_PROBE460
    always @ (posedge clk)
    begin
      shift_probe460 <= probe460;
      mem_shift_probe460 <= shift_probe460;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 461) begin : FF_MEM_PROBE461
    always @ (posedge clk)
    begin
      shift_probe461 <= probe461;
      mem_shift_probe461 <= shift_probe461;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 462) begin : FF_MEM_PROBE462
    always @ (posedge clk)
    begin
      shift_probe462 <= probe462;
      mem_shift_probe462 <= shift_probe462;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 463) begin : FF_MEM_PROBE463
    always @ (posedge clk)
    begin
      shift_probe463 <= probe463;
      mem_shift_probe463 <= shift_probe463;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 464) begin : FF_MEM_PROBE464
    always @ (posedge clk)
    begin
      shift_probe464 <= probe464;
      mem_shift_probe464 <= shift_probe464;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 465) begin : FF_MEM_PROBE465
    always @ (posedge clk)
    begin
      shift_probe465 <= probe465;
      mem_shift_probe465 <= shift_probe465;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 466) begin : FF_MEM_PROBE466
    always @ (posedge clk)
    begin
      shift_probe466 <= probe466;
      mem_shift_probe466 <= shift_probe466;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 467) begin : FF_MEM_PROBE467
    always @ (posedge clk)
    begin
      shift_probe467 <= probe467;
      mem_shift_probe467 <= shift_probe467;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 468) begin : FF_MEM_PROBE468
    always @ (posedge clk)
    begin
      shift_probe468 <= probe468;
      mem_shift_probe468 <= shift_probe468;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 469) begin : FF_MEM_PROBE469
    always @ (posedge clk)
    begin
      shift_probe469 <= probe469;
      mem_shift_probe469 <= shift_probe469;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 470) begin : FF_MEM_PROBE470
    always @ (posedge clk)
    begin
      shift_probe470 <= probe470;
      mem_shift_probe470 <= shift_probe470;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 471) begin : FF_MEM_PROBE471
    always @ (posedge clk)
    begin
      shift_probe471 <= probe471;
      mem_shift_probe471 <= shift_probe471;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 472) begin : FF_MEM_PROBE472
    always @ (posedge clk)
    begin
      shift_probe472 <= probe472;
      mem_shift_probe472 <= shift_probe472;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 473) begin : FF_MEM_PROBE473
    always @ (posedge clk)
    begin
      shift_probe473 <= probe473;
      mem_shift_probe473 <= shift_probe473;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 474) begin : FF_MEM_PROBE474
    always @ (posedge clk)
    begin
      shift_probe474 <= probe474;
      mem_shift_probe474 <= shift_probe474;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 475) begin : FF_MEM_PROBE475
    always @ (posedge clk)
    begin
      shift_probe475 <= probe475;
      mem_shift_probe475 <= shift_probe475;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 476) begin : FF_MEM_PROBE476
    always @ (posedge clk)
    begin
      shift_probe476 <= probe476;
      mem_shift_probe476 <= shift_probe476;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 477) begin : FF_MEM_PROBE477
    always @ (posedge clk)
    begin
      shift_probe477 <= probe477;
      mem_shift_probe477 <= shift_probe477;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 478) begin : FF_MEM_PROBE478
    always @ (posedge clk)
    begin
      shift_probe478 <= probe478;
      mem_shift_probe478 <= shift_probe478;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 479) begin : FF_MEM_PROBE479
    always @ (posedge clk)
    begin
      shift_probe479 <= probe479;
      mem_shift_probe479 <= shift_probe479;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 480) begin : FF_MEM_PROBE480
    always @ (posedge clk)
    begin
      shift_probe480 <= probe480;
      mem_shift_probe480 <= shift_probe480;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 481) begin : FF_MEM_PROBE481
    always @ (posedge clk)
    begin
      shift_probe481 <= probe481;
      mem_shift_probe481 <= shift_probe481;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 482) begin : FF_MEM_PROBE482
    always @ (posedge clk)
    begin
      shift_probe482 <= probe482;
      mem_shift_probe482 <= shift_probe482;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 483) begin : FF_MEM_PROBE483
    always @ (posedge clk)
    begin
      shift_probe483 <= probe483;
      mem_shift_probe483 <= shift_probe483;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 484) begin : FF_MEM_PROBE484
    always @ (posedge clk)
    begin
      shift_probe484 <= probe484;
      mem_shift_probe484 <= shift_probe484;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 485) begin : FF_MEM_PROBE485
    always @ (posedge clk)
    begin
      shift_probe485 <= probe485;
      mem_shift_probe485 <= shift_probe485;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 486) begin : FF_MEM_PROBE486
    always @ (posedge clk)
    begin
      shift_probe486 <= probe486;
      mem_shift_probe486 <= shift_probe486;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 487) begin : FF_MEM_PROBE487
    always @ (posedge clk)
    begin
      shift_probe487 <= probe487;
      mem_shift_probe487 <= shift_probe487;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 488) begin : FF_MEM_PROBE488
    always @ (posedge clk)
    begin
      shift_probe488 <= probe488;
      mem_shift_probe488 <= shift_probe488;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 489) begin : FF_MEM_PROBE489
    always @ (posedge clk)
    begin
      shift_probe489 <= probe489;
      mem_shift_probe489 <= shift_probe489;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 490) begin : FF_MEM_PROBE490
    always @ (posedge clk)
    begin
      shift_probe490 <= probe490;
      mem_shift_probe490 <= shift_probe490;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 491) begin : FF_MEM_PROBE491
    always @ (posedge clk)
    begin
      shift_probe491 <= probe491;
      mem_shift_probe491 <= shift_probe491;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 492) begin : FF_MEM_PROBE492
    always @ (posedge clk)
    begin
      shift_probe492 <= probe492;
      mem_shift_probe492 <= shift_probe492;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 493) begin : FF_MEM_PROBE493
    always @ (posedge clk)
    begin
      shift_probe493 <= probe493;
      mem_shift_probe493 <= shift_probe493;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 494) begin : FF_MEM_PROBE494
    always @ (posedge clk)
    begin
      shift_probe494 <= probe494;
      mem_shift_probe494 <= shift_probe494;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 495) begin : FF_MEM_PROBE495
    always @ (posedge clk)
    begin
      shift_probe495 <= probe495;
      mem_shift_probe495 <= shift_probe495;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 496) begin : FF_MEM_PROBE496
    always @ (posedge clk)
    begin
      shift_probe496 <= probe496;
      mem_shift_probe496 <= shift_probe496;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 497) begin : FF_MEM_PROBE497
    always @ (posedge clk)
    begin
      shift_probe497 <= probe497;
      mem_shift_probe497 <= shift_probe497;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 498) begin : FF_MEM_PROBE498
    always @ (posedge clk)
    begin
      shift_probe498 <= probe498;
      mem_shift_probe498 <= shift_probe498;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 499) begin : FF_MEM_PROBE499
    always @ (posedge clk)
    begin
      shift_probe499 <= probe499;
      mem_shift_probe499 <= shift_probe499;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 500) begin : FF_MEM_PROBE500
    always @ (posedge clk)
    begin
      shift_probe500 <= probe500;
      mem_shift_probe500 <= shift_probe500;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 501) begin : FF_MEM_PROBE501
    always @ (posedge clk)
    begin
      shift_probe501 <= probe501;
      mem_shift_probe501 <= shift_probe501;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 502) begin : FF_MEM_PROBE502
    always @ (posedge clk)
    begin
      shift_probe502 <= probe502;
      mem_shift_probe502 <= shift_probe502;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 503) begin : FF_MEM_PROBE503
    always @ (posedge clk)
    begin
      shift_probe503 <= probe503;
      mem_shift_probe503 <= shift_probe503;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 504) begin : FF_MEM_PROBE504
    always @ (posedge clk)
    begin
      shift_probe504 <= probe504;
      mem_shift_probe504 <= shift_probe504;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 505) begin : FF_MEM_PROBE505
    always @ (posedge clk)
    begin
      shift_probe505 <= probe505;
      mem_shift_probe505 <= shift_probe505;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 506) begin : FF_MEM_PROBE506
    always @ (posedge clk)
    begin
      shift_probe506 <= probe506;
      mem_shift_probe506 <= shift_probe506;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 507) begin : FF_MEM_PROBE507
    always @ (posedge clk)
    begin
      shift_probe507 <= probe507;
      mem_shift_probe507 <= shift_probe507;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 508) begin : FF_MEM_PROBE508
    always @ (posedge clk)
    begin
      shift_probe508 <= probe508;
      mem_shift_probe508 <= shift_probe508;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 509) begin : FF_MEM_PROBE509
    always @ (posedge clk)
    begin
      shift_probe509 <= probe509;
      mem_shift_probe509 <= shift_probe509;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 510) begin : FF_MEM_PROBE510
    always @ (posedge clk)
    begin
      shift_probe510 <= probe510;
      mem_shift_probe510 <= shift_probe510;
    end
  end
endgenerate
generate
  if (C_NUM_PROBES > 511) begin : FF_MEM_PROBE511
    always @ (posedge clk)
    begin
      shift_probe511 <= probe511;
      mem_shift_probe511 <= shift_probe511;
    end
  end
endgenerate


generate 
  if (C_NUM_PROBES == 1) begin : MEM_DAT_1
   assign mem_data_i = {mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 2) begin : MEM_DATA_2
    assign mem_data_i = {mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 3) begin : MEM_DATA_3
    assign mem_data_i = {mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 4) begin : MEM_DATA_4
    assign mem_data_i = {mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 5) begin : MEM_DATA_5
    assign mem_data_i = {mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 6) begin : MEM_DATA_6
    assign mem_data_i = {mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 7) begin : MEM_DATA_7
    assign mem_data_i = {mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 8) begin : MEM_DATA_8
    assign mem_data_i = {mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 9) begin : MEM_DATA_9
    assign mem_data_i = {mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 10) begin : MEM_DATA_10
    assign mem_data_i = {mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 11) begin : MEM_DATA_11
    assign mem_data_i = {mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 12) begin : MEM_DATA_12
    assign mem_data_i = {mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 13) begin : MEM_DATA_13
    assign mem_data_i = {mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 14) begin : MEM_DATA_14
    assign mem_data_i = {mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 15) begin : MEM_DATA_15
    assign mem_data_i = {mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 16) begin : MEM_DATA_16
    assign mem_data_i = {mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 17) begin : MEM_DATA_17
    assign mem_data_i = {mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 18) begin : MEM_DATA_18
    assign mem_data_i = {mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 19) begin : MEM_DATA_19
    assign mem_data_i = {mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 20) begin : MEM_DATA_20
    assign mem_data_i = {mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 21) begin : MEM_DATA_21
    assign mem_data_i = {mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 22) begin : MEM_DATA_22
    assign mem_data_i = {mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 23) begin : MEM_DATA_23
    assign mem_data_i = {mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 24) begin : MEM_DATA_24
    assign mem_data_i = {mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 25) begin : MEM_DATA_25
    assign mem_data_i = {mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 26) begin : MEM_DATA_26
    assign mem_data_i = {mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 27) begin : MEM_DATA_27
    assign mem_data_i = {mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 28) begin : MEM_DATA_28
    assign mem_data_i = {mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 29) begin : MEM_DATA_29
    assign mem_data_i = {mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 30) begin : MEM_DATA_30
    assign mem_data_i = {mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 31) begin : MEM_DATA_31
    assign mem_data_i = {mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 32) begin : MEM_DATA_32
    assign mem_data_i = {mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 33) begin : MEM_DATA_33
    assign mem_data_i = {mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 34) begin : MEM_DATA_34
    assign mem_data_i = {mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 35) begin : MEM_DATA_35
    assign mem_data_i = {mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 36) begin : MEM_DATA_36
    assign mem_data_i = {mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 37) begin : MEM_DATA_37
    assign mem_data_i = {mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 38) begin : MEM_DATA_38
    assign mem_data_i = {mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 39) begin : MEM_DATA_39
    assign mem_data_i = {mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 40) begin : MEM_DATA_40
    assign mem_data_i = {mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 41) begin : MEM_DATA_41
    assign mem_data_i = {mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 42) begin : MEM_DATA_42
    assign mem_data_i = {mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 43) begin : MEM_DATA_43
    assign mem_data_i = {mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 44) begin : MEM_DATA_44
    assign mem_data_i = {mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 45) begin : MEM_DATA_45
    assign mem_data_i = {mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 46) begin : MEM_DATA_46
    assign mem_data_i = {mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 47) begin : MEM_DATA_47
    assign mem_data_i = {mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 48) begin : MEM_DATA_48
    assign mem_data_i = {mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 49) begin : MEM_DATA_49
    assign mem_data_i = {mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 50) begin : MEM_DATA_50
    assign mem_data_i = {mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 51) begin : MEM_DATA_51
    assign mem_data_i = {mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 52) begin : MEM_DATA_52
    assign mem_data_i = {mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 53) begin : MEM_DATA_53
    assign mem_data_i = {mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 54) begin : MEM_DATA_54
    assign mem_data_i = {mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 55) begin : MEM_DATA_55
    assign mem_data_i = {mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 56) begin : MEM_DATA_56
    assign mem_data_i = {mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 57) begin : MEM_DATA_57
    assign mem_data_i = {mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 58) begin : MEM_DATA_58
    assign mem_data_i = {mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 59) begin : MEM_DATA_59
    assign mem_data_i = {mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 60) begin : MEM_DATA_60
    assign mem_data_i = {mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 61) begin : MEM_DATA_61
    assign mem_data_i = {mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 62) begin : MEM_DATA_62
    assign mem_data_i = {mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 63) begin : MEM_DATA_63
    assign mem_data_i = {mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 64) begin : MEM_DATA_64
    assign mem_data_i = {mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 65) begin : MEM_DATA_65
    assign mem_data_i = {mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 66) begin : MEM_DATA_66
    assign mem_data_i = {mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 67) begin : MEM_DATA_67
    assign mem_data_i = {mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 68) begin : MEM_DATA_68
    assign mem_data_i = {mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 69) begin : MEM_DATA_69
    assign mem_data_i = {mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 70) begin : MEM_DATA_70
    assign mem_data_i = {mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 71) begin : MEM_DATA_71
    assign mem_data_i = {mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 72) begin : MEM_DATA_72
    assign mem_data_i = {mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 73) begin : MEM_DATA_73
    assign mem_data_i = {mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 74) begin : MEM_DATA_74
    assign mem_data_i = {mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 75) begin : MEM_DATA_75
    assign mem_data_i = {mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 76) begin : MEM_DATA_76
    assign mem_data_i = {mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 77) begin : MEM_DATA_77
    assign mem_data_i = {mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 78) begin : MEM_DATA_78
    assign mem_data_i = {mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 79) begin : MEM_DATA_79
    assign mem_data_i = {mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 80) begin : MEM_DATA_80
    assign mem_data_i = {mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 81) begin : MEM_DATA_81
    assign mem_data_i = {mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 82) begin : MEM_DATA_82
    assign mem_data_i = {mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 83) begin : MEM_DATA_83
    assign mem_data_i = {mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 84) begin : MEM_DATA_84
    assign mem_data_i = {mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 85) begin : MEM_DATA_85
    assign mem_data_i = {mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 86) begin : MEM_DATA_86
    assign mem_data_i = {mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 87) begin : MEM_DATA_87
    assign mem_data_i = {mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 88) begin : MEM_DATA_88
    assign mem_data_i = {mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 89) begin : MEM_DATA_89
    assign mem_data_i = {mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 90) begin : MEM_DATA_90
    assign mem_data_i = {mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 91) begin : MEM_DATA_91
    assign mem_data_i = {mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 92) begin : MEM_DATA_92
    assign mem_data_i = {mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 93) begin : MEM_DATA_93
    assign mem_data_i = {mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 94) begin : MEM_DATA_94
    assign mem_data_i = {mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 95) begin : MEM_DATA_95
    assign mem_data_i = {mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 96) begin : MEM_DATA_96
    assign mem_data_i = {mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 97) begin : MEM_DATA_97
    assign mem_data_i = {mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 98) begin : MEM_DATA_98
    assign mem_data_i = {mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 99) begin : MEM_DATA_99
    assign mem_data_i = {mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 100) begin : MEM_DATA_100
    assign mem_data_i = {mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 101) begin : MEM_DATA_101
    assign mem_data_i = {mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 102) begin : MEM_DATA_102
    assign mem_data_i = {mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 103) begin : MEM_DATA_103
    assign mem_data_i = {mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 104) begin : MEM_DATA_104
    assign mem_data_i = {mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 105) begin : MEM_DATA_105
    assign mem_data_i = {mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 106) begin : MEM_DATA_106
    assign mem_data_i = {mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 107) begin : MEM_DATA_107
    assign mem_data_i = {mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 108) begin : MEM_DATA_108
    assign mem_data_i = {mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 109) begin : MEM_DATA_109
    assign mem_data_i = {mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 110) begin : MEM_DATA_110
    assign mem_data_i = {mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 111) begin : MEM_DATA_111
    assign mem_data_i = {mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 112) begin : MEM_DATA_112
    assign mem_data_i = {mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 113) begin : MEM_DATA_113
    assign mem_data_i = {mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 114) begin : MEM_DATA_114
    assign mem_data_i = {mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 115) begin : MEM_DATA_115
    assign mem_data_i = {mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 116) begin : MEM_DATA_116
    assign mem_data_i = {mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 117) begin : MEM_DATA_117
    assign mem_data_i = {mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 118) begin : MEM_DATA_118
    assign mem_data_i = {mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 119) begin : MEM_DATA_119
    assign mem_data_i = {mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 120) begin : MEM_DATA_120
    assign mem_data_i = {mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 121) begin : MEM_DATA_121
    assign mem_data_i = {mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 122) begin : MEM_DATA_122
    assign mem_data_i = {mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 123) begin : MEM_DATA_123
    assign mem_data_i = {mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 124) begin : MEM_DATA_124
    assign mem_data_i = {mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 125) begin : MEM_DATA_125
    assign mem_data_i = {mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 126) begin : MEM_DATA_126
    assign mem_data_i = {mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 127) begin : MEM_DATA_127
    assign mem_data_i = {mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 128) begin : MEM_DATA_128
    assign mem_data_i = {mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 129) begin : MEM_DATA_129
    assign mem_data_i = {mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 130) begin : MEM_DATA_130
    assign mem_data_i = {mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 131) begin : MEM_DATA_131
    assign mem_data_i = {mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 132) begin : MEM_DATA_132
    assign mem_data_i = {mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 133) begin : MEM_DATA_133
    assign mem_data_i = {mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 134) begin : MEM_DATA_134
    assign mem_data_i = {mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 135) begin : MEM_DATA_135
    assign mem_data_i = {mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 136) begin : MEM_DATA_136
    assign mem_data_i = {mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 137) begin : MEM_DATA_137
    assign mem_data_i = {mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 138) begin : MEM_DATA_138
    assign mem_data_i = {mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 139) begin : MEM_DATA_139
    assign mem_data_i = {mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 140) begin : MEM_DATA_140
    assign mem_data_i = {mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 141) begin : MEM_DATA_141
    assign mem_data_i = {mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 142) begin : MEM_DATA_142
    assign mem_data_i = {mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 143) begin : MEM_DATA_143
    assign mem_data_i = {mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 144) begin : MEM_DATA_144
    assign mem_data_i = {mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 145) begin : MEM_DATA_145
    assign mem_data_i = {mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 146) begin : MEM_DATA_146
    assign mem_data_i = {mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 147) begin : MEM_DATA_147
    assign mem_data_i = {mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 148) begin : MEM_DATA_148
    assign mem_data_i = {mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 149) begin : MEM_DATA_149
    assign mem_data_i = {mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 150) begin : MEM_DATA_150
    assign mem_data_i = {mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 151) begin : MEM_DATA_151
    assign mem_data_i = {mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 152) begin : MEM_DATA_152
    assign mem_data_i = {mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 153) begin : MEM_DATA_153
    assign mem_data_i = {mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 154) begin : MEM_DATA_154
    assign mem_data_i = {mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 155) begin : MEM_DATA_155
    assign mem_data_i = {mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 156) begin : MEM_DATA_156
    assign mem_data_i = {mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 157) begin : MEM_DATA_157
    assign mem_data_i = {mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 158) begin : MEM_DATA_158
    assign mem_data_i = {mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 159) begin : MEM_DATA_159
    assign mem_data_i = {mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 160) begin : MEM_DATA_160
    assign mem_data_i = {mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 161) begin : MEM_DATA_161
    assign mem_data_i = {mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 162) begin : MEM_DATA_162
    assign mem_data_i = {mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 163) begin : MEM_DATA_163
    assign mem_data_i = {mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 164) begin : MEM_DATA_164
    assign mem_data_i = {mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 165) begin : MEM_DATA_165
    assign mem_data_i = {mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 166) begin : MEM_DATA_166
    assign mem_data_i = {mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 167) begin : MEM_DATA_167
    assign mem_data_i = {mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 168) begin : MEM_DATA_168
    assign mem_data_i = {mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 169) begin : MEM_DATA_169
    assign mem_data_i = {mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 170) begin : MEM_DATA_170
    assign mem_data_i = {mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 171) begin : MEM_DATA_171
    assign mem_data_i = {mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 172) begin : MEM_DATA_172
    assign mem_data_i = {mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 173) begin : MEM_DATA_173
    assign mem_data_i = {mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 174) begin : MEM_DATA_174
    assign mem_data_i = {mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 175) begin : MEM_DATA_175
    assign mem_data_i = {mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 176) begin : MEM_DATA_176
    assign mem_data_i = {mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 177) begin : MEM_DATA_177
    assign mem_data_i = {mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 178) begin : MEM_DATA_178
    assign mem_data_i = {mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 179) begin : MEM_DATA_179
    assign mem_data_i = {mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 180) begin : MEM_DATA_180
    assign mem_data_i = {mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 181) begin : MEM_DATA_181
    assign mem_data_i = {mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 182) begin : MEM_DATA_182
    assign mem_data_i = {mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 183) begin : MEM_DATA_183
    assign mem_data_i = {mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 184) begin : MEM_DATA_184
    assign mem_data_i = {mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 185) begin : MEM_DATA_185
    assign mem_data_i = {mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 186) begin : MEM_DATA_186
    assign mem_data_i = {mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 187) begin : MEM_DATA_187
    assign mem_data_i = {mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 188) begin : MEM_DATA_188
    assign mem_data_i = {mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 189) begin : MEM_DATA_189
    assign mem_data_i = {mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 190) begin : MEM_DATA_190
    assign mem_data_i = {mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 191) begin : MEM_DATA_191
    assign mem_data_i = {mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 192) begin : MEM_DATA_192
    assign mem_data_i = {mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 193) begin : MEM_DATA_193
    assign mem_data_i = {mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 194) begin : MEM_DATA_194
    assign mem_data_i = {mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 195) begin : MEM_DATA_195
    assign mem_data_i = {mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 196) begin : MEM_DATA_196
    assign mem_data_i = {mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 197) begin : MEM_DATA_197
    assign mem_data_i = {mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 198) begin : MEM_DATA_198
    assign mem_data_i = {mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 199) begin : MEM_DATA_199
    assign mem_data_i = {mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 200) begin : MEM_DATA_200
    assign mem_data_i = {mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 201) begin : MEM_DATA_201
    assign mem_data_i = {mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 202) begin : MEM_DATA_202
    assign mem_data_i = {mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 203) begin : MEM_DATA_203
    assign mem_data_i = {mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 204) begin : MEM_DATA_204
    assign mem_data_i = {mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 205) begin : MEM_DATA_205
    assign mem_data_i = {mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 206) begin : MEM_DATA_206
    assign mem_data_i = {mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 207) begin : MEM_DATA_207
    assign mem_data_i = {mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 208) begin : MEM_DATA_208
    assign mem_data_i = {mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 209) begin : MEM_DATA_209
    assign mem_data_i = {mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 210) begin : MEM_DATA_210
    assign mem_data_i = {mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 211) begin : MEM_DATA_211
    assign mem_data_i = {mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 212) begin : MEM_DATA_212
    assign mem_data_i = {mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 213) begin : MEM_DATA_213
    assign mem_data_i = {mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 214) begin : MEM_DATA_214
    assign mem_data_i = {mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 215) begin : MEM_DATA_215
    assign mem_data_i = {mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 216) begin : MEM_DATA_216
    assign mem_data_i = {mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 217) begin : MEM_DATA_217
    assign mem_data_i = {mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 218) begin : MEM_DATA_218
    assign mem_data_i = {mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 219) begin : MEM_DATA_219
    assign mem_data_i = {mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 220) begin : MEM_DATA_220
    assign mem_data_i = {mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 221) begin : MEM_DATA_221
    assign mem_data_i = {mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 222) begin : MEM_DATA_222
    assign mem_data_i = {mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 223) begin : MEM_DATA_223
    assign mem_data_i = {mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 224) begin : MEM_DATA_224
    assign mem_data_i = {mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 225) begin : MEM_DATA_225
    assign mem_data_i = {mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 226) begin : MEM_DATA_226
    assign mem_data_i = {mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 227) begin : MEM_DATA_227
    assign mem_data_i = {mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 228) begin : MEM_DATA_228
    assign mem_data_i = {mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 229) begin : MEM_DATA_229
    assign mem_data_i = {mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 230) begin : MEM_DATA_230
    assign mem_data_i = {mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1,
mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 231) begin : MEM_DATA_231
    assign mem_data_i = {mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2,
mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 232) begin : MEM_DATA_232
    assign mem_data_i = {mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3,
mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 233) begin : MEM_DATA_233
    assign mem_data_i = {mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4,
mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 234) begin : MEM_DATA_234
    assign mem_data_i = {mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5,
mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 235) begin : MEM_DATA_235
    assign mem_data_i = {mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6,
mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 236) begin : MEM_DATA_236
    assign mem_data_i = {mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7,
mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 237) begin : MEM_DATA_237
    assign mem_data_i = {mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8,
mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 238) begin : MEM_DATA_238
    assign mem_data_i = {mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9,
mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 239) begin : MEM_DATA_239
    assign mem_data_i = {mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10,
mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 240) begin : MEM_DATA_240
    assign mem_data_i = {mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11,
mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 241) begin : MEM_DATA_241
    assign mem_data_i = {mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12,
mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 242) begin : MEM_DATA_242
    assign mem_data_i = {mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14,
mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 243) begin : MEM_DATA_243
    assign mem_data_i = {mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15,
mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 244) begin : MEM_DATA_244
    assign mem_data_i = {mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16,
mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 245) begin : MEM_DATA_245
    assign mem_data_i = {mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17,
mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 246) begin : MEM_DATA_246
    assign mem_data_i = {mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18,
mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 247) begin : MEM_DATA_247
    assign mem_data_i = {mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19,
mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 248) begin : MEM_DATA_248
    assign mem_data_i = {mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20,
mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 249) begin : MEM_DATA_249
    assign mem_data_i = {mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21,
mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 250) begin : MEM_DATA_250
    assign mem_data_i = {mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22,
mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 251) begin : MEM_DATA_251
    assign mem_data_i = {mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23,
mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 252) begin : MEM_DATA_252
    assign mem_data_i = {mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24,
mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 253) begin : MEM_DATA_253
    assign mem_data_i = {mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25,
mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 254) begin : MEM_DATA_254
    assign mem_data_i = {mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26,
mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 255) begin : MEM_DATA_255
    assign mem_data_i = {mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27,
mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 256) begin : MEM_DATA_256
    assign mem_data_i = {mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28,
mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 257) begin : MEM_DATA_257
    assign mem_data_i = {mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29,
mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 258) begin : MEM_DATA_258
    assign mem_data_i = {mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30,
mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 259) begin : MEM_DATA_259
    assign mem_data_i = {mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31,
mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 260) begin : MEM_DATA_260
    assign mem_data_i = {mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32,
mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 261) begin : MEM_DATA_261
    assign mem_data_i = {mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34,
mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 262) begin : MEM_DATA_262
    assign mem_data_i = {mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35,
mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 263) begin : MEM_DATA_263
    assign mem_data_i = {mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36,
mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 264) begin : MEM_DATA_264
    assign mem_data_i = {mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37,
mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 265) begin : MEM_DATA_265
    assign mem_data_i = {mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38,
mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 266) begin : MEM_DATA_266
    assign mem_data_i = {mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39,
mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 267) begin : MEM_DATA_267
    assign mem_data_i = {mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40,
mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 268) begin : MEM_DATA_268
    assign mem_data_i = {mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41,
mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 269) begin : MEM_DATA_269
    assign mem_data_i = {mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42,
mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 270) begin : MEM_DATA_270
    assign mem_data_i = {mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43,
mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 271) begin : MEM_DATA_271
    assign mem_data_i = {mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44,
mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 272) begin : MEM_DATA_272
    assign mem_data_i = {mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45,
mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 273) begin : MEM_DATA_273
    assign mem_data_i = {mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46,
mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 274) begin : MEM_DATA_274
    assign mem_data_i = {mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47,
mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 275) begin : MEM_DATA_275
    assign mem_data_i = {mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48,
mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 276) begin : MEM_DATA_276
    assign mem_data_i = {mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49,
mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 277) begin : MEM_DATA_277
    assign mem_data_i = {mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50,
mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 278) begin : MEM_DATA_278
    assign mem_data_i = {mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51,
mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 279) begin : MEM_DATA_279
    assign mem_data_i = {mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52,
mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 280) begin : MEM_DATA_280
    assign mem_data_i = {mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54,
mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 281) begin : MEM_DATA_281
    assign mem_data_i = {mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55,
mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 282) begin : MEM_DATA_282
    assign mem_data_i = {mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56,
mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 283) begin : MEM_DATA_283
    assign mem_data_i = {mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57,
mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 284) begin : MEM_DATA_284
    assign mem_data_i = {mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58,
mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 285) begin : MEM_DATA_285
    assign mem_data_i = {mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59,
mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 286) begin : MEM_DATA_286
    assign mem_data_i = {mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60,
mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 287) begin : MEM_DATA_287
    assign mem_data_i = {mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61,
mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 288) begin : MEM_DATA_288
    assign mem_data_i = {mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62,
mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 289) begin : MEM_DATA_289
    assign mem_data_i = {mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63,
mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 290) begin : MEM_DATA_290
    assign mem_data_i = {mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64,
mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 291) begin : MEM_DATA_291
    assign mem_data_i = {mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65,
mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 292) begin : MEM_DATA_292
    assign mem_data_i = {mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66,
mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 293) begin : MEM_DATA_293
    assign mem_data_i = {mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67,
mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 294) begin : MEM_DATA_294
    assign mem_data_i = {mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68,
mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 295) begin : MEM_DATA_295
    assign mem_data_i = {mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69,
mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 296) begin : MEM_DATA_296
    assign mem_data_i = {mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70,
mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 297) begin : MEM_DATA_297
    assign mem_data_i = {mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71,
mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 298) begin : MEM_DATA_298
    assign mem_data_i = {mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72,
mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 299) begin : MEM_DATA_299
    assign mem_data_i = {mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74,
mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 300) begin : MEM_DATA_300
    assign mem_data_i = {mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75,
mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 301) begin : MEM_DATA_301
    assign mem_data_i = {mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76,
mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 302) begin : MEM_DATA_302
    assign mem_data_i = {mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77,
mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 303) begin : MEM_DATA_303
    assign mem_data_i = {mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78,
mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 304) begin : MEM_DATA_304
    assign mem_data_i = {mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79,
mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 305) begin : MEM_DATA_305
    assign mem_data_i = {mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80,
mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 306) begin : MEM_DATA_306
    assign mem_data_i = {mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81,
mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 307) begin : MEM_DATA_307
    assign mem_data_i = {mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82,
mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 308) begin : MEM_DATA_308
    assign mem_data_i = {mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83,
mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 309) begin : MEM_DATA_309
    assign mem_data_i = {mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84,
mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 310) begin : MEM_DATA_310
    assign mem_data_i = {mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85,
mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 311) begin : MEM_DATA_311
    assign mem_data_i = {mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86,
mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 312) begin : MEM_DATA_312
    assign mem_data_i = {mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87,
mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 313) begin : MEM_DATA_313
    assign mem_data_i = {mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88,
mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 314) begin : MEM_DATA_314
    assign mem_data_i = {mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89,
mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 315) begin : MEM_DATA_315
    assign mem_data_i = {mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90,
mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 316) begin : MEM_DATA_316
    assign mem_data_i = {mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91,
mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 317) begin : MEM_DATA_317
    assign mem_data_i = {mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92,
mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 318) begin : MEM_DATA_318
    assign mem_data_i = {mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94,
mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 319) begin : MEM_DATA_319
    assign mem_data_i = {mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95,
mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 320) begin : MEM_DATA_320
    assign mem_data_i = {mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96,
mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 321) begin : MEM_DATA_321
    assign mem_data_i = {mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97,
mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 322) begin : MEM_DATA_322
    assign mem_data_i = {mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98,
mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 323) begin : MEM_DATA_323
    assign mem_data_i = {mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99,
mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 324) begin : MEM_DATA_324
    assign mem_data_i = {mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100,
mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 325) begin : MEM_DATA_325
    assign mem_data_i = {mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101,
mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 326) begin : MEM_DATA_326
    assign mem_data_i = {mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102,
mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 327) begin : MEM_DATA_327
    assign mem_data_i = {mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103,
mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 328) begin : MEM_DATA_328
    assign mem_data_i = {mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104,
mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 329) begin : MEM_DATA_329
    assign mem_data_i = {mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105,
mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 330) begin : MEM_DATA_330
    assign mem_data_i = {mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106,
mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 331) begin : MEM_DATA_331
    assign mem_data_i = {mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107,
mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 332) begin : MEM_DATA_332
    assign mem_data_i = {mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108,
mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 333) begin : MEM_DATA_333
    assign mem_data_i = {mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109,
mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 334) begin : MEM_DATA_334
    assign mem_data_i = {mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110,
mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 335) begin : MEM_DATA_335
    assign mem_data_i = {mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111,
mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 336) begin : MEM_DATA_336
    assign mem_data_i = {mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112,
mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 337) begin : MEM_DATA_337
    assign mem_data_i = {mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113,
mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 338) begin : MEM_DATA_338
    assign mem_data_i = {mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114,
mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 339) begin : MEM_DATA_339
    assign mem_data_i = {mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115,
mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 340) begin : MEM_DATA_340
    assign mem_data_i = {mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116,
mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 341) begin : MEM_DATA_341
    assign mem_data_i = {mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117,
mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 342) begin : MEM_DATA_342
    assign mem_data_i = {mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118,
mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 343) begin : MEM_DATA_343
    assign mem_data_i = {mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119,
mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 344) begin : MEM_DATA_344
    assign mem_data_i = {mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120,
mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 345) begin : MEM_DATA_345
    assign mem_data_i = {mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121,
mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 346) begin : MEM_DATA_346
    assign mem_data_i = {mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122,
mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 347) begin : MEM_DATA_347
    assign mem_data_i = {mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123,
mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 348) begin : MEM_DATA_348
    assign mem_data_i = {mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124,
mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 349) begin : MEM_DATA_349
    assign mem_data_i = {mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125,
mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 350) begin : MEM_DATA_350
    assign mem_data_i = {mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126,
mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 351) begin : MEM_DATA_351
    assign mem_data_i = {mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127,
mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 352) begin : MEM_DATA_352
    assign mem_data_i = {mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128,
mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 353) begin : MEM_DATA_353
    assign mem_data_i = {mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129,
mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 354) begin : MEM_DATA_354
    assign mem_data_i = {mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130,
mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 355) begin : MEM_DATA_355
    assign mem_data_i = {mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131,
mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 356) begin : MEM_DATA_356
    assign mem_data_i = {mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132,
mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 357) begin : MEM_DATA_357
    assign mem_data_i = {mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133,
mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 358) begin : MEM_DATA_358
    assign mem_data_i = {mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134,
mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 359) begin : MEM_DATA_359
    assign mem_data_i = {mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135,
mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 360) begin : MEM_DATA_360
    assign mem_data_i = {mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136,
mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 361) begin : MEM_DATA_361
    assign mem_data_i = {mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137,
mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 362) begin : MEM_DATA_362
    assign mem_data_i = {mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138,
mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 363) begin : MEM_DATA_363
    assign mem_data_i = {mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139,
mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 364) begin : MEM_DATA_364
    assign mem_data_i = {mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140,
mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 365) begin : MEM_DATA_365
    assign mem_data_i = {mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141,
mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 366) begin : MEM_DATA_366
    assign mem_data_i = {mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142,
mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 367) begin : MEM_DATA_367
    assign mem_data_i = {mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143,
mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 368) begin : MEM_DATA_368
    assign mem_data_i = {mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144,
mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 369) begin : MEM_DATA_369
    assign mem_data_i = {mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145,
mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 370) begin : MEM_DATA_370
    assign mem_data_i = {mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146,
mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 371) begin : MEM_DATA_371
    assign mem_data_i = {mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147,
mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 372) begin : MEM_DATA_372
    assign mem_data_i = {mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148,
mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 373) begin : MEM_DATA_373
    assign mem_data_i = {mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149,
mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 374) begin : MEM_DATA_374
    assign mem_data_i = {mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150,
mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 375) begin : MEM_DATA_375
    assign mem_data_i = {mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151,
mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 376) begin : MEM_DATA_376
    assign mem_data_i = {mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152,
mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 377) begin : MEM_DATA_377
    assign mem_data_i = {mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153,
mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 378) begin : MEM_DATA_378
    assign mem_data_i = {mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154,
mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 379) begin : MEM_DATA_379
    assign mem_data_i = {mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155,
mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 380) begin : MEM_DATA_380
    assign mem_data_i = {mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156,
mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 381) begin : MEM_DATA_381
    assign mem_data_i = {mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157,
mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 382) begin : MEM_DATA_382
    assign mem_data_i = {mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158,
mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 383) begin : MEM_DATA_383
    assign mem_data_i = {mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159,
mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 384) begin : MEM_DATA_384
    assign mem_data_i = {mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160,
mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 385) begin : MEM_DATA_385
    assign mem_data_i = {mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161,
mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 386) begin : MEM_DATA_386
    assign mem_data_i = {mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162,
mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 387) begin : MEM_DATA_387
    assign mem_data_i = {mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163,
mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 388) begin : MEM_DATA_388
    assign mem_data_i = {mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164,
mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 389) begin : MEM_DATA_389
    assign mem_data_i = {mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165,
mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 390) begin : MEM_DATA_390
    assign mem_data_i = {mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166,
mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 391) begin : MEM_DATA_391
    assign mem_data_i = {mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167,
mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 392) begin : MEM_DATA_392
    assign mem_data_i = {mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168,
mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 393) begin : MEM_DATA_393
    assign mem_data_i = {mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169,
mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 394) begin : MEM_DATA_394
    assign mem_data_i = {mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170,
mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 395) begin : MEM_DATA_395
    assign mem_data_i = {mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171,
mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 396) begin : MEM_DATA_396
    assign mem_data_i = {mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172,
mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 397) begin : MEM_DATA_397
    assign mem_data_i = {mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173,
mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 398) begin : MEM_DATA_398
    assign mem_data_i = {mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174,
mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 399) begin : MEM_DATA_399
    assign mem_data_i = {mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175,
mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 400) begin : MEM_DATA_400
    assign mem_data_i = {mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176,
mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 401) begin : MEM_DATA_401
    assign mem_data_i = {mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177,
mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 402) begin : MEM_DATA_402
    assign mem_data_i = {mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178,
mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 403) begin : MEM_DATA_403
    assign mem_data_i = {mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179,
mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 404) begin : MEM_DATA_404
    assign mem_data_i = {mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180,
mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 405) begin : MEM_DATA_405
    assign mem_data_i = {mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181,
mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 406) begin : MEM_DATA_406
    assign mem_data_i = {mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182,
mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 407) begin : MEM_DATA_407
    assign mem_data_i = {mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183,
mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 408) begin : MEM_DATA_408
    assign mem_data_i = {mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184,
mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 409) begin : MEM_DATA_409
    assign mem_data_i = {mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185,
mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 410) begin : MEM_DATA_410
    assign mem_data_i = {mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186,
mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 411) begin : MEM_DATA_411
    assign mem_data_i = {mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187,
mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 412) begin : MEM_DATA_412
    assign mem_data_i = {mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188,
mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 413) begin : MEM_DATA_413
    assign mem_data_i = {mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189,
mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 414) begin : MEM_DATA_414
    assign mem_data_i = {mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190,
mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 415) begin : MEM_DATA_415
    assign mem_data_i = {mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191,
mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 416) begin : MEM_DATA_416
    assign mem_data_i = {mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192,
mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 417) begin : MEM_DATA_417
    assign mem_data_i = {mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193,
mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 418) begin : MEM_DATA_418
    assign mem_data_i = {mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194,
mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 419) begin : MEM_DATA_419
    assign mem_data_i = {mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195,
mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 420) begin : MEM_DATA_420
    assign mem_data_i = {mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196,
mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 421) begin : MEM_DATA_421
    assign mem_data_i = {mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197,
mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 422) begin : MEM_DATA_422
    assign mem_data_i = {mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198,
mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 423) begin : MEM_DATA_423
    assign mem_data_i = {mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199,
mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 424) begin : MEM_DATA_424
    assign mem_data_i = {mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200,
mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 425) begin : MEM_DATA_425
    assign mem_data_i = {mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201,
mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 426) begin : MEM_DATA_426
    assign mem_data_i = {mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202,
mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 427) begin : MEM_DATA_427
    assign mem_data_i = {mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203,
mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 428) begin : MEM_DATA_428
    assign mem_data_i = {mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204,
mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 429) begin : MEM_DATA_429
    assign mem_data_i = {mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205,
mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 430) begin : MEM_DATA_430
    assign mem_data_i = {mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206,
mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 431) begin : MEM_DATA_431
    assign mem_data_i = {mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207,
mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 432) begin : MEM_DATA_432
    assign mem_data_i = {mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208,
mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 433) begin : MEM_DATA_433
    assign mem_data_i = {mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209,
mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 434) begin : MEM_DATA_434
    assign mem_data_i = {mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210,
mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 435) begin : MEM_DATA_435
    assign mem_data_i = {mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211,
mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 436) begin : MEM_DATA_436
    assign mem_data_i = {mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212,
mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 437) begin : MEM_DATA_437
    assign mem_data_i = {mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213,
mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 438) begin : MEM_DATA_438
    assign mem_data_i = {mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214,
mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 439) begin : MEM_DATA_439
    assign mem_data_i = {mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215,
mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 440) begin : MEM_DATA_440
    assign mem_data_i = {mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216,
mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 441) begin : MEM_DATA_441
    assign mem_data_i = {mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217,
mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 442) begin : MEM_DATA_442
    assign mem_data_i = {mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218,
mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 443) begin : MEM_DATA_443
    assign mem_data_i = {mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219,
mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 444) begin : MEM_DATA_444
    assign mem_data_i = {mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220,
mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 445) begin : MEM_DATA_445
    assign mem_data_i = {mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221,
mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 446) begin : MEM_DATA_446
    assign mem_data_i = {mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222,
mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 447) begin : MEM_DATA_447
    assign mem_data_i = {mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223,
mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 448) begin : MEM_DATA_448
    assign mem_data_i = {mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224,
mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 449) begin : MEM_DATA_449
    assign mem_data_i = {mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225,
mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 450) begin : MEM_DATA_450
    assign mem_data_i = {mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226,
mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 451) begin : MEM_DATA_451
    assign mem_data_i = {mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227,
mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 452) begin : MEM_DATA_452
    assign mem_data_i = {mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228,
mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 453) begin : MEM_DATA_453
    assign mem_data_i = {mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229,
mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 454) begin : MEM_DATA_454
    assign mem_data_i = {mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230,
mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 455) begin : MEM_DATA_455
    assign mem_data_i = {mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231,
mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 456) begin : MEM_DATA_456
    assign mem_data_i = {mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232,
mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 457) begin : MEM_DATA_457
    assign mem_data_i = {mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233,
mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 458) begin : MEM_DATA_458
    assign mem_data_i = {mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234,
mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1,
mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 459) begin : MEM_DATA_459
    assign mem_data_i = {mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235,
mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2,
mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 460) begin : MEM_DATA_460
    assign mem_data_i = {mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236,
mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3,
mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 461) begin : MEM_DATA_461
    assign mem_data_i = {mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237,
mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4,
mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 462) begin : MEM_DATA_462
    assign mem_data_i = {mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238,
mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6,
mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 463) begin : MEM_DATA_463
    assign mem_data_i = {mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239,
mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7,
mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 464) begin : MEM_DATA_464
    assign mem_data_i = {mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240,
mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8,
mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 465) begin : MEM_DATA_465
    assign mem_data_i = {mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241,
mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9,
mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 466) begin : MEM_DATA_466
    assign mem_data_i = {mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242,
mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10,
mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 467) begin : MEM_DATA_467
    assign mem_data_i = {mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243,
mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11,
mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 468) begin : MEM_DATA_468
    assign mem_data_i = {mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244,
mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12,
mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 469) begin : MEM_DATA_469
    assign mem_data_i = {mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245,
mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13,
mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 470) begin : MEM_DATA_470
    assign mem_data_i = {mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246,
mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14,
mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 471) begin : MEM_DATA_471
    assign mem_data_i = {mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247,
mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15,
mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 472) begin : MEM_DATA_472
    assign mem_data_i = {mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248,
mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16,
mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 473) begin : MEM_DATA_473
    assign mem_data_i = {mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249,
mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17,
mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 474) begin : MEM_DATA_474
    assign mem_data_i = {mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250,
mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18,
mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 475) begin : MEM_DATA_475
    assign mem_data_i = {mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251,
mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19,
mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 476) begin : MEM_DATA_476
    assign mem_data_i = {mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252,
mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20,
mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 477) begin : MEM_DATA_477
    assign mem_data_i = {mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253,
mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22,
mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 478) begin : MEM_DATA_478
    assign mem_data_i = {mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254,
mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23,
mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 479) begin : MEM_DATA_479
    assign mem_data_i = {mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255,
mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24,
mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 480) begin : MEM_DATA_480
    assign mem_data_i = {mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256,
mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25,
mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 481) begin : MEM_DATA_481
    assign mem_data_i = {mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257,
mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26,
mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 482) begin : MEM_DATA_482
    assign mem_data_i = {mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258,
mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27,
mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 483) begin : MEM_DATA_483
    assign mem_data_i = {mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259,
mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28,
mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 484) begin : MEM_DATA_484
    assign mem_data_i = {mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260,
mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29,
mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 485) begin : MEM_DATA_485
    assign mem_data_i = {mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261,
mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30,
mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 486) begin : MEM_DATA_486
    assign mem_data_i = {mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262,
mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31,
mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 487) begin : MEM_DATA_487
    assign mem_data_i = {mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263,
mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32,
mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 488) begin : MEM_DATA_488
    assign mem_data_i = {mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264,
mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33,
mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 489) begin : MEM_DATA_489
    assign mem_data_i = {mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265,
mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34,
mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 490) begin : MEM_DATA_490
    assign mem_data_i = {mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266,
mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35,
mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 491) begin : MEM_DATA_491
    assign mem_data_i = {mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267,
mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36,
mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 492) begin : MEM_DATA_492
    assign mem_data_i = {mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268,
mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37,
mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 493) begin : MEM_DATA_493
    assign mem_data_i = {mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269,
mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38,
mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 494) begin : MEM_DATA_494
    assign mem_data_i = {mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270,
mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39,
mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 495) begin : MEM_DATA_495
    assign mem_data_i = {mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271,
mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40,
mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 496) begin : MEM_DATA_496
    assign mem_data_i = {mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272,
mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42,
mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 497) begin : MEM_DATA_497
    assign mem_data_i = {mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273,
mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43,
mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 498) begin : MEM_DATA_498
    assign mem_data_i = {mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274,
mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44,
mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 499) begin : MEM_DATA_499
    assign mem_data_i = {mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275,
mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45,
mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 500) begin : MEM_DATA_500
    assign mem_data_i = {mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276,
mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46,
mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 501) begin : MEM_DATA_501
    assign mem_data_i = {mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277,
mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47,
mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 502) begin : MEM_DATA_502
    assign mem_data_i = {mem_shift_probe501, mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278,
mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48,
mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 503) begin : MEM_DATA_503
    assign mem_data_i = {mem_shift_probe502, mem_shift_probe501, mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279,
mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49,
mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 504) begin : MEM_DATA_504
    assign mem_data_i = {mem_shift_probe503, mem_shift_probe502, mem_shift_probe501, mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280,
mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50,
mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 505) begin : MEM_DATA_505
    assign mem_data_i = {mem_shift_probe504, mem_shift_probe503, mem_shift_probe502, mem_shift_probe501, mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281,
mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51,
mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 506) begin : MEM_DATA_506
    assign mem_data_i = {mem_shift_probe505, mem_shift_probe504, mem_shift_probe503, mem_shift_probe502, mem_shift_probe501, mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282,
mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52,
mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 507) begin : MEM_DATA_507
    assign mem_data_i = {mem_shift_probe506, mem_shift_probe505, mem_shift_probe504, mem_shift_probe503, mem_shift_probe502, mem_shift_probe501, mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283,
mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53,
mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 508) begin : MEM_DATA_508
    assign mem_data_i = {mem_shift_probe507, mem_shift_probe506, mem_shift_probe505, mem_shift_probe504, mem_shift_probe503, mem_shift_probe502, mem_shift_probe501, mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284,
mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54,
mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 509) begin : MEM_DATA_509
    assign mem_data_i = {mem_shift_probe508, mem_shift_probe507, mem_shift_probe506, mem_shift_probe505, mem_shift_probe504, mem_shift_probe503, mem_shift_probe502, mem_shift_probe501, mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286, mem_shift_probe285,
mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56, mem_shift_probe55,
mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 510) begin : MEM_DATA_510
    assign mem_data_i = {mem_shift_probe509, mem_shift_probe508, mem_shift_probe507, mem_shift_probe506, mem_shift_probe505, mem_shift_probe504, mem_shift_probe503, mem_shift_probe502, mem_shift_probe501, mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287, mem_shift_probe286,
mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57, mem_shift_probe56,
mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 511) begin : MEM_DATA_511
    assign mem_data_i = {mem_shift_probe510, mem_shift_probe509, mem_shift_probe508, mem_shift_probe507, mem_shift_probe506, mem_shift_probe505, mem_shift_probe504, mem_shift_probe503, mem_shift_probe502, mem_shift_probe501, mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288, mem_shift_probe287,
mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58, mem_shift_probe57,
mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end 
 if (C_NUM_PROBES == 512) begin : MEM_DATA_512
    assign mem_data_i = {mem_shift_probe511, mem_shift_probe510, mem_shift_probe509, mem_shift_probe508, mem_shift_probe507, mem_shift_probe506, mem_shift_probe505, mem_shift_probe504, mem_shift_probe503, mem_shift_probe502, mem_shift_probe501, mem_shift_probe500, mem_shift_probe499, mem_shift_probe498, mem_shift_probe497, mem_shift_probe496, mem_shift_probe495, mem_shift_probe494, mem_shift_probe493, mem_shift_probe492, mem_shift_probe491, mem_shift_probe490, mem_shift_probe489, mem_shift_probe488, mem_shift_probe487, mem_shift_probe486, mem_shift_probe485, mem_shift_probe484, mem_shift_probe483, mem_shift_probe482, mem_shift_probe481, mem_shift_probe480, mem_shift_probe479, mem_shift_probe478, mem_shift_probe477, mem_shift_probe476, mem_shift_probe475, mem_shift_probe474, mem_shift_probe473, mem_shift_probe472, mem_shift_probe471, mem_shift_probe470, mem_shift_probe469, mem_shift_probe468, mem_shift_probe467, mem_shift_probe466, mem_shift_probe465, mem_shift_probe464, mem_shift_probe463, mem_shift_probe462, mem_shift_probe461, mem_shift_probe460, mem_shift_probe459, mem_shift_probe458, mem_shift_probe457, mem_shift_probe456, mem_shift_probe455, mem_shift_probe454, mem_shift_probe453, mem_shift_probe452, mem_shift_probe451, mem_shift_probe450, mem_shift_probe449, mem_shift_probe448, mem_shift_probe447, mem_shift_probe446, mem_shift_probe445, mem_shift_probe444, mem_shift_probe443, mem_shift_probe442, mem_shift_probe441, mem_shift_probe440, mem_shift_probe439, mem_shift_probe438, mem_shift_probe437, mem_shift_probe436, mem_shift_probe435, mem_shift_probe434, mem_shift_probe433, mem_shift_probe432, mem_shift_probe431, mem_shift_probe430, mem_shift_probe429, mem_shift_probe428, mem_shift_probe427, mem_shift_probe426, mem_shift_probe425, mem_shift_probe424, mem_shift_probe423, mem_shift_probe422, mem_shift_probe421, mem_shift_probe420, mem_shift_probe419, mem_shift_probe418, mem_shift_probe417, mem_shift_probe416, mem_shift_probe415, mem_shift_probe414, mem_shift_probe413, mem_shift_probe412, mem_shift_probe411, mem_shift_probe410, mem_shift_probe409, mem_shift_probe408, mem_shift_probe407, mem_shift_probe406, mem_shift_probe405, mem_shift_probe404, mem_shift_probe403, mem_shift_probe402, mem_shift_probe401, mem_shift_probe400, mem_shift_probe399, mem_shift_probe398, mem_shift_probe397, mem_shift_probe396, mem_shift_probe395, mem_shift_probe394, mem_shift_probe393, mem_shift_probe392, mem_shift_probe391, mem_shift_probe390, mem_shift_probe389, mem_shift_probe388, mem_shift_probe387, mem_shift_probe386, mem_shift_probe385, mem_shift_probe384, mem_shift_probe383, mem_shift_probe382, mem_shift_probe381, mem_shift_probe380, mem_shift_probe379, mem_shift_probe378, mem_shift_probe377, mem_shift_probe376, mem_shift_probe375, mem_shift_probe374, mem_shift_probe373, mem_shift_probe372, mem_shift_probe371, mem_shift_probe370, mem_shift_probe369, mem_shift_probe368, mem_shift_probe367, mem_shift_probe366, mem_shift_probe365, mem_shift_probe364, mem_shift_probe363, mem_shift_probe362, mem_shift_probe361, mem_shift_probe360, mem_shift_probe359, mem_shift_probe358, mem_shift_probe357, mem_shift_probe356, mem_shift_probe355, mem_shift_probe354, mem_shift_probe353, mem_shift_probe352, mem_shift_probe351, mem_shift_probe350, mem_shift_probe349, mem_shift_probe348, mem_shift_probe347, mem_shift_probe346, mem_shift_probe345, mem_shift_probe344, mem_shift_probe343, mem_shift_probe342, mem_shift_probe341, mem_shift_probe340, mem_shift_probe339, mem_shift_probe338, mem_shift_probe337, mem_shift_probe336, mem_shift_probe335, mem_shift_probe334, mem_shift_probe333, mem_shift_probe332, mem_shift_probe331, mem_shift_probe330, mem_shift_probe329, mem_shift_probe328, mem_shift_probe327, mem_shift_probe326, mem_shift_probe325, mem_shift_probe324, mem_shift_probe323, mem_shift_probe322, mem_shift_probe321, mem_shift_probe320, mem_shift_probe319, mem_shift_probe318, mem_shift_probe317, mem_shift_probe316, mem_shift_probe315, mem_shift_probe314, mem_shift_probe313, mem_shift_probe312, mem_shift_probe311, mem_shift_probe310, mem_shift_probe309, mem_shift_probe308, mem_shift_probe307, mem_shift_probe306, mem_shift_probe305, mem_shift_probe304, mem_shift_probe303, mem_shift_probe302, mem_shift_probe301, mem_shift_probe300, mem_shift_probe299, mem_shift_probe298, mem_shift_probe297, mem_shift_probe296, mem_shift_probe295, mem_shift_probe294, mem_shift_probe293, mem_shift_probe292, mem_shift_probe291, mem_shift_probe290, mem_shift_probe289, mem_shift_probe288,
mem_shift_probe287, mem_shift_probe286, mem_shift_probe285, mem_shift_probe284, mem_shift_probe283, mem_shift_probe282, mem_shift_probe281, mem_shift_probe280, mem_shift_probe279, mem_shift_probe278, mem_shift_probe277, mem_shift_probe276, mem_shift_probe275, mem_shift_probe274, mem_shift_probe273, mem_shift_probe272, mem_shift_probe271, mem_shift_probe270, mem_shift_probe269, mem_shift_probe268, mem_shift_probe267, mem_shift_probe266, mem_shift_probe265, mem_shift_probe264, mem_shift_probe263, mem_shift_probe262, mem_shift_probe261, mem_shift_probe260, mem_shift_probe259, mem_shift_probe258, mem_shift_probe257, mem_shift_probe256, mem_shift_probe255, mem_shift_probe254, mem_shift_probe253, mem_shift_probe252, mem_shift_probe251, mem_shift_probe250, mem_shift_probe249, mem_shift_probe248, mem_shift_probe247, mem_shift_probe246, mem_shift_probe245, mem_shift_probe244, mem_shift_probe243, mem_shift_probe242, mem_shift_probe241, mem_shift_probe240, mem_shift_probe239, mem_shift_probe238, mem_shift_probe237, mem_shift_probe236, mem_shift_probe235, mem_shift_probe234, mem_shift_probe233, mem_shift_probe232, mem_shift_probe231, mem_shift_probe230, mem_shift_probe229, mem_shift_probe228, mem_shift_probe227, mem_shift_probe226, mem_shift_probe225, mem_shift_probe224, mem_shift_probe223, mem_shift_probe222, mem_shift_probe221, mem_shift_probe220, mem_shift_probe219, mem_shift_probe218, mem_shift_probe217, mem_shift_probe216, mem_shift_probe215, mem_shift_probe214, mem_shift_probe213, mem_shift_probe212, mem_shift_probe211, mem_shift_probe210, mem_shift_probe209, mem_shift_probe208, mem_shift_probe207, mem_shift_probe206, mem_shift_probe205, mem_shift_probe204, mem_shift_probe203, mem_shift_probe202, mem_shift_probe201, mem_shift_probe200, mem_shift_probe199, mem_shift_probe198, mem_shift_probe197, mem_shift_probe196, mem_shift_probe195, mem_shift_probe194, mem_shift_probe193, mem_shift_probe192, mem_shift_probe191, mem_shift_probe190, mem_shift_probe189, mem_shift_probe188, mem_shift_probe187, mem_shift_probe186, mem_shift_probe185, mem_shift_probe184, mem_shift_probe183, mem_shift_probe182, mem_shift_probe181, mem_shift_probe180, mem_shift_probe179, mem_shift_probe178, mem_shift_probe177, mem_shift_probe176, mem_shift_probe175, mem_shift_probe174, mem_shift_probe173, mem_shift_probe172, mem_shift_probe171, mem_shift_probe170, mem_shift_probe169, mem_shift_probe168, mem_shift_probe167, mem_shift_probe166, mem_shift_probe165, mem_shift_probe164, mem_shift_probe163, mem_shift_probe162, mem_shift_probe161, mem_shift_probe160, mem_shift_probe159, mem_shift_probe158, mem_shift_probe157, mem_shift_probe156, mem_shift_probe155, mem_shift_probe154, mem_shift_probe153, mem_shift_probe152, mem_shift_probe151, mem_shift_probe150, mem_shift_probe149, mem_shift_probe148, mem_shift_probe147, mem_shift_probe146, mem_shift_probe145, mem_shift_probe144, mem_shift_probe143, mem_shift_probe142, mem_shift_probe141, mem_shift_probe140, mem_shift_probe139, mem_shift_probe138, mem_shift_probe137, mem_shift_probe136, mem_shift_probe135, mem_shift_probe134, mem_shift_probe133, mem_shift_probe132, mem_shift_probe131, mem_shift_probe130, mem_shift_probe129, mem_shift_probe128, mem_shift_probe127, mem_shift_probe126, mem_shift_probe125, mem_shift_probe124, mem_shift_probe123, mem_shift_probe122, mem_shift_probe121, mem_shift_probe120, mem_shift_probe119, mem_shift_probe118, mem_shift_probe117, mem_shift_probe116, mem_shift_probe115, mem_shift_probe114, mem_shift_probe113, mem_shift_probe112, mem_shift_probe111, mem_shift_probe110, mem_shift_probe109, mem_shift_probe108, mem_shift_probe107, mem_shift_probe106, mem_shift_probe105, mem_shift_probe104, mem_shift_probe103, mem_shift_probe102, mem_shift_probe101, mem_shift_probe100, mem_shift_probe99, mem_shift_probe98, mem_shift_probe97, mem_shift_probe96, mem_shift_probe95, mem_shift_probe94, mem_shift_probe93, mem_shift_probe92, mem_shift_probe91, mem_shift_probe90, mem_shift_probe89, mem_shift_probe88, mem_shift_probe87, mem_shift_probe86, mem_shift_probe85, mem_shift_probe84, mem_shift_probe83, mem_shift_probe82, mem_shift_probe81, mem_shift_probe80, mem_shift_probe79, mem_shift_probe78, mem_shift_probe77, mem_shift_probe76, mem_shift_probe75, mem_shift_probe74, mem_shift_probe73, mem_shift_probe72, mem_shift_probe71, mem_shift_probe70, mem_shift_probe69, mem_shift_probe68, mem_shift_probe67, mem_shift_probe66, mem_shift_probe65, mem_shift_probe64, mem_shift_probe63, mem_shift_probe62, mem_shift_probe61, mem_shift_probe60, mem_shift_probe59, mem_shift_probe58,
mem_shift_probe57, mem_shift_probe56, mem_shift_probe55, mem_shift_probe54, mem_shift_probe53, mem_shift_probe52, mem_shift_probe51, mem_shift_probe50, mem_shift_probe49, mem_shift_probe48, mem_shift_probe47, mem_shift_probe46, mem_shift_probe45, mem_shift_probe44, mem_shift_probe43, mem_shift_probe42, mem_shift_probe41, mem_shift_probe40, mem_shift_probe39, mem_shift_probe38, mem_shift_probe37, mem_shift_probe36, mem_shift_probe35, mem_shift_probe34, mem_shift_probe33, mem_shift_probe32, mem_shift_probe31, mem_shift_probe30, mem_shift_probe29, mem_shift_probe28, mem_shift_probe27, mem_shift_probe26, mem_shift_probe25, mem_shift_probe24, mem_shift_probe23, mem_shift_probe22, mem_shift_probe21, mem_shift_probe20, mem_shift_probe19, mem_shift_probe18, mem_shift_probe17, mem_shift_probe16, mem_shift_probe15, mem_shift_probe14, mem_shift_probe13, mem_shift_probe12, mem_shift_probe11, mem_shift_probe10, mem_shift_probe9, mem_shift_probe8, mem_shift_probe7, mem_shift_probe6, mem_shift_probe5, mem_shift_probe4, mem_shift_probe3, mem_shift_probe2, mem_shift_probe1, mem_shift_probe0};
 end
endgenerate

