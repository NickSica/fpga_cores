`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16448)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5IKuj8mgBxS3/HebTMVlzJ1vjfj1ijx3SLL65K/xYdCiFAUCidOrmzed
2+4h/MahfwPHHMNoNd2K5w/ntf59RBL6Ao3gKoB3wvgtdZE6eauMLuqs/POeP0XaMXm90lnihFxX
ounqzySjiVjdYTs5sIXKx3bY1Zx/5qZDuswepE+BPgdoZrCFCaTd9UBfp5yMzdJ1QJI0qA7+goYQ
PJekp6jv4/wONqgXdrWuYSrnV5mLRxm+teMEHYPLGp8Oh65SMJN8RmQt/LNPv/bYCceGsflioHHT
pg8i+y2PqK14T6h3HOLEuJqqoq57stHvJ1eeQkKq6X5l60zoD3H8/BkJcUZKlZb3HBM8Fjx0XMXS
T0YFne1deQjwG+GC7n1pgYUrYmQ97cVlWrE5Gs1vx5IgsQtwzdjf2xbK61vbejCvIPtixIaKrv65
rwZ9yWbIe+yABskr3VCz0iUbAh0Zdh5pmoIQZDoahEOeeW/LNlFQbnru2V41YLEBvCEYOraU4vZm
pObIF3lidxlfWriCeKit8w+RpyTGAGgVlybwU3AkYP0z0B1IKJks/2Jj6rRP7xps7iAk56B+JWQx
G5AHJWwN+lgCkt6D5kLmLzfomaOhiI9y+5jyo3f6m7gtXnd9UD0aQF2yQ8YwX0XOchvGkmVGSm54
3/i4YKbOSWdMVwuB/q1+4WKMd22gylq6B7mCOxU1filYQWmB+EpaX5YwOkJ6c9srQjLC02RLhcqN
NhmkWAXQBaHITrwI+pZ9dx4Wu/0ceiw6muqaX299OO7jQcfWD2Tb40PBiXZfBu4qoz0QJp0ThnVr
2COQ4bSJmyjH6kcHbM+EO0Ix/XF8S1NAKfaCuGwlQhzXiyjiWnDvbKjTdN0EGPUWIWfL3EoVnU+W
i0TBhxUgwzJ5TkfUZb9TuAQCnUz83vqmTimM6v48TgtDoUVOCjK9XvLbmqpGcLa7wsGamd1JdHnW
SC57HDdYebcO3Rjy66uYEWvhXaF+/V8B8FS5P7ICxku08xd4MVtY9+NgGXJZzp9FP+RW0Oc96qAa
MDfcPE9ovqdI7hsvyWnhVP3Xb2u6R8+oc8CzYuoJfwyz74ADvg4torFTdc7zN3TqdbRjETBCxZTI
bbJx2f54QRwLDxJ/IgPkPBI6bk0AODkbgidba5LEM3mRopjrBx9o6WT5tam3fx/5sdEwEQHEq+kK
3xAhDcrcf2DufgWs/PacSn+1zYnhaoqADVzXkg3xLKAM4/iFen5BCYZvDHO5oJsxLHSuy/5nZ4s9
FeqIL4PkwfhC4mWcUzkE4sXQZNvgMDpGUR4J4S1F02+MIuou1ysQfCrYOVfqtlxfrCZdclRurmKz
YCEPDW11oNOBYSTwSVU5VbBaxdYUE6M9Ipy3vXZGUpGeEj/15RbtNVDb0W0UdHvX3+7pOSP/GHX3
elbuhfP8ZtCh1WT3D6N6g543pUNc34aX0tlF2IlHPFUxAN9CYwZx5IFuSSlcJZNULNzW7qChL+sy
Lyj+DSV4Jk2ck45m/LQTAR0ayfoLr+lsO113KGH3qi3euWQcA5axPcKqoCExzkO81q2vlMfjPnYQ
WUr2eGdxn91HB9GH5edgyA89wAzVBmlqamxnQJTNvvA+rf/hF9MPY5YaNvnlQr6HsUYO47vaRdsD
MzYF3vM9w5UowLt/6rKgB5lTvAQulfErZKt2hpOQyOOOVQIcK2XdbQjKBImAlI0hRuqx3yontzVK
PGrD5tSH0nsIc0wRAqIFce4LJsPbEFLHnAISWPYTSVCA2rDpvgaObBZPoK0eL5pBQmHOL6DcacGq
TxcN7mZL1XvD1KWF4f7pNAiZYrlWN91vWpbJSwKp9kzx2OiCmqSRPyV5B7iYal6RPOjMkGrykzOb
l81eNhL7s4pWOC8hD86bbU39YcUJwWtyH+cdZWztU+aZCGbC0Qpslaxt0eC+t6Ic2owmOjofXNjk
bB/oZozY+/Cb2KiAjGXE9qFuPIVm+Ab894ZqB4r32SjjCkluKSBp42w4VGaSEQCxwl5ktqsUnOEl
KYwiV3VTxUId/MN45rvC01Po5XiTi/Ael+B40e9OzvkdBfsLh3FCEmTK0pSA8DbO2QqrXVP/8GKF
IAeXOuVLoFzL8Ub7GJ4dFNIQoGjCFFA/Wd5PR1Gy0Rc/inahVNwDUAORYd4RhXvmhncgdchvsfUf
lsvJNrbJTYryu2RhRBkd9UFxtJ55VTqKlnU8TKI7FxZTC0EF60s5jCfbdcauGvGmnBbnnfGdQSM1
yBkfJycYVYlaubLZH/iUM9Oqck7qA0r937SIMIAApLaq7NAv6yb2GKORIOxefJQ5eqeVrhhlUOWK
MoVIOZ04uLZhD+Et6wEIpTEsgbEy5iC+Gz8eAnUk9s2r8CKX185VRNku42ebyp0Qxc1FXqVfZ2z+
4pvcN5Fn4t2PLVITI7XmUfnXMLTlCEX4oR/Uk/FehcpNGTvBdXnPkw/YvG1UdD+/bA3SDEiQIa6l
ooqv9VawKCvYEDDymxmFslnIgU9/zVZnzb8AONkf5NWNbEICFK1yueO7fCCgqI1ycVFMzJNLtPaQ
un9Ew54xdGhR6tjTD9kwzo7TXhB0vQLo3PVVAhD8R/wqWYlYVLYFX41YDrsRbmqL+1W95bRdTYed
NFodogDRraR8pKXuNpaGFKxL/BGWk6mWdsNLeLda7JlZ0IrQcWS+HFgga7K7GYs7QG5CmQ9uEIwp
z9qEIhxXv/tHN4U1KDyrFW82u6pvYpPvctmuAFKlLYDXgdcQxETIgmwJDFt11B2bCtzzwATv11rI
Ro5d95xI3YHqZm3YSND2Uow8+qh1efO7/oor1FKnEHSNrjvIuTcrlvnDY/pgXbx5Kk/dQbojmQTW
0ck364ZbpEYeHQF5tzLSiiNHlcBVuoiS6u0JelF0fBbQULyC0jr7THgMIWO64kjdIK9+e4U2Dr53
of/5qtNfBcXx5IyPKWArS4dfeRGZvOLFCzGItYpPrWA6eM7S9cDIjZ6498qhZzeVvlE2/bjq/ERk
p2Phai+9CILRp/ftTA2CUi42ZhDBv5+HsPrK/B8UOKxBO0h5Q0GPIPtTTjPnGDm/8IfQlvaiR0zv
fXuih2y8TuGsjUMgKuGCtPwIjTGzRrw3vbUSNeWZMHnraXqGcBcmh1u7GwONN7gCfXaZ2gO95lA3
vWYBfNDBW7xzi1Iyy7ikxNpzcxlAKlnhXCmaye12CQ3xbTwXmKW3SxWu9J8RDFnAOtrRUVQBr6lB
z0fkkNe6FXtLKHcIcoMoTdjlqwH3P+A06zL1ZYfhw0tYmNv4cZAdSfRy2pxij9GishmfufHxExKv
DJ6F2bUr55qHQr0w2OjaXOkt1Cvg+K8/55SLfuNVOq9WoEIYBBCqtcWGfdCLvLRZ/y9BIOcuRUeL
0eiX9GUz/wcIGdGxmKeGGKwyZUkVceXDp6bNo/Y67KmiA4xgQz3fp+0S7uaazr09Cd0cQGMXofGj
kTHkrt8wGnyjtUANZeVn5O1cqra1F1sgupPT7nn8J2OfIaZv+q7HHa2dcbSJMsOgZ2BZUb1WNLrq
1ciLDxeZTPMY541aUPVPyx5CDCjzxUb9P6rg0Sml+aMzdHvKFN7EapKgAolv+Xug23Vdh2B2N2PL
O3CCkDMAZrul6klgNWaGWfDJizU6oiRyjx4XeQB/nKCiXNOiKAtrui1FOKwigt8EtyhvBO19p/tZ
EPRdLTY69r8P1KCwMbgyhqG2bjvC3Yrjm4WaF8NaHr1lrTqtFK5ZN0ae8irpoCYnZoaR5iHwvH8M
BekOT5OjgjiOsRlrdbd//f4bC4iv+5VXkQOkOV+YPsfV85V4GyMXcFszOK65OOP98QA+NLts8MGc
l2zHnWYF7VTtDc0YMMyxORzbpuoLbgPuFKXm/Pqo8hrE5CAM43ZsMFTA05YKG6u4ifVj/eC4qYc8
0YfKWnP0S7/nyJEkvwVeXeo7trVLxdKyj/emkmWKVmNSy9VziqBj5WbApwKT6ZCqx9yDz9KX4hsL
XZ/UCY5pK9u5vwfLHfVmEwgFVRNjulJlOU74nfZnMh7nbZal0EcI9VURbuQr2Yltt/azVbcuUhHx
rsyJ0H2quF/glIaX7Ecel8vGcwJDXOVk3xQOS89/YVmser2RRJsOTYpUFuUW4L5ZHK8fA3p0P8Pz
OVtOX10m8mhsG5F4s1G+qacR7ISIWB/udnUrsLrm7A+mU2JgghtafN8F3rz0tf0/HyGqed19esTN
PRdZGV8M/hl9RZc+fpIAJp2e5Nladtlq96/spAo1+X/4yAHu24P9igZS9e8wC0cU8g4dZOnAp+JP
qTBH3TGWK8OL8YtdgMOXHahVJbTBMWjzah7GM7YfxSUtbrKNoNT6U1v3mT+9DO7PPtN9VyDFxV5t
x5THYOotIYMz3F/GA+L/CWbSkFUb6qBzPL5PAFI8i0RRqvs27RIyIDLo2//lro0WJo7WUlts9CMD
iEf3NahfH1d9yaXcLNHJgI2WS6vP/HbHdQVjlkHDd4DBaH+FqiKc7/d4gC1qrMjbZ3x/BNe5L3io
aUF2lIT9a+PE/8ATgrAFINXjVC29EOdr96LhjDOLwRRKpe6ayyrIxu/9G1EN+k1catCg4tKvO5Ze
TaWSqVc3XrnFMm5ghMtoGAOx/L5RS/vpOrv4GJQ9x0A1SGBTjgWNP+9O6OjPItQlxMLr462CE9ht
EWnk1URjj3/WFeJ5X63MBLmRCzoxIpwDXNANkECflBC9A/U0wj8IuNlIZI9vbs/wM5H0sNERYB07
unLRGSFUdH0JtzkGhLxsBbHCfjuZVTpEPSQEBu83AxbMQS124rdhUUYHAfViMt8mh+ZIDUh4m235
IOUhaAe6Srj7uuBj/SK+0NarFdRpCCv7V1cHWQyGP8NH1wFrhbITCICKDt3Q+k9jkCRul3WnvHql
NaLZz57KXN+iLDUqlDeW09LwH5V79NWMVFTXUWvr/LQvZGyAkPwmpQyFDs7uyGezmQW5L8eo3HAF
6Yd0zvt/KCNK0CYaeQ2yMtj407Ghczg1NcS76iKtV6rsifcNH9REu0+cHAHk8qm8M0PLsiAObgAk
NzQiNLOjmKsJ8mNK2WweWPhOLPiDhbbdwN9aX2hF+glXALG0nHH0NNbfxZ6ii1t0WlVe+vaDptf6
EmnC4CpY0T8535AqdZkDdoo+TTraIKsKZFuRY5tscWyQbPakd7VKTxBwnvEsXuEaLp46xddgBa4g
ox9nH2F5Fk3wYpqJynW/mXuylc1SdkYz00MvC1vbmyY6niu9GpJ+3fiavalzHFNsXfEvfaLSjk2T
4KKfYETILHgjjKDQR5kPGEG134coBD1S7N6QIU/mj3guZZDJWpflGrcn3/Kim40d9qlgVMO/qZp7
qW5CqWFieUKPazfDf/MwCPpDzVcQS4hlCx4/pSKOjFdMUcrLzzcqx3qNijxPabCaodDGWOcq9XK6
PV81G5GP/yP2cLt8RI/4X7iDc4KRzTR1l4pJNydd8QE9zo4YTYukbmZs1iz1/jwvRQNriRg92MTH
5UTm+XEq0hAFkCv70FMahmzvvHObkzYPgx44NoS+etbpTUAdUfJuqYTZC8xR1EdlYUU4h4nnfj4+
Ky3eZNYJ+EN1lZ18PGMuM2rperYsDHu7apJSHL1OHSPR4BJEjTEM/VzKStCHwEypkHD+AJ4SiXS4
5sISdtznN7BhcmMknKoZiYrNJLMpDWjEHtEVCQkwajRoUmDCE8wR/k88QGmOO+K/GQcw7QdsHHKm
k2sPVk3f9botZNvTci8tCFQ2JKRnYW9Ys3nOeB0YXMWV9gVPDYlkp5p52WbasSpuLLvnVET2PZag
GsjPMLC6L+QrH/bCCBPM6bZTJrj+uNW29UDeVzs6kbi37fnoIgWcDs9VM4OlLEBxnq4dB9RubMVR
yqVY2nS+hVSWgIejWto0B3LkwwQTAsThVouWExbEnk0LY8bFf+ibw4xcpIvUyXtDt0KWf87oHK+5
6tdjBSfpWIxfXxEjDFgUYVvPLblDyRFUdo1HTripRKPcypjyzR12L7fc4y7rV9VtUt/j4LZHnaWj
OzgkxW7LDllf/4Cbk79T3Yic4e4IV8Z76poJZP+kg32HBtQ2kzLeW7oydssvN2iknetUq4DXVmzf
RbZiBYAm1Cjhufxw0IMOEz4hCBq19/i1aTRBxZvSFkWvStU6R3gc3PCHLFZjtDcNtsP5V8psSOZ0
YouoiXfSXvcNnrfi3FPz2IWulNTvWt6T4rmfIwX22fF7H+0PLn8zfzRTi8iXCXaTgv6j1xXYGP63
ot1p2vrHRUjNgYkpfpcXoDcHtjDYrLJiNdymbe+U0QBsz76PXw7xxQpUgdjJ2BqUSealm9GPf+Il
MKbjzHGbSjsi+4OF2hgeXMBk8CdRRx2hAz83ITrk9liJDwq8aGbhop0Q4To9uOFejx/vhn2SpROJ
m6pJ9zhqhqlRmPtEbCcOT90oVfn7Ltj4EjA/1kuo6jPoUC287iLthj6DtyiGui353H+xpUA1CcaB
N0PZmGmEe1QPeMCgbHPm/dcIH5efmGzvRCBaaOGFXpl7aii7lnkRtt+eQ9A+LUkcji/+L7Fj2psS
dLoqccwgiHDQI+7lxRdcwAVNEEqbnkUFZwpFW3GqS7mAkq8uWKHEBDeagAjRscY0FaXbRwO9jZs8
Ls6yLFtnIBwbVg2DcdtXj0aJTk23hHswqdQw8R0/EU8iLaQ0UHvKlo7nvXv+zQ1Jy4tvPi5rB756
zWL4obAKsOnwgqpPL3V0NXW4v/qHmrcVbVTWYO1wC1xuo7+I6sNnbiTfAWFchIav4LFYJmxANM2G
cgtdpT+4CAtFAO7eifn4LDxBhcDLOh8BukldTIGBQIxmB22P6Qz8AMg4WZnH5ziTjnSDG3WPg4ni
RYW8+xPLTYsyT14YiHaBtLfCcnujEEA8KmDVH4k0Y/H7EKgFz6ND7HWcmD2dV4WLPC0crufR9K6y
5Qs7MwsrntHmA0Bthjt1d9GRwSML2/VYpscAYAZGddRy/JiMojIqDEzGl0YLndMCR0jAzDrEv5mX
l+YJuGfSJBapFwJw94EbgRRzCRtkM2PYTzXl/or/0Dex17x5cbzQ8+RSG9zqwaUxMcTfBPgD4OLC
bcRlpFBiCH+jHtK4fNs5u6ienJ1F2gsCSFTANlZAFuFk5jyPv/MgmiCw6TxSh9KmEE2IQ/BwUk3X
VhBjAnUFecnpcw5yo6Yx5+EF4lQ3BIKdd9/yXYzzAFcGwzo691SjDxkow/XK87MaN67Nh+/2Gs85
+bVdEv/0WIz1k9DwupmLXmHmfTbLnDqRt475x/tFtWaTdlp3h8rcqmPuXjBhYxPsxHVJlYH697dh
cgO/nQ23ojpZiUB3D5cP62LIfTLPuVeERuk/l/GPK8PVE5oik0oH3Pix54gvBfRU2Y4asY2LjBFa
Cf0P0QZcLCFgKZP4mfW1M8HDLvcAOOfEEDm4pAeEskJGodKHLMiAo1Chc94KawAXprVvypY6wBzC
PvhkOkxDP5TWewSQjAiiE2wlHXunb/MJTfVEL02wR9lMX5jfD21LyL9kum85dQK2DJZ3CfknEW89
fXfoOYWBNmzbHZPfVjkjIZwTxlP8BLmjSO02HNkrFCoQPm7VbHOGC1bFKd+91VZhhteqIJupJeWB
cLHgDnvOwv2P8uy33u71EYu4UJ7nfaAYy/A/+J5xVbDPGdOUP28P27tbZ0b/pIgeUZTG/TFMNRnL
WLUhYDISE2kr5jZ+7jVwUC8fenNFiYlQ5OJzx3owJ7s2f+dUUs8FjdPInQZgSuvxxWQGVoIZ7WpZ
0OwYFLyppniFCPJQ4YtlVX2UkxOgmBq2YwVi32Med7dBsk8PJ54d6o01U0Pa6mL/w0NYkDy5EFGp
LEbdHOq8vMSB3J8STfhVD+o/wtO2WBN5HTvTSSUVwUW5X7qTcIgg3ClOjbC5KqGBEHcxQVHxybsN
A4Sr+aDFNRghmCLMR4rt8Ujjd9u49XKrivyoE/qJIZ95iekA4wsg4YusON9OAWJROPze6JnCpC+b
Inlyj8RmsP6LvnMd2PUln2KzvQEbvKicDYOaFRw2H7edt5EgHJ2Wt6iE3ERnUi38UYObcxt6+Pw4
uF4rXou2mJQOoqqPliCMZ5nUmMNcUp75xKZxERLN9yKxtHDlCAPF99dpX2hiMTt/9MTjod16gha7
Y1H5H/VsQdTcVRQkBi5s1wUa3xkCb7JkHCgaxy8qGpb5dWw2n15suPoQ8e0308GgcVmwZlh1abA4
aH8YjZb2iASZgqC8uzNPy3lw2TAO6Br7qlp4WAfuYKRLy9UfVKRj+kRCM3y+RNF2psXuPWhC76od
wrdeXhhfssMX9/HlQkmUVZIvPgd3E/3x02PbX348keZy6xX7bBm1R2/Yi1OzgZuybIU2VAp2YCt9
DV9AXvp7ngCWPcO4a3CORlrmqYAfUbNy+B9nFzlox+KRFfwhYXKa2oOd1GmgvVVxjRIOnyW0bewn
UG6B0K9z3ZGrb6mXznTB387jrAGiHoadme5RhFrDR4ZeNwNcIxspZ0mc/72GCY3szL2S00PaZVym
JoWkofrlMW30SgBZ9IzC5sY7FJ3/u3PHSw+8dUiAxB8bf2C78j0ODTovSuY8NhV/6ohnml3OziF5
Cm2GiQ8ruZ6ur7AubV+oXIjNIbNh4uhP+WwrOJBNac4QTE/mJ9ZX/rYDuqvhcqnG/TF9bOp2aGbw
Seg2xlmF5Y8/gF6ZoRPPZlr1rqAS3uAkLs1sMQaijz8YubxBl8Jjsoo3LKNNufCJrADeBT4HE4VY
h/O1Qy1n3TIm9gv8zGEVI7TPTnJ3NOH2V7nafafdobxjlwHyPtqQhpWgsqzW1cCpLd8nIbBT4Ced
C2W3N+ENpYasGS4noPD2JtY6kRavmg+ujA1TBjLGnSDrj5iG30rr6xQETotXtJwtFT3J4zlMSZFZ
TQbw6CevH/tkso9ebcl7oiQlla0ORv3bV3RH4glYuuwJDhhvvmqyzIhrOyBMCA1jksUWouDKDU4X
8yX9Dk0QAsYjsX/ZF3PX9B+jSIXhpF+fCW7LANAvYmuGqAO4BilQpuX6iM4wWI2ISDWxBMFL35Ka
gaOyVSP+H/vZj/Y5p9vy9/jd5DwwrX7IJXjZ0QtDd453E7UIT6cQO4Jg0W1qOlYeAz3z1TJokTCM
dvzoHgXup1SWgi/lbNp1IP/HzI9BxZHo0SNZ3Djb2vyrtgAjFFr0t/tWX0ukirPUxKEV9Q6dZDWC
mthRIcs/RZ5EE9LSq2ish0gqPop5RudLvuCFzOqwdLRdTtBGoyYaOq8AXriUyiRuwiCTJPaiGzON
6GJ/1bXN7NAMWnXausfTX24wzS8/OXIRdvB0AWo4c6LoPTTJH/4627c40/3QhO/Rsili0/JyDTbM
fr/W6DqdnGvOb5xHtnTifEWRjH/0HWIsDRZ8LAz0GHzsH4I1wu+Tr0aTJVvKjtv+iBS9SzlkF6Fb
bddmWqh0S2+Atj8y5BHhDC4Y6PpFFV/Lo5FDc1i5KVcduQwh7EFxUqy+YjWkl7dhXbvX8jKG9Ydk
Ih1ETarxa3xTfXO6hZb8UVKxHZ2XVUdQOs1ubf/HGpzoZuu0Sfia1E5b2IYDwg1uT+bCbQMwmvgV
AL8fMBC+XQerhBK+MlTrmcyGBuHMYR3oT15M/hn6ParX8agVhGJjfFE8Drj1IEaWhYBoJug1M7lY
Vs0PUdpnJxRQbzDDxi4YA/4FRlr8TrRL4te2+RrdmqXhcgXeF3C397P9zHd2glpp4Z++MuQiBej7
4o+EKvqAAzT4AkV8DbBpCHoy27N/IjwfKXdaxWn87XMSYBPVdy7SFyOEJc0JWn1VHHpAIclkmxZL
AAob962aJLTEqT0QuT1rv97r6bbhBm6hC9NxBjlqQUKQ1m4EW0xCrFtcxCXFHt5OL/Of74rApc4u
4n1mBAhw7qQp5qOYatpq7acrpgYYd9S8mNprTiDhHEiGpkhloPDPDMRjsidAmwbwNncbRZNEuqtQ
0lpvn8yqKJApDDCpekBcdybO5WfT183lcWxTmZX3EYh9I4Dj5V6uA2izNjGl22DwgCt2rTM9x4zc
r8qpO9epEc0eWUQLvNI4aAtUyIyrYIsLcMDGi6yUtJ5zXQ+Izdv4tPCUpPDeHD8uPPDsz95OhIMY
jZk1ITaACRPcoctVrFmmvi8PpiuXcSqa0eKtvK68pnX6FbzwmctPcAyvvV6Ia1aDBMLfAhQ4bXZG
hFoLEyJwQbgtK14JO3kUf0S+MMSMHou3g4UoY72CmRp5mfZtdRU7WOT8XJ1wO5JOkSM175/khxWY
aiYtTBykiKDn9cfiXVazY7yEaqQMs6IqE2TOVA20m8egyH8/t9AMT1UFyzrLHViaOZSxgQXFmOyM
GYxDWqvKKprO2DAJIkp/U+su4vHV/vnWpmP/QT8hDlGS6/artgrSBQvgyVWqrGQ0o0GpBXMqyqQc
nASVBMe3MwrghB7wmi6F2zcRxpG1i4tW9sIi2eEUptJ6CV30an2re7Aa6u0/+Cn8pWoX+UsLJlCX
ZKoDMb0rjwvnyCeGAg+7KuWSP025OtRmKgxAiEtv7c7OPXuxypCnUghONANXAdfEypnEvu1UjFpV
5pl3PtbBoA5M992/QNNrKW0+4XiA4jr/LZlQOK5BULXNbcJ35gCGKzMPz4ng3Ao8AH+zyi9Nmrjr
hARgwTSQNWizb7WaKYn8YhVcWA6h9wwSLHeayiI5Qojd4o3oylsHOvCtGvPqpzoDRE1Hah7zBybP
pL1nG9yQTzFfF9Uq5RBQ2C7ljoAGdJLrI5XvuzIr9hliCd1NhZzgRXtIFOxtw1bEjFWc9ufrmCzH
IuwzQi9iPDw1Get4jqlz61YBIvPtgggE4b2uin6u5bjThCk48s8r4otskYN+uvtBjr8YHHGf5Woo
Zaa5ft1UiNpQv/3t5v9MqtpfklPzJGFjw7UgZQQ/qfi/dtEP+jK7cmxbLEWbsuOtsNWgPjgQtkbS
a2GQ66fEreBx6wWChCFsbCtqsrzod2FEUwXNDcpN6gALH+d5SILUBVhZYW7Lpvatl/+CLI5CHp8i
1JpJ4NmKYuCciCE4FB9IYfKrLtG9oi/mE5XsFrUvuRF9HgECL/Z52cJLUCgc1TmWyw4R+GiW9JRN
f33YZlRh7+Jxp80QV7YDP+rY+0ES4Zq9RWtMWQUYxOaPN4Okdfv8f13r0FJawGcXTlVaD0tMEoqA
+e5y9a/EOxXq03pvuPxq9iV+Un116hpyNtzhhXknfqtte3OSJnNfAd878SHHP+vS/Szv8RRG9t4+
Y8afRwrRx8xhyNjpjbKTgClCUN9j52CyCSKpHIaUNfeburye12XnWOQsW1zZogwademW0g1vFfpE
lQCjhoGrKHAv7ES1EEAN2RYDnzkulmx3otUEgkPZFYYOl1r2joAOdd2UkuIV97l75lF7h7WQHaer
1pX0e9/Kr2Diwo7dRfP3VKhPsDsLwDOyZCrbBC6IM5wbpS9qfzfezDJFIRMrQ0nXfVYCUKmKuou6
87O7CvxQmcI57PRWbfBYOllZFZRAgjzM7c9F/bzQSEOPzHFCkGOH3PUfQDZ/5NkFc2qP/D6ofmEK
vKl6kWiGhIiHNDknO+c0J4xvBRssfHVCvKdQdk6r+kRql+vGfkMYMzJMzA3erQXdoIkSji7tliYW
xhHTSzUdXr/nRSIfbBUbeKQmIW5wckDtWfwdBFI2j4vMgO51mPIOHYBMEPlyHEO5ZFjHxXAxooL5
iPEUdxCIVEP/Zkr7EngrkaTL6bvs4ZUbkuooDmV1cYqs4IBRH92BJGQBhHdgAucrnL/Y9EGLxJaf
qQU2cOgSS9fUHzF9kcbfK+XQUTkb46jXXCDvAvmGVJf49g26qDQQu79RKJsWOZI8PqK/qWwKlnFY
SMIWWt7nD4ZRXDyi8sxkHQBLBFucmxG6bdxHcbDlujWyZbqQRZRo+ZXKHx23iQSLNbSTCQkJg4lk
n84R9jDVtHxv/dpK0A4FvEGNmAWuA6RBYA6PRIGd5dEh4salq9an4Vie9Pk9Cuqm7g+KYvem4U4H
Xsz1Ad7kFxesqBxCsuG4L+b3sfrc8OOOvoEwndqnswxeo1scwCTtrr/Ru+qQdYgiygjYwEM8SVyB
X6etP6en/Hz/wpY6Xa7Qjv6ij1meWmz+KdSjLeN/83rqlmrDe+VQhsdNAEPTkOBhlhS9AEaWjFy1
RLMVSED5zGiTklhR0Hti+XfyKpP8a1HPqKfPPOOfVUzHxmMHc+nL2p67FGkaq8w1tA84beO38QJe
sEkpVkqx/2ue4egfdwl/LpRD1J5WeqVcZlDRgfi+XQzWAVRIzVjskRmIW+eNo1o5YhHHshkvZSJ0
8FzMwVJsGLbcgzXVsVrRkhLhuJtgOFGFvLsqZGh9WxPEqAjWfwB2uWUGulIqBYvCzhS5L+m9Fuye
2llMdNjexBBd35kzHYs+bm2v06bgBRNUQr65Gd6NrnUBWiughxzAFZNHsPu+aRcN+OoxdiIQBxaj
IOpR3HSsCrNNZFgyPQMRDXz1qxCznz2TM1GmHzqZTbx6Kqr1RglbXvL4MopddHGf4+ByMsdNnldp
2nooeQFhRaN/gCElagTO74w1j5u02Qpe7DwuetShqzxI0euP92h+G9/nU8lmVtoi3lM5qkasIViB
js4GT3xbucXYGd2T2Z2km0MvGI+36TwxjV1JxS5xfHZ5tY6ahJzNQKMA3Dug5SDMK+ttCyikTm+b
tKdVUj8IBEByAgCjcttgMP/XZV5Wx30a29hnBB1iVxazJe14NIrgRAhzc6Ms75mzJhXjETM74g0b
z239QBz0+/a9u3VVpXItC9nhVcGbHDezSr1ytOc60e/7W135oOtXmkJBtzvUq1GvzSWwaQrjR8PG
U8piFO5lnQbLX7y8r6Il1I6mTyfZkyFEdM9xMQLop8Vw/B+u5CVd/l7ZAZnyQ0cPTUP90kmqhNF7
C7t9aYQP/N1wmIrh3tQD9xxiK0zC775+AQZ/heYj2AswoEWdywO85hZW1SbmeMgoDAf/yHKP591G
YtTmZrRLVeUcIXiR2Fl99whe3LI1GW9AuVT9SJvVpL/tZTbBlfk1/cfmX/s3fEtEUn34LloD2lgp
eSCXIYsbzJvKigdpwDpnJaxc7z5ksK70EhbUN2blsUDNLKVic31Ob0S9fkBct3TUJEKhsxNabDUN
8vcj+ZduB0/vovTKqfJiZR8AZNy/LaZvfdN2ltrirjPFXSlQO2xOvO9JBzhkBt+NyHiF6hXR2Hza
7oU3FCIlKZQj6mGEETMk57jbNXRnPJJSdvBEfvUivY+BaCdrW5We9NWMEut1PTXe4ApQuT2TwbEb
cZ30qOOmYPYyOGMmU0dNoPo6a7dFlLSU16tjuy9d3+N0RDkv5uC+36bTBzFy5G2acL4j5Hvk9BmR
xHqpI7Exjr+/R1zJQCMSRVjrqKG5OLkZXC6PYUTRaiB3SIngVxv9usIEdnOPZpz2M4hyTwEfo+QN
56lRWiw0n9NfVhe5rYGsnmio9bb6Z2uh2ef0q/3MTab28rLK18AlwrQXOi8DT4IAhqFPi7l2sRe2
+gmAx3+sBTuG2V8vp0pQQFC4p3hQKXW97mQtd25ZncHA81u8VD/5ZgAO99flSLYXN5SkV/2nrTTM
8qRrigz0j7en4/Cz3SG69RPy+CNbtKik3GufVdBf557yKyTHm8oBkXX9mN0wpfmsCY1TNC0fSqwj
qXbNDF/T1QlIufje6fvN59/lJSHGyz1y6WeDFfgAlwvj6MBY7VVNk9stor2Y5/8BVVThi2yMh6Cb
k9QdZ5Cg7t5vKmJeFEZKs9q0G9U86ZkWuqyTiIz5QgY+QGD3V/rT4iK0hbBsir+cMdNikEZIEise
scH0S6MDIEJNeV3f3M84TRCrdyon/WyNRuUFMV0rvEAPfr7T0D62YalzmRhQtT1jbnBLjSLMRc4V
I9MCMMU1jkJu5VZi2D6DBNbtSoI/YRiwdFNy9wT2JzkLVV8JYIOA/1YJjoMtWS3CutFc70k1rs7V
lWBqKkHTJVD2npDC/258fCDWPliQXWDyTmr5/reoBUvqUprwBAFnpBvKTM7Z/aBs6TePI4V5isJu
WwfxbXLPqaQ4URVEGzWKOfDzwvyf++U75nSAm0KuJc3Fub2YNYrNql4F5NqUY6pDHkzl7bFxFhSd
LREziydbyVXByOMYfoVehSR4WtOaaJNlK/8cE76Il6esAbdtBYNYPTpE07Mnm5x81oTB/u0H1qWy
jsVONpK3Y7yfhOpHxOyDhaYqhg8YIRx6zFrzYLN+EyR1Rw93SweC/BLkm8aCxWlbALNo5HrKsp6A
nWKsuHvMhCaGY+upBZu4HrV7SK1pisvKmc69orZ3QEh34ehyya8oTzN0LmTk3Cvb5zNWKod+XTVV
nKIlORz50xiiO8HhbKeix1Z0V7la/ghFv1HlAnzx55sSTMDA+ekAD8qdLsfBVydeHtWSRj0aCF97
H59GErb30MnrpHgacT2p0HD8gM6brbeYFeYEe+YE3eDfWGhNIK1UjSNonkZQIPJnzSIrov5KLHnB
2CbK4DR5UpeX5tuDMvWb3MVdxCuOhono39EMR2pEQJ2CvLmfk7Dpf8FHxnh0mrbEwY2xnSYd8Dp5
N6jEX2BiXqev3OZmCeu5exDkZGSvXJt+4m2it0J6LTFTlfgjFXYhKfL63j9FXmb1M0o0Q5Z6ZvEv
YIrH1jWZi6oiAdUpDP6SFlM8edMXrYDi0Nap2DEifmcA9J7BxC9pDqSQMEW1wkQiW99eFFjsyVaz
9Gn2Rq/UyerWs6P5/I3ptLWt4qO4S8Gqdz91PLXFluXyqewyWseKJP+cS41bgvYB7slcLxLHlG+P
N+2BtMxVdgDTlv+qE/GehXujJ7CMhbE9mYBXYjWe/d4VIztyreyXFi/noXR+WCIZQxSIrs2VvkRv
s+y1DGCC4xm6lmQOmVh5ltvKSZrv8sKR7ADgPQVNOiZzrdRKLtzVJrr+8V2XY99EhBwglv8Jj70M
7Lr7qBib3HRR1wKaePrs1dLIPREXqXNymXYdQ89BFsLAujrcBVZyjdss0+uVaaPuAdO/wu75xvHz
OfNqIkvdoNxH49CalaUXQ0bdgJfKaX/FM7Yqk3XrgX/P4N8C+zHi+6W/lgan9PQRvL7qKszOMPWa
hSUHHWmGuSHZKo+B3FcoglCiUPHZ5vNJ4hwBTI78BlsW1N9NbrA89sy2uIk34AE10he7TjBE5tU2
Y/L0WWSFXGqMp3erVKXJ9VHR00SsOzUPfqBvL/szR+9YFpUL00vwcrxu++coV9EHn8abFOD5DYcZ
B86VJ/IZP/Ls7TH4ljgy/28dbeya58pxBjpgHwqHJCnxXy88Cb1IQFdRVcMDzxWVDrjU344NPbiX
K2IWv+oZ1GStLkZwdWJb5xzZrQQ3OUnro6W5MKWrzZ+5BoDpEY+OlmnONcCUVzDXESutbQzG5u+h
mFHQs6YwLhpNIEHIlprAok/fspfINC4xproqhA102IzC9uR2HGlwxxmFX2Q/QWxoB26qll2IOBfe
R2YqBY8LWmViQuYzJFWwhNfXd6tvB5K6AFq62WkRBbOc7Vefgukhcy0dGU/oZtIebevpdEvl9L1f
b3bxZwbVdO9dRBT1HCa1OdGdutKT4iOFJwbeE6r7+q4X9uOG+GuzF1OgrdobH1/SOOJdzRvZfqYl
HDetMFvQwfNiIGFQ+wF2cFn6gt/IbiTpyXNDC/x84kKm5KyisFHE5VIxoiz0GW7+Aq7F/FjKUk7C
ixAd7LMUWqDMquVoQnQqCJl7icU/7ooikjuRM3eqrEjDZJ0nv1YGIP2R8m57RTrQgtnCWj/+ifZQ
5GLTHl+iwAPhmyeBKDqrzsDsJA0GMVOpEgFJp15O1MqB37j7jZ0sJd+fhEeNhXC5NQooh8/1UNuO
QCy3RaMoVxns4Z7AKJeA0PczGRvRsAUWXdse34Ra7I59EPTJ5uOHks/oIYN3GTLdB3NDGN8E3Bw8
ZxTyWLP8zXv+IPdj4Okp5N1OI1QR3+HzHpdt9rdJxXGMTrYI5VJtLyQHQpPG68kOF+YPaq2VbYPk
9A9lq/itwC4D/qfjfBQfyQLaxFy+hd/U7qjP8znOCFI+YcppjZSm2AkOeNRq2cddNbmgl1CmoG52
/eqlOyBh8NfhcpJrSuTKtShu9YWtlYl0ASJrJujREFGQXByrzCWo3SImMLR/056w8nm+kpfJG82c
ncq7+cxl8jGb1qhtAjY/Y6VjZuR261d9fxAZcKLpEIx8pLoQcgYpiDZwu23sKXUZemH3i7pfIu/O
aT/bkJthZmOAHGATxnD5OjlNq7z/Uw7aLwNphILfP0HldVPYfBmBCL5uM/79yaLCVGl1hPNTgIQI
An+zy+Bbj7IQppRpwPBf1jY9HtG1QvZsKxzRtPciMyUFV9i2CpG3d2D2IZVbNEVj0BlkM/knFptR
Zm081F/XJCS3NRYTtDU6SdDqqvgBIUFKum7o98/5J08NJEEcXVNt/dxnRHihqa3Cl5SU7FEGNgcr
Nv3Zf3ADZbdIDUcc/VjHHZVsBjVsj5Ccvy6F1NhRZW04P0CenT6KqJ1T6duWJCjRh9IvjlNVfXOo
5L91KmIl0ylPlRrkOlfmcWkHHFcTgHYbAJVprNtRzRF2Emfn57a9WBLv1SJGqNA19j5SwNnFUkNN
RlvOCXiwpFoFFA2+e34M5TvfvMKn/469/VH85NP+SgEMiNQfNxKhN94GoIh1ulqx7vgafmE7q4sM
UB7o0HCANpwPudcfEihdRf21bb2/BSuO8t7F8QFDTK434FATq6+/twYg7Bx5FFy1+xuxrXneQjkU
7yBDPyj+V4FUyzLMoT475xISi2HKiX7nKUHfC9dU9fofD7r08swO/0abPqQ4341kBBhyCVk4ncEp
NNcEDi0O1nMnlVVh/fcJd291p5WSx9M19MuOM1xjZ0nXcoBcftTzcz/WypFEViPM3E9X0Yk1SrW8
Yfh+GI2og+6lbipq0xkmalnNwVm6ygDOWmsPKzdj2C7v3yZztVMiT58AuMwqnznzTMuMEIZNJYCB
qZk6wBRqFKa/9US+m66sUu+7UDqxBqSPmE5/SSwnlCxo2dKMqOSM3bjkVQY3ag7Xm+gWzjy7NR+C
drP86JZM1IlNIOpzMP4aySTf8PYFCXwg8/FLoNYYr0PbeIM8hD3xXN8cYhWMw8DYB5I67eT0ZfBj
dAvQL1zz4/8FUvtOGqFk4ki4Tf6yWYmLvdyi40+TIeE3Sj3dgzK9KiA0gtrH72ybfbNSis4qfOYY
WLt0m1EwH1UpS51KdkB/JxVuWmuD2tN32CkLnGQAPkORC4PF9pZFXcjRC+Nu2udRJ1w6TaTK1kIq
oePgRqy1LMMLXv1x4DDm24TG/HqPZlPfYmEQ3TPpC3o3ViOoQl6Uz7+N4EdruwIaLgzNT8eLwlmR
DmBA9txzUXlFFjpqHQ5rRIPJMAez4DG7EmD+kpgybwo1Z09fuBi5FPCEiHEn/qTz7Q4QsCDMGTIQ
mqSPd4gRmtyLZTcbkYShfQhBKhSljjj43VreAtqPeq18wjFuB7ozvLeqRmtYYksyq+g/xGqq2VFc
UQZ3+TccX9PG2rULyHibwG3dxFAyXzVfKF0tqfn1suzIcRkjQK3i+WOiKDRHXAGWcYkexoExCbE6
vNzWskygpNtQ6DCRX9uuckXsfr3P4jAeFKg6BJhFK6g8T6PyItO1Z/czjXQw93XU5pe6tGjZYvM7
zRa0Faeyye/ATMK4xIGDfZf6IVTl8LA3AQuzx+ljk1/QTglewmwsqdW7rOydbISTjmhpLfbm18z+
WpLytPUFv3dktiX+n3KsZgATnTzid+2qeFLzCZpKyr0kpzOYu6yGrjof1DXB8BezqUM3CK8lIEsK
O39RqtWBapV9OH/bpu1j98TFklUfbP10C8HXVmp0GTQevkx0T9uqYV/Imsxr+4WIOV/sr/HmctIm
9at93Jv8HVvkTz34Iost7vLoy70zYUXcJKYmh3vdNgAcqygUzsIUuQZJ5Wf4ImcapuUaXfOj6r6Q
J0pvtwdsva4XC3paQTOh2zXCTN7kgfnXqa9k4ZGDRFqbENP04Fn1TxnS7pxOyrCdLQnB3Pvj7OjV
qs1+285IGKudJLWMCHOiYCBBmMCoHqVNaKMMsOqm/JwBR68RTd+yD/U6iLh5wmHe5IoCg9ZS2LbX
2W9C218ew7hfBNuQiL586BqutS0zQ/H3yHJ8GuPzyKpkU11l9yJKfNt7O2mUY17D/EB/AhrrnArv
exc/HuOkjKeqxJKtxdxyY7MxFeyNJT2gYAFD+TlF2jd5DmHwlj3RS459LlBh2ZTLQK+8sfpbqHH+
jwDj7SZt3+9iNCeJRY6qUSmGQpaJGXEx4rlGBtulI8XqQmm5RmGkwjnshVdPOd03OF7nxwZpMOVd
s0ELJ4k/JqfrE1onYDSQ1NUQVySw7WqzJlXcyBkohz/6tSfgit/6lraN1sL8dHayLNa01sCi+Oq/
jCNtZwnWEt9FhRGriwim6+tM1HGGrBp9RxxgMeMrWzDJQhamEiZ+7MkgbabXgjCB5nVfoWHtkYOz
+DhLT8YjqlWBCpbh8gHqZ09yYhqEs86V2bRbsk/6oZFX/wklCIyST9yqowlhsjH9dvbmaSjQsuer
HPIKkivhAuev6/Gp/um7znkHFk9yS3HwOSQIfPMpONkNCXF3WwIaUIO4RGeKER34iAMf1Z6K+Lqa
Le9BakZox+xWsjdUJCttlTILul/rcxF5hVYprQyp9rKKLd1i3ceUHYFLlMVWW84AQP033VJWg7XE
3gEKrxuNzSZ6wU3xKCdbINwB9Ah7v8+KlPIPzgDxEJ4jCpafF4nKMY+Bdzn7OUXRanqOpGCLtuwl
zlPJSHrRF3G8JbIsSsL/9Mwt/ffKeM0UY0SS8SYCw2Iij6PHBwhrllmYAs4wX3LCi3g2hc+ZmZ+F
+8RRFIB98hoQNxiwbXJJR7nvGr1Tb5KtutKGffFZHZQQjwxBg1zwa1mtqnw3lpDimt6EqV8YyT+S
45ByYkL2LTd81i+DA/UQQ9roUxIJRYa2MaXaYbfzm5CVY1sHQD4gvLSJ/qgXt52ySuUXzjx4SYb8
A/xPGJ0DB3qk6fttHGp0zDFjZ8ni05HCVpFET1GSOMkjqwkMNB20kGPUxAk8ywE2wCEQ0IOhag8j
bdZfY8rqi6UQcsHeY9uJ6talwUu3F4dSRK4oMIiKJq1GO0tx8pE0Mfc2hFsUGHR4y4/jffuMpwtu
D6qu02kNRs81Sk+49jua3fOzqht70KTyQ6TRgD13qq3lIe3mROf80VhsWWljnyvrUDOiGMYuo/Ha
h5FGfYeFbR+WnxoLNl6VrCp7kR/w+BGAaLAYlW8XevEjf+9YGjE34KGyqmgBksGvPPY9RbBzVnym
UtargzMM9mUEokSJbBpj7rKc9HyXLwfmJRhGxD4mtqyomuOw758zcpNRD4flwao68G8DUw294kJO
RLjZPYRCXPh5NBhZspp6yUjeE1RwPyFy9RZlOik1pebDF7twWlBTynkbtrMeG7N12EBsgvG2NqHe
6sxj5bsYdkLFDQViivhsLgsgvirTcapAl6RGK4WFj2vEIPf+cW5MCs8b6XHBAH4xDM2dZVLPheKD
D7y4dh0CuoeC3FgNVIurSqpBvDF5+PME/zpclHeSCzeQR4JkssYt+l9BTNTlOMnSS0Rx0sZxd8Ol
iHUoDFZtyq5/J2rYq9O5zEpJ7X5unto9C38tUTviJR8EiIQVHCec4R89jjSpnyGAqPPpY9lC/l2o
nuGVE/LRr7vjvmJsaJipyh/u495kLVDSRJTpYbWGwT7lCNm3VgcGsO0VFQNPnhyRsznIkZRTuwnV
xdoIAk1+hIUjVpABaGZxoA2ScYoAHRFmwdxxDbhi5FQKH4jLSVyGX+sEYH9BnXSAU6MbN9vJMxoU
73EYq2bt3dcvwnXhzuudcp6h9iwfP1aqeXWHA6pkgaCbyeDPoHfHaJy/ygTicM+XL6QsxEcCc4OH
a4DoMYYaVPp8on2V9eM4mhpeO0pb/ZgLMeA6vtW2j4WJkxe88PzvkQiyi07ivcIdSWquE0PWKeNU
jHzUlElMa77vh47hlFydRvsFh5YI4Ag+afe3vtJbxkt4B56KdNqr93eVTUJAqa+urcA+beyFmnX+
YY7SQk6IFzZO9g0X7i5UvkOyLXOSK9R2pzNHmJ+xzwO3MDuF8BmNYveq60DciC5KcIs7vrFNzzRK
6b3aaoN3A4cEQKNtfDBy/jfYM0UHQyOnwd0kxdFGaV5Ysvz0ixKQajExjqPx4k+nA6hN+dmO9A+W
4nHcYQZfe1yQV3e9471ibDh0E9OQlkkOR0v58NkjpG0HKJIVqBrI5ZB/QnSjZ6Zbb0y4JZ8QQl6r
+RPXDuv8U9t06gIWzV50sr0pwnroJHVdUFI+gqO+QOIviWX06UoV02gCzsx7H3uxP8YNHLOAMMAB
aRpgZNfVzCKlUeEI7h42SsASAdF8/wuS+3akzAkqAGPZG0vtzmbPF5k5J8rblvW4Mwm7qQRIb3e+
NP2dmLbfzFguebrDnbxA0sgj1WkqmCHEYlju9Pppka6OWfLCcMch+JdqiraBPdfdkFzhZ5bQ+wM9
ZsF8XlUNOWy41RFkjgOZnJdsvIMsTNse1nrFuuXc969HXhU3TYS9Tz+T8ucivFunVwtvYSLYQtdS
ZDj6xudPrXnirarnA7SQLTqbwPICbBRBIQ8Zzq46oy6V3Z/ZyJRP44bN3s9F8uKQhC/miQIvocwx
zPnuDjysN/PtKVPx0HQ1uZ9ZGSMSvRfgy/D4xnKPsb3NmuMQvO6m4LYKjmoezBSU58d8I3MxQzHM
Qx/uCyyZzEKOlR6U6Wevvru9/bNh28lkr8sEzWA05LddIAKqJALNUdVUhRe5oDsh96zeD6FhdrzR
osY5F1t9ENk6Z5KPhu410Yk8txE7HY1HfKk1DidKHAW/gxN/6zBayQvBDMRLAQ+Lx1lNm27N/UXt
/Sw+bdiJQIK2xVN6sAgXN58x2Sia6vyI4BHNggf6NBxroFAJNdCP4gM+zulIRjHRYVdpb7gMVF9R
J+xIUPcavRMvViCr28za9bPo+hwXSbV0YoksAiHjIaGsWqr3DpQd/1Zq22WVE20k8Jp+m+znjVJt
I3sGdZnulvCFDvqPemG+howC25ri9NqQmqRg7A5Vo27OgDgV5qYY8b0Y0Ba2CWIP8djT0RZ0k89p
Q1XrGpLz6btSgY++kQiRNK2XkgQPtCrl43jW5GkcuDnkoQXh5s9ta/gQoKHuPGYhhHtH9r595HfZ
yrXsPgAJzJHmS65F/nITTTencBO1MfMPau0k0UZNC/HBt9C/JwEoM5/+6mo1m7ogMGaO1xc2u1rU
WdAZhOBqSMktmHPpJifFC6XJ0flmD1KdCkumUTrUhIfG8w+72sIK4dxYnnPJWW/m5i++kNXqZXeV
ConhH6nFtduM6oSBqLxM6SikegqQhS7SnEw3KYpDwT+wqTJevYx/3IMFO+shnYzfKXwbWKbrIg+0
il7lsxvUrYyfss1m3OKvePtFqOKOkweo4nWiz28unmnfkuduffKQFI3tqyizB6fFnM3xbvCUVBAT
1nMq3wxKA6TDjnRdn3QKwpObKG9ACZTslPAA9gRk2oA9U6je0mSAWu6wz4j8+5v9NmuE4m4EIYiP
L9PQ6ZCDMEYxvGSM7o07wPkSMSAPiQLlR9x8wujwBdBnAodtM+GoUxbfFZPH0/EMcaWjeR1W4NVv
C+qFlD/XOGWO4sJJ+uKx4KjhhBjgIXBJfrjE/5NFqX7HgYx2R1Vmulfdprafxu5sgYmdUx7D/GPJ
eNK4rTPBTn/5zgHNiz+XicjRPDRFpWQ5e8zo6JiogwI=
`pragma protect end_protected
