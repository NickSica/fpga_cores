`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
V82h/mp8FbHcv3//3zVZ5VW10Mue/LSt5dvjsUkiSGtG5WaH8H9Fv7j37k+xy+3/pQvfXcpqBF/k
iaz4/vETUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n4WSOWV3uUjyMD/l4IGcKD1bHONRRplCKgax9lu4YRYlORLHEpckVBvOD9geZHtnlLIjTLNUcuHS
rc4oO2K5x66eEf5+m+hNzaPYWCrVKWQI7/tyX0imMAsD4JQXzU2CP3ATsQoldRyYOQZmggmbIMiB
stLQ3uoRuVc4t0kXI7U=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zgo3FUzRcS1G0FRTCr4C/JBs44dp3dv5CUvkYU2vM2fDyGtu9ekJcjDXnFGi3Qx2X0BV1gEyWxsJ
xqQkFlu/f/1mutspkUjOMtKZNCgPGDHkGfwBEPN/xT22fOBwQJUR+Oj5KSeDWe2U4t5UJ4XXcGMb
ZV9syPFreDWYOTWkkl85cAKcf/WXC6oz+tOUowqV4nSLA1PaSrK4ohf8oaOGNVX+4Ji/w6ViTIJJ
OqmPJQ151npm7Kbt4RW80tp1OmABkNI+o6h4rwtTS1IHzM6bJ1Krrp0V+2aEmmqoZkuKINjX5Pw3
P4Vi6iUmJI0uMpdsCPr3MEC8HH4v95WCnjh0Qg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A45QQ9IEoKpoNXpmniz3AuFZmGAAZIhtA2hP4/pi+Iwurx8nPI4ZkKpYXPnn4DfH42bSsec35aiS
Ve+A8f1Q00bmFgtclspinRe4YgFesk40ftn1mzy6g6sLCNXhUm/IIjCSNk+ie6jVQS7STfOdio+z
cvSm8QQePoJjzlJz/jkNhsD110PhDAevJWb+C5fforY6kT0k7ZmJmE7btahod6wU3o7t2HM6+XGU
DDNZ5E+RLS+IiJYVCOwsdqQFDuRaWwS0k8Mk4UuDiVWtU0+QLFZ/8UGJhy2ZDSYlL/8TrrsWcD/1
Vku2N+fkWCj38RSMWEEe5TmUHSSzP7uBI6QwVQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b+wEsHDGMmVXUM545W/2toIjDItLsHFsIOyFDid8Fv6KhzBePVZlc9t2c1LfdAa6UEpdqcx5kgIr
+oVEglJG3R/fb6dRp2mvlu6+x0AYh7FK0My5t84q7uKZ6EPBxHnDds9FLGQdMDUFv8E10WtGrG31
lkto5q+L5WLAzYgiD3//MgdbP+aqLc/75XWIRhw/PfRn4OqyBU7xSBeoK9TDxBwOscUv0cQ+dauJ
dUQ0W2ZCXwF6cP5c47k76Ikfu69J0/IO+FTLKMkjAB7Wzsyqbpl6RMVdJ/iYscNROh1xxo2k+52w
4l9VnVKN7wTWZdW75B3V/MsNTrKb2I6dBdveDg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyn/owx08GdB/M0CwlYM5XwpK1DLRGgNdNGvCa53fvz5ftb1LM2R7yhWTTXlm8iqXlg1S70wvPmw
WVO2ZNZ0csmDdQcX4HNMiokrI2gpR08Dk8n3nzdOhqyFyh79/eVJzQItyKMQmJZNCvFfww0mtX5K
FbNe2x6ria5jEBEBp3U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J8WwILioFJtk4e6vNsFHYZhWTjvAMbsqHcnvhYKYzsY6fpaoYuWnjTNNNxS6JYZj7bKOFgPjdnBA
rKaGPLghV6UU9fx6UcBVLjNOj95AU3CZPEjWGC/GqjGRPxOkhGtDka91PZuOBRTBqJT8F+5qIgQR
vO7WJHaKezpaUm2zbeC7+ShM5p4Wm9L4dzJ1OuUGZNm39p9FbORAZNzAWa35wpfJ6PPOgATFMi7Z
sN0Hg00oxMFCKSg1bxvN3p4iC3rVT+wV6yuzOecq97B7Fu+tfvP+shqnUhodTpF0WYfGWHeK9ocM
Mg7nt62XJybi4Tm5rgYGMIIM0i67934etK5Aig==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AF8EDKLpUnsf5U27caIfzjHsL1dKCT4FvrlOxjBwD3ZJ9vsXwbWO+EJTOJOFymKnoSSFnuslr7C8
ZCAbkJJLJrLXJwfvC9hiPRksxuYzuxWrtwsjJd+5KWtue3gL5kHClD8Tbo/V+Dnr3gvKzMRNdFRz
i+4p8dC6/32xR0/NITJMYT1uOYu0oBFDHGLR02Wn4PqghcTR3gQMVeL0RsDhJibeNnf4Q0NsKqCF
7OscDpis6r9ZAFao+mdpLGI93rreTlZvJBUPh2RcpqOjL/8IUv0iM922KOCZ6j1LtvD0igXehvHa
5hOx0DDcMjOoejqJiwIqLij0FB13lDBsu+fjWw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 129888)
`pragma protect data_block
BMP9G5RAk03qFRu5UmzfhPRa2E8EtqJjN3D5ol0ioUjHNFu5U09LfZJLTtZ2WeKpuNopUgPzEZau
anpChD9EnV8nm1MLenTq5eHvoWB8v8Mw1EdwONhAajSxv/gGFLfXNRuliXucexLG/rL4QTS38KTs
gK1rgT3LK+sis2Sn5Rbh8AHQNr55gHoEmrFSt05Rc5LTSxmX25sHFY+oXgX+JbBAk9VSxOW7Wxtu
/BO67hQyA5J2wAe760Zb6pzAquexX5tIji+h2OuVwVkMtOvCO8SezVMBrdlLi6SUnumXA8FT9UrE
Ju7I3l+G0ekYY2vl+AcCy3t/07ReHAg+8XKcwQ/qC8MrYLO370PL6G25zvVo5m8ytn4fs6oqxn4A
g3TwHScvhI6zdoaWIYhw+uR8EVd+lpIaljr5q6KqWMND4U1J1x14QuReq2VocBr4wpnRzPJSuufE
OwtFrzeySgusEAZPzBNJMj7CAHLrzrqPH6S4c1F80xFy0kvvgAwshzxNezCdgIdJ9jBAyC2psArK
UE8dEhYEAgDrLBdsozzODa85vSImMFl1HVHI0SCNBhcy46Uf+azIM7jxaZ/8t3h4eT2NLTn9XUW6
yWzZuv9PXZ6TlWyTN22hnCH4niIfUHQ9adVZ0BlhT6jSf6eCOCs3PMxr2l/lp8+NYJreK5/ljSvw
iTE/dU4OBcqg1vRztILNPj/W9X0GpaEv82n1kfyCdO/xM1FbPyHlNE2I5r1KINAcFG8Rui1JF//c
zVPWJe780Tt12hKHwPYvyBrDCRggFovNtwy96wJICgqYguaQyTLwfAWiPpP7rdIHpTzAq/El3OFm
RojwY+h8K7qgpCd2VXtSirfL7SJg2kINle5b8ka3r7HS+grvub1Gm73Vc8iioVVolkcDJzqHfDP5
gCMsyM+8C/q7TsYAQ6guslp/KXR7F/KvOYFObnf6ktkRcsFhZ2JB0gg/oaD/cSvn335V1LgOt8K0
wp9SsL1IrzSrFGUh+H8rhwHvkMoKI3To0J+Qe1uY7mdonlEkxgDj3F5QpVqdC4nZedCDoBsf6Df5
AzfYlUqtIk0FJGJV7cLvaSgeztMpLw6RDY9Y+EXN3eCviPyQLmTYbcZ3iRUQbGU5lYxMurMtf4Di
RjTqJUPM0jJMV6kbs+d0WwCcX+5bXB/hszbuWqNe5foa3ytEqVn0s8/JccaDrc4uMa9raHVhoxTx
cYvR4bsxcjLuaGjWE7ICyYKUsCDq+4+3u2IA+knaMAyf7LL5ZLoA6u2/WpRQPtIaEj5waEFepxxg
BUYCI1kkzZSxE23xa7bhg0YvbSKZ3PuNoxiU1m211IZETrqgwA+rD9y/0vOsaQpKjOOXwr8n1fv8
KT+6rIRcQ+GPRdAkF7tu+Vz7dMTJZOyz5glbSkINCmy/LEX1HPkWFNX5JPwmDgfYDLrigb9Zm13/
qpiiRfQ9zGixjyUILEl8eDvaiHMQNGMBQvnzLunGEfmyaxTPg26nagTrzeVosb/ZUW5bE2OCs9US
iVj5Apj+bIn7H7mo8Io7VcakwUK15RXka0WNeGqSrdSKUJCtQjS+FBpVDnAVZXfxxny0MT38YIYn
IiMVWRBXHk6p76tGoFTb7njOAKIHIRaXoTSKeWw6Xn4fQRTIElyBJGK6yHPSCfuI9IXsjxh4qmpA
u4A2kknK74FBcH7reJfoHRxll2Zd6yDTrq40labvqvKtvkg46dToszgNwfKPf7irliD8Pv2mxxPY
eFkKA0Y0tXtucTb1RoREaJjDMSWk4BtHGaM76gEFmgHZuc2BzuToT2Ga2zeEXxZBgyb6MTM+B8+x
H32maH/7hOHEbYsH+p5RoENdQ/vbQqq3iTsGQ8EMW8WSA2lIXQiSI6AQx1D4kIBS1SeqH1Tu14gH
LwYZVEwpXKR6Zpc6n8sLDOQHvzvDmPlw9+DvYaziBzP6mnEBawxcipnq36c+4MwQSHiipNUHwVYx
yqHLr21w0MZQcZwjhQTVFsJ9DAuGT32Pg23hjlnovkZjEpUs333z21kYoSXFs5fZ8ATRd7cB8NOU
Tit9XgM7U5DJ6dEJg63/8EDRa6HXJL3sdNKmyKPgTvlbtThEKi4DjRP9GyCffsQ8nAWo9M6MCP1f
w3eyh6DoJnVq3YW9GzbXnzM/85NqUiM9+tt33RbYNwZEWgpeDt1F1Rni5QXWANRHlKsbfOwKo2W3
oZBmaSofiVwIZKu2aIeBt6znDTEU7nL8+eG7swB/45SMEyH2mDnKfUUo2iYiJ4K9mwoz4emXkgG4
4aL7BI9pt6feexq75ebZccykNO5pN4iBF5ScKGrKtBuxGkCMJhfQO9iSwt6lhqXiBMn7IveI7KRW
ixNG2guhIuJok+5MTLcXjKW0YkUSz2BAI0mq05lRXKTmNBrroVWKbGIg1zWM6Y8uJq/TyTdvyWHF
II+C/LU4mY3jc+b5zqRHLN2R5RYC3KGsrGuaqLtBkItWrwI9hQtAlX4X+zPJl19BD6nzdUIfRo7B
6RjDDag/tXYos5JM3ttQs/QCkdXVgf4U0tszChcmaodpmSyUOJt5m7jAqUYcYtjG+wO4sNlSKAS+
b9+P2uXSchdw/fnXiM6U492troQbL/M4rwYU2qJ6cSB4uvfQpuXNfdg6k4GGu8IgB2y2iclgRKc3
+2Qp8A74M9bd1r779/ItBoHzHG/NXxCBlhVt511hS5fcj47w0HcgxVtj1ywxJel0mfpIX1VbO4XZ
lbTc6gWgyjB8lTI8jJ2XeRSlCFx29hOLsdWCbOgKDemWqpTVnlqIWGAccgIBL5qvLobF/51ZDUV5
feIrAlStjC0KzgGOdMYlsJXpN/3pg2LuD1wSRsgNYedlHu7fgvx+FMBnPCMrN+3n1kVDkbDupozP
tuS6NNxFTx0i5o/Uq5KYGEY06JlhOFKih4jdGfWVYRnxSWVc8YhDj8eEMPHniciLUXmiAok/oX7P
Tz0vEfPH7W/dlZLZ7Xdnm4Q/3LCcnGOPEnS0J8RnyVqtxYueiECSugUxrZyu0589HPaQ5aQXjU0U
Bm6gxQH4gGg2SKxPi+JlG4A6ul62xM/kdy7X17v9tgatIh6Bq69F2ybE3N0BgIKDg/eVEIz+Q7Hw
RCgsmk+zRzWigm+Y6+ou6ZkKM5GQpg+/fhKqwND3bZwZutu14gHZYbnDtCHeKoxC0BGbYeUIHlWm
OJ2XprTS19lzJw/hsNQH0H0jf6h0zWea13ZA4LkO4GfmvbSjtT1lofY6+vXbPTR8UsdlY2Nd8m1x
4xYFZxXpUxFoM4TduwJyrpdbd+A13+sF6fdjM98RBqh88sTHWheuRePUF/UBDS7XFJWHykgo3b9Q
vdwlEVHIK4X1LXK20yGbbwRVdSrepZPRKj8tfXgBhXcyN08SE2y3uG3t/BNiGUlABpvsZjhHAkQc
4jGWvxvW4cWrSEUZpTBY6mtAHpt+34hwgQ3iuha81o6I4gORGXsW8hHJsA/x8RcliIlev+J+8HeT
FZSd05mFQaSLdeJX7CpHGzNm91u3RnMV2pd7qZEMx0/JWTowlXNmYuRuuHiWSpUSTgSRYcOQFwxe
HHQ7M0cKvsRn3wq155Z/eNIHBFiIzq0lYJg1I2tgbbrBM3zAFh372E54jCWJyxTm0UB4zeuvgXrb
2JVPTbuAqf+YuJMph49zv8HCoIvxlKfD0SzS+ihwggkHG+/19aG8S6P2e3RcXN286piOelqnGeDh
vVGvRC2jm7USJOIHNfwrIfGTgIriyAjcTdzgX3pOKNPS6Sy0GNDI8uhCYz0ke3lqUO3BoL3pBBRg
+x5T6bRi0LUC2duOgyHejPgLr02Av2bCEHJJX7VZT8MEHv0TtSOHVhYE5JXwOwxYBdHLGdhqEGAW
wtkVm6IvkGfIKpywZwYrE2auX9x9Nq0yungsCdzWDd1nzefPvevPRpLG1c58+lHA8WHYkLNlwCwG
0RMbiSNr6swaJpsCn0eRtCm3PVBgkyFRfDQ36IZmbBQavxc4p/Kg1uwv0/eo8IhtZw9iUpdk4qkJ
O2MMo7MgD7xzBtUqJNNlGLfm+WlUMwA+6BkmwcrQT00VlVB8Ccz4zZ9SA7TBYeoqa7LmDXuS97i7
pZCBjF9vIyB6R1NLoXJ2fPPZlGmYLSkEAtMBtd5cxD/YhZNEhCbWK8M0PJcxm/Paf5MMjemmYruf
nt3a+a4pjWpAxl12RjlAjjm++ZM87pUPXTIDp721mRB2TmA/LNNhOrEM3m8cIs5jHh87trF6QwOh
9oggUFkdLejWVNWvQhhaVPyoxMgjqIneqA6HSt5iUrfeDEzFIyRKUQG+9gzT0ye+V1YK0pRFJIm8
wkCcmbcrX6c634bj+NzJ5Wl0r+rwml8kWtVC95g9NriOVBxKX7FRaLavtKBpT5a4A9ZaAzxKzwPH
Xvd7R3wO1m0ihYHABkOSVJvdLEcmozOroQCXZV9VOB4x+7LQ7NQtRRbA5yjjKVMj+167BDN+R1WQ
OI9ZrJbAm5Iqs+DTI8oB3JM+LxSZiJxXiWV9ePksXDDYPin1OPuqXKAxwmSWlObvZJ6+H/B33pdA
P1PBEQMn+xYuXJdHUFEMdKcLjOsA/Kb1m1/afyENSBcOULWd0WgZGCtwABWlfop1AJYp8dl345SV
quH3hkar8qWyeBDzrc3SaOCUj0y7FySUCbHkCnFCpDEsGJAbLG8ecMgVgyuIDtOmhNFPhm79u4BU
a3TQGOXi3Y+P6FGwmuKBZGnnyZUXNRtaE+kwToqhFo6zqCHF2hKBxRTPNRLdYraKOkb5yPR8KIvT
JJZuJaluNfQQDoun6eyPdaus3Ynbs9YruQDI+s3+hM7ahSqAuy1ndZT28jTOczA2jEPAaMU9P54A
XArzz/KnfqqFdc3Je/XrLFowpeZsYd64XCAOCfQPMfAbU5VS9fYdPODfLFnl7uniAsdiUECDELXZ
b1iob+GzHqpV8qBkqx/HEzThcD59OOuhaaj+OKTuuczJLhbXulnyAKgpLqHLYEh04X3rf6GNP2CZ
bsQ/zekdF6tCjaZh86z3OyJw3edH/UYjOdm17g2LvE0BDUB2MumoyksN343KWfbnkY5OhTl4Eimg
L4lpTgd8fgDlW01qquHuXWGTXJjfSKmwB57xGrsyiPvPWBVY+OLwnBBOZ81UYZ/EiKRgD62ZKGxj
/geu9gSdduC9/cNZeV/Jdq58H6v6UodGDSgwPMpTTTPx/EIqQHwLWi045YOjt91hZGhaJeDxsEQf
BB8seKU4w9uwCFK0lKPetgH+smDIjoOa/mW4lslwKUiIVzlFoL3NkO4vrPv5qAfc3ZwNzKhnRgen
xK4GMM3CVnGPZA4D+bSUxt86L/Rhrmh3XQt5xGv4Kp0yVhFHOPK43AP2je7Hd3tlSILZSCjeOJpT
zHxXxRCktZnpeWwJYIjPFKJSZsnmL1hIWaIvjdHOOULbcalluOMHzkPZhEOsUjmgbTe5dYzaysbs
uQPJMbEwxkypf9Ceudmy6hd1UxE97IJGwVzaVgCJNcHULAk1C1rIddqHepRsJsh3htVtkcTB1Woz
AQgV53pMOw+wjjBxzQinLFT7DFrTPk7+qa+FDwG8UAXTSrcXnORQD0f46FYNfBbdpLizHO/Nvn34
UuYN8VoaMpRKRz1DZUPJtcpZCieHveBPb3lUp4lSToAd2QOTYVKfXHF63H5uutwsyaSqEDOk0UhT
Z8+AmsA7lJF+6JD/EV4UGjxz17sbb6CpMsOXYP3DDeyRH/KfALWkF+hDn/6Nqzpo9t4qR73cEMFd
YYjHvuDaKPJxOYtugu2Z935lzmvhLsZmoRJJDVholrbGNikZCUe7RRSu2czSyPmH7EMr5d1RjphQ
iv7Mpgl34Sj1AH3VnIvyqcknL5QJdsQsZ4xkbrjSP8Md8PqNpzPZ6Gsuc8ULsNlirm/8nZtNp3Jj
n+1rOGFQTtSVm/mEKPyKvHsVlbuDyGutoCMRdVSdFZg22gEmNkuOChKC+Kkaog639Jj1IKen90yj
noqTC7V2bSlJB9JiwiZND7hnjxiPpXPFqnT3YrSzBOZGKfykJamr8dDoJ+riCtkGn0SgxDsdu8Eh
rQw8R7wR9Ox0QR/tRanJE4iRaO+bKgGexjVA6Dgb7LZF1vMyAk/ZVlD6tNDVaaRQEi5CEcaoH88P
EvEwiBtZHnQpi1ZiomGh2DLI28WJfE/OyyDufvGj4nsmCAqfyss0Exq0QZMJenB0O0kRzQf2yohk
nceu8e8guZHh46Ruvdg7Mu5dnXRw9jqaDIo0oondKYjPHZnAt6ryh69K3Ig/peGgBBOBqiNT3/ra
UQjpXWQxYkItV0lIyV/GMy2g31cF8zSwLorUr11B5UleuQzGVJp4mrE0FULidZ/BzWSehNjoTE5k
uJyGe25OIbZwjU0DvJacmQZ1JYYNPMsovzAXlebgoGKDNjSDDT/OFhATjo1lxElKFCzvh5dRSi1S
Auma6fq+6HL3GuDtp5DWYhWMpqvyKGB6oIr/G7YKXW/VVa61aFSYBYVeeI2I33Hj4Lwxr4nbSf3m
FdAj9hk2TsSlwurKNTBKk1tBWkJFU4AbiXD+5C3Rq2ZQNC6zn3b42UfbfdhGrnUXh52IZBiaS9do
qXtj6A/s4C+ebH+L765zjJO49Muo1LN6AfIh1+aXpIcP+rV5V+htx1Gfd59YfWcs03gbRERuJaxU
iUbYwRMM2AcbebZH/nmDZjtticN510lckBTsIpnfOKhUPXAPOfbBm9BMw3OlNdGuPIagKf8YQMg7
i+XItDNYtWvTN+oZMz2DfvDsupmndxAP6V/t1h/pEb3tYzxAtCiq0jRuFSORJwWVVF0VXJ3y99DF
pYIwucGZJ3aeHQJhsE6Ct80BvBN2n8UVW2srR2rEYRgye76LpfU3J06Q9pWUWHULA+ow/HEqx6gz
r5ODLJG05M73xp+WAYWXFTr/XZBQF30bx6lhCqgFxzpxB7TlPHKMaymQevR+8++dYfr1OVhcOfzb
ygJNX6MGSaabc9SSpFgzVwra+rH5QoDDMI47/2Nv+sebZwrcItg/pCsJSAwzCZtdzl218dO+bYS4
4+VXnT8PCnFEI4I70Jj4xjNE8mC51EQAWvsUkk+gFnMNA/dM6q3aI6D48dlvFZj4MpKgvw9YSx20
tzDqHWYnBguf5H6bo2+qKm/mSrB5sAwktfNB0gva3nKY4GW4JRLWgYlaTWOIaBd4CN5cMgpNj738
GZdsoqXpZlwyzyP4xaLcDIwEA/EwqJL/ucw9vBHvi3aqPAIV2KioOtRKElLsa2HtrpNsJzL89nIf
Mgbn52BpVQlooA9pX9EygucOpOn5hO65IZab6gFetE5nVfCH1U6hl4uiaQHhD15vYuszPgiEPDBR
xOJGJBGzhAOadOOkDKmSmzbqCMVpnOJXkleiRjdzI+5m1bVYekJnz29zW7GTpwbPfLEve7hjzq65
lYoOvgZKk0hJ8CxtFGpDPZ9HMdum+jjRmzlkL515Kx4h1y4rEfV0NTaX7OX0vl1Z6VnxIZ/nBt4j
FXxg84eghKBqGu/KpLNV5JZUnotrxxLENaUqGTfqD0BtfHkCHo+0prz8tRw52Znh4ThrykqKR4Yu
uf0IwvdOxeEY3Pf7K25hkvkhnGHyDuztMTwi5l8bs1ay0R2xPTuIHrWqzgNxLlVMrL8m5rrZw9Vz
4KOP3+0nnfzeFxrxIRHzTUVBlLZgaRCgL7LAFidltMkA11LMo+bDh/O/1RLcueslJ+mZhHklyvW9
lUixsoXA9MYAIpc9aMTYvdO1Kr8WITUacVenqjo4FwMzNkh/qcY+LA1B7bfWlU1uQ8Ipt8MsKqYW
F+/vvkCJ9CzzXHquclk/ZmQ7cjNnsPgZnOJIaORO7RLHOePZeI3Ohnh49aqfMotDgDb4mdu6/3cK
SN8JqRE7jPFdTDwm4igLX6PTuHhpTwKwE6glEZ5/a+b7ks5lkVlnAUw6sYWLuxm4hqZ8obZnWqQ/
AFOl0BVtdgJdF764B5+rmjIEF4pXLd7EhLryPDcza24PfIgY49F+RvSpND50IJBqjZVwC6DL6KXw
1fNuEuTW2r0vkzYfbSYZQpWSBhGIAkyADOPdaLn+8UF8Jfgl+pW3leBJifNYAvzuEeOPDIbJKCdA
mXk//c+UgmZSP4US1y/xEaK3Jp5J6bBsdcadmzhAiHYZyg4PdITfyvqLNOi9K/WuJGLRr9h43B5/
cQ7jJIOWYwX9jnyo+2xmxPPvPcyQfZp5H3oZpxQfvs1hZ5Kwv0biwp37Joj+tOGpvoqb6olsUkw4
PJ6HVjtXs71X9TjczFU8PWJWTNVapXZE0nnhNuZjb8DLl5rXNbcxd6c+O0/jMunLiRtKhhmjSqsw
lS04ff8HwltmOos6l2t+lyD19AQj1dyRi/GtRjXa9Do1zPzFVlxztvUGO5MiafMxPmuMH5vFnOYC
BmR1Jt1rN6qWR3oRiFrCScNm9QJrQFX6YCZSgZQFpsw0ikxMlSmmChK56+8yTaOPwPp7SjvMgfR7
6ZzLh6fcqxcsK2tKpZc9KcKVoU2l3YVAoCLayfWtHaECJghIofA9r3BrVhEimh1Ac1EJ4ZvZfL4v
xt8ZBpozVYBBT9xqCKA1v2TuB0do3ug37lC6Q2jEeR/6tLLgDYVkhCQMSIgZ45jRQKOMaNGrYNf7
G3+JaqVgNWW9Z4XqcwSMkYVW2bD28MvsQIcLH5IcqkSePW7Nn5r2UnQDZbw/3AVmKvvD5lMqpHzs
w73VM4Lw1tp3mB/PJYgnwxKpNrrE8nP5T84hHmeVAabGJYO+zNESaGUqi34jyEpHduQW0kykD6uF
j8Jp247P4J3irdlAaZ3ynxGuvnAmRZX+b26aOoFR6WYozLmHtOJW1PX3/4rgbbD+OiWXyojI8v2M
6MRqDHh8iuG7Z3MNbY/LO2W6Wxt4PdYOVYz4oMFNJcxMSB+TubbiX153d2siPp6OQdgZvmvKDwBp
ks0zvgS+MZAMiwZWpTAl1Sm4kU7++0Lwj/6jqeyeiJd9pE5S29CH8vZNDyWGskge2yE356teICHH
qXvdrgc13q/AzNMg227n32FUU/U5KqlevhH55tio2AWRpr/pKKOcFgmTuJcBvhhZunfOqbHk11Gr
eGxSEFIZ1/qiJRasaMPSb9m31t4LtyN5ib+5Kye17tbe8hW9JufUFOLs66MU8GvFhqTz7EkLdSBc
sI3sOffF6nOvxDU10H73DXzezPUURuHwlFze49SZGvUURNG2YZ1R8vieN2JTRzXg36OHxw/lrgDe
TZOClgenK7JqR2DKpjeDv3pYkcQ2E31V56T/apZ5SExt2fiDt25gfWhWS7Xj7YXCvHFY4zXqvKc4
FtUK4rx8423Uy6DwgY/FJfFUvUdb0AeR98TgI+Ra/LFJed/XcjVI9riwzs7ko6GyrwGBWRw6IKHL
j/obhcBEe0CAfDKMtEi0G3FowTjZawtHy/PpPXgWkaVKgvo0ShF25uK5Urwe7tOmJZS3y2XVjXHf
Mq5dUVXx/7clpR7pIXDcUa1SG311FAROfhdCM8aZMcvnMkk8xtSFpBsvjGIZGCNbfaPN9/aldmux
RAZMQiek7VUdoCBHZ3qIYowYENOCmXfsaSnUsptg0kaUlCL8gdxMtgRILRDm3YdMJp1IAqJypwdn
MCRYGS3c13hsjAxYU+UBK0qMDEP6nGa2LzgpripuuS/6Gig3ECjJrifdWp4gsDYIQBZgWEbcKeR2
EpPVVHHPqg9RfSWfW7lacunuc8Cp466qiUU/gzB19hxgih9IlLksXkp/eZLeTf2S0wjwik8LbGVG
17DBfxIKt6720cTofvmpc22RHM7jk6qZe+mNw/W7fgRY7KyFzMOqwPwdyH2ScX7sPbQmGWF6RqdZ
vEhNakz5No4ePYCgKFqPU5tqqVI+eQ3j+jlwUuqE+Cd0Wkx8myVKnShNiPyGH8dN+p/KxBgcTcPb
RXfLjmEWxqzn9kXLe0UpibDbrO2XPprEAJa5hZo4XomGvPTg0zlewyFOKOwveZs7A9bs36e54ctC
RdKT8BBGvxJVqYoayFMmPlafXnicjKQnbTJ/bx9FSZTqELZ87loABu2ksqDC0hJ/ljd5ff1RjQ8M
TmRn8dEe4gO+LbAAOwpxz2qa196yjxUU7LTC+59DwLaL7g2Hg5bDwIkU9rCKagw2D6KK+b8ilEga
rDCJp6pGbqFC9hfZ1eFlCeug1a2l9BQxIrMoB1vRsSMX9v0a2ThK4blln7vewV/JpRf42rCw0bfb
XaZLYVDA8pFCmX2V9CJt1g49zyrn/KJubYb1yL8Dm2jQEhoV8jsH/lY15ikCI3oAL8k/cbvEJ7aa
+USExY3thzx0do9/tZ/nVQID3HqWtF0k7etlGai2aY+VumTpM1gHRewxbwkDAlGQkE4fSYNs4Efh
qV1zY6CjhhXVp3lEq8gZV/lj7OV5R3SN1k6wEHorhIvZdoHSQ2EOsr183WR0C+4ZvtAZxW0ULhJE
X4bvWryQwZgDWFz2g3pmCWL9/9SqPw7hWO6eXbWoUd9JrGM7ogvQRTLP7u0LQjJHPacRAznjaHeW
Or7q8iFWSs2qRh63clUxOr9i47ofpf+6NlHb54A5V2CeALWbdFO8Itd2BAWiYqAeEDE4zUO6QOaB
qo4sDgwVFmCUD1jbk6n1PhoMJjKua1Uf76zY44flCktADaCiF8r5cF3NwWR/ETuKBH8SUKJD+E/x
e4VFs4qWhiYFwFwkMfTR2DqnOIMETk5TTaNBLAGhPaLcdm5HMD8KA86yxY3bCAEHip5z7rtEuj8h
ZiEEjyjFjdgBO9MJv3SUxBmNQN8lhs7ZscQ676aZlcRyMVGjVcXqkNfuVb0fRuulHNHykRI8/GZO
5t5aleIKpZzs2PPMVwYP6aDG1KNcJVu7kRnTxvBNmbk/+4AFt7+0bERD3wqqs7VE1rxxxLS5S6dK
r1u9BUKIFBFuwi3zvtioZXAOpCr2FMSNxX6yvi8ik2g2VwgFycvoazwff6a5ZdATAk5w+KXGTntP
q4UnVJ7zCGtcCTO7yF8pScsgvSQkNl/jKu4NeQP7LZhi7EZ1rUDnv7DuM+2IZ2eMKEDfm+SWZql9
IGbWm+Al31JbpOHCFTtuUY81Zdp3ykze7GBvvNaR/NOyr0i8o4maYnlNH7JljfZMMcC1TIMS3T1j
Fd3mhrq7GcC1Sj/AMmp+rSgIM6kkECpT8rXfFHYuAr5ycYuGX5hBxQBUYswWyOOgJcUEDaMY9lEQ
mKiexoLqUt60Q8qG0n3Pw6Xle11Qwy/vUagE9dBkeCmGsrY4HKMi4tK891oi0Svn17K5EfPlNxPm
Ocr5MCdLvLGYOi6TWCoimvEYgdcjxVQElSgajMf8UcIPg2un5loOkbs91t0lOAiGnc4niqOQIpVd
tqVeOLJYRnSGvz7dDe1fhlwNJZGYMjnejNkGJQfbPxusLf3cnHWp05OG7fOCwLPZE+nSQO47o8ax
Xdmgi5ZJWqiwaIQvteGMD2hIjJ0iOPnXPfjY4RO4pReVRN03RJQCFCNxCMLuLV7VKRFXj7M593Ge
YMJuhbxHLJG8wvX9Z0yV8xJeDYBUjxJqL8zfAGap5KIpyc73SFiqXb2keqpEnjqd9sJ/KK8CHDPf
1z4ky0EgmLgkxEoaEEy8yW/FQAHXv/Ke7jmqwTc8viblrlK0TLC+u8OTRVal5qz8TcmcBtqRES1y
DijC1Q6QpUJO5Uw2x6b5aH26RGA52/5y9O/3E3P13oy/KPE51ld2SPJccSwXHHHcs7NMgF6uhbCI
imILni9iCueTV9aiTSUDPZR3Sm/SwL62oLIK53CdGJp8pOCJDvwM/Zzmcl8NRAo90nn/jcf3rvR6
etDnsWzPq+YS7zpxVmX5zA6BrayVCBpL8D179A9r/+OdtJ0T1vX0YTzXI6WarYKpewwtfFfLhWst
SOYi+0FzDO3j9Xe0l2qhekfVGUtmUnkmdhpP/cMQuQCc9s7RthGbVxfkZP+eP/Ah/Ci3ETQmEYl4
GkmTFbXNiPcrboEl+5z2bh5QJWkWZl7Man7Xs3OOZylYP3Qcsj/sYP+0KHeuIcLeCumdxAlXZXeh
A+kESe6b1bWNfSaoBbokCaTbOIL9Od1ZiFjJQbuZA/XqJQsx6IjtV+3d1Mft9juADPkHvfB6mRwg
HWrqHSW31vTjuSJCG+Np6CCkdfNs0jGD0lxI7EhAtTryufQQpPj3EPQDym4i5ZSed9XN06EtQTsa
CKnIdsrBGoMlqd3f+T9jvc7lN1KdMyxCtrZp0/Nkls0we5YkMydJEtnft6IOax1OGifCmAFuDUn2
O/vpceXVi6SokJS0fa6NhUDbkHrNbEQY1aG73K6RWawQnUPuM3SiqtDzkD11WK2Kkys9gO4DKr6P
mkFs1KulSY5YxfNygoSDBUGTBb508xk0lAZpQV/aB7awpB0Z9OXIo4HAWJ4f8PkXZwOOtjE/oaQB
MrK/LLksu3mJUWjPfzxu4dQw+lVPHE1m/JLNwsrZ/AQcljuJFkJj1HsYMurPYuwgvwb5x9rrTDwa
COnCUdgUs5UP0iXj4kH4j1wUk3FCo26xwkNb0Rkwh5M+lCMgsi2eBa6eiZFiw2+jIzNZe2HxOjQc
e5uQmc/wqUKHYn+uPWDhCZr/G3iRIci22+m9/UEms1J95bYxhjCR2GOSPYKwIQV6/DRTZXqQaCzk
SZcaScr8yJpgKCLZgbxsZc7uNLktLJI1+ujZJcFeH/Db/crMPF3JfoXwtH0tlLjFZE5pGgrgrFGl
O+FMydkVAyS65KVQ36uMUmwPzUF3DA/Tio0sKhsgWKNFFYhEkkIVl/TtBNS6Wd6FM+cjWLXgmiJ6
hWX7CbSHs/2MatvvbJI7jShHU4RmUAXuWMa/13zxSE8IDqq+pC6dIyBRTBPxLJkaUx1tUKUtlwGq
87pKnuZ9eSyHe/teNdWEi9YNuP7KjxpeGP/1mfDvQP3g8dO6A+LexMlgJY0Qe3Hjzoe6yzvPhmXx
AI/9pOb62wHEfaD87gcHuKLA0audTsTcJnyrqwSbuIoGdbmU5/ZKJcYveg/sOeTkTmj01NxEFC1/
8QwVZ3omLrlO0Vzc1Zc499u85jxJ1/bxJcXWOO4x0isXrf1OTs4N7TS3bLNpLO22cxFEgGXHsQ85
PYssoz7uRZ363yNwrQwZcW13skF4wE8AhbG6mZAAOP4sI8txIQevw76FvQqzt++Xilsdu+A+tWQ+
4RfG3s105IrJA438+k20EGvZPbw1EIlEke0kVyAu5OGm6F1lrp4mQmDUi59pRU8pWWBtsG9/f8Lt
Wub/cGFL/TgQ0Wj8Z7PB2eR0X28k1XFETmioxZPMmhmvc3Dx5zZsM4w8U6Mbne33nVPLFFbt3VcZ
yiWBfbNt49LV0QDd5v0ffcOh4KcF6Ss6JQAHeUrulS6euFsdn2h54OTov89I4LWNY9+Md+7k4O4A
mSoD1wTDSfgQKpsgcvtPHzAHFguPVZNYmRXeZEUKNAscfsDEefp5pN9WZdayANeBw12Y//yyEZPY
X2fw1iylWHDhJ2iANBhBdOzwbMY64KDyIWjZVsUqiKqSlHfBYMdU4YX9mjlzYXp5sbqMJ8QJT2Cp
EMbUzw0nxUvS/7R32+C3tny/WxTW8XyeVjtYNZMEgn/EuUJCSu+28YuvBBrcD2v6N1wcJIJDljS4
YrdpgI+GU/wYNJItUe6r8Zx74jeotx9fyCmYP9sLxyWTmxx8IhftwfejvF+jDHNuo0avdeLtYzSe
KZSNomD+FINDCqiOtKE+pD8Gg4V1j/gjZDRuYbpbxGEDGGaoMN05EOJj2N6BbxA+J6emoLS/ageu
WknmrJGwAPyQxkostBHw63rjRxhi2pS9QfBqt0UucRWaFA6fvoP4921VwAI7hIZY1Y2SHBQFSxUX
+2TVk2qg0jUhzrdd/R8pgVlSeFZfDn/aUYqMsZz/y+j25TDbBUyMXo5eoGRkKflh8BdKz3w4a7ar
RLcAueTAwlbOfRNmQ+gCxusRTkfUzkz0S5DiGt2ZxA1iNhbJ9agasq685JR3u6htLi5Y+xVZlJeG
hN5hQVufw6Fy7cMc+d6Ur9hfXMkfXRXZWHfz6L2LB2UFrxnnRDr067N1OtN6WDOxZ0mAoU1PNHn8
cEyjRjS7OWd7cNKwDSCfBxp2utpyef4Ov0k15IZUqX4vtuL9bsDqrSkKrxq4ITkT4gml3hH8E7c+
KkSpx0CQEBa37qWOdV6DKMWT4XL2QocH6lkWGpcZxvBpuHvLUZe8/cUsoUe7Hx1I2xGj5tpdP5Rn
upuGm8IKWCOXzkJtFi01jnMdAwjzhaEx/YzY48zCElq4Z8ISMeTnJtrYdPL//ACGQuLf+MKhC2p2
DxG/uJRMWCNlwtII/FAhG7rKrZ6vqP/msIbzlL6+QBwwX9E+4/VMGAh3HCglF2A22zlp6aof0Fwv
cuH50wuUq8uUvqKhXKMmcjn85tUd9y1+86wiOPC13uUujet6OXDDXgbURpRj/qohY3cZ+1ZeQyxn
oD1Dj73SBykcgDVqxH7L/K4lhuxRPcAfrJ9kUcoXmOGNKECgYkpKaobCuCrXel+KVirsy/0eRsIu
1jplq7xvf1rh2Fx+uyxXzstcWuSEqgtKtcvPOLuT6aePXe0Jz44UuENchLBHRDkIKvJOOqsU1LQR
tVrF6eu05cFV1Mc6QE24Ddv5/1Z1cjJSVMi+5TiBI9Oa1OKPPRrSPG2fiSHjKtq1248FssLSis/4
4c8lgAPLrHHIgUjHDcFgNnP7WDvrzMZNFO6It0vj3M7uKjFqqSgI3Ia2wTiCZYyY8OQsA/GMuHaQ
QeIbcd/ukghm2+qOGGOWDsAqNhxgFqS7Bp9P1mtTUh78pSCrjPOA1E63ZX7e9pJLxAKan9UbAMGy
hQlXgljqTlgoiNDpsyTiq/qeV089RGChqmJuAb92VASaqgVF2cl6l21xF2gsuo8oRO86Ar8x0qlQ
m5ORcfzfGuArWm9ynYx6j0oof1Ij+hGjprUtgEq55mwbmhNTPuwGry32rr5e/JeP3uryekIDYkw8
+93KcStK1CdytARzMwdn3dVC2jPwmTZzBzSEuE0UMMWvr82U6+MEsH4Y9X1cxL5yuaneKtMjuSAB
Y0Z1BKR8weuNw46HSw+Oum8SMrJZGVxLLXci+cMRM2KWrv7N8YW+XYW+QdOq+nwaqZ6gouWopOhk
GRT/GkqEiTML4HMNmzg8d8mkH38aCSmrPgUJr7dQl+GcOHHWQLRNzwlxWqIbigpMcdurTiorjTmr
EWtjBxWBmxbsKguopopHI6RY4B1FUcQVUt9B3B/rOZEgPZqAXlEKT+3u7G2Xqu0xrc4u0Ovr4mLA
lZKs+1fSnIXiOlwT8mUkzqBSTkhKw+yTZvokdP1rca7Uyyf4GJi8MoMTuBHnqFttbddOUwujO/um
V4RLfCpTbGH1P361wgELyjuOY4vHiXwWzL+MPQcCx5L2SIoARRgQ1kAg3o6xKvlNDBorZDYDtWVX
/zCojEW3ard9ZCLsBa1k/mIkRAxDtkVZaERwdA04LfgISjM/rmIvUaLtkZAmV1Rvfo07IDrLTqt5
Jr//U7fHoOS2srRyuXstVhP6liocEOBAZmybQ/buzZzZo3z7IHjHnVltkrjs3WrOHDEXqzYyy49i
fWuM0pvQdjwaSKhSOJHPs6nPved3+J6ZASY52SDTU50FTLPk+Kglj+DjN9xHn5C9lQOld095TslN
oCJUTmYWgrWkJyKa04R+B6zN3b17OnRby5wv4o1FKL01GcadTl2s7HPc5uBYv43v+3Csupx8I8MS
Saf3cqMjinOWO4ICHtlgNT/i0FBa1kYNct7eyRa7qSycm3MXwjYpkWe4HqJ//hbNOyCB0naHsHrj
CJZo2wiCF4OOqR3fGoM+0f+z1AYXBEgSDB7HGPkXeebyEBSzsgm/Y1PwnTnLotbKMH173eduKLNL
zWR1/RYSm0JfaIF0qDfWzBGbZo+QGp8U/jiFZRCI8/pWZm8eNqYELTUZnjpJwrFcYe2Ermk4cVZe
hJr8uwB4PSwgDzjEPb82dDPGGXHRWPNWcztVcTprsuXEHPcgksNRhBNB+SNfmNqiW4tL0YEygFf0
Os9D+TWQ7Bc0mWF23LYzd9MKmTokD9hzaU0ndMaWer0A2LWlIH9VqDN1sBH779YxiyGsowOYrRBB
PeEsiv5Mbs294N1bMhpxE9NurH8mpbeZjGcLpv6eW35H4QBvCzJvjbBNe0Xz1KLgl/yWbS6pt8ZV
tD1ShmfF1COfDm7fJ/t5tImj2xxl713g28KfyQ6Ss5uKAr1iFPkCQUquraEfIM44PBLO2cu8bcMV
/TBfCQBKs99rAROmnkkBnttBi2vimf8qBDUEyvCrgZOY9IidnzNWFo19kUOXNDLcxl7MmE8CseJ0
OZQaQPo/8FekjjsFEib4u3lJURSHHQp9XIRzEE2N+72eUGPNCinBTtejt1J2762UirAoD9kjRIve
vfwXO2QkjX/1DDbmIQ/58YwYJNdQnCcQX3oIuWLVsh4JA9bDN6vr2m+U/1OGvQb5ZuByONtOEYmh
YeAoBKxlDRhhtkyWcApvuh2bRE+nJfIMZcZJdouczecySwOU8P8Mo3XWdfiu38iNGoJfqJGs005J
OWEH/UeU0DiaicEJyE71Dc7etHDg3C2ZSworS166+HvZYEJfbbVEhnz9o5BGRLYoZr6SYU3SQfYB
kr7YCNvQ8hzuthnuox+9fErUsxWjiMmq03zAeVM8cHOm4k/5Ehv6WCJxECIkc6NN9yr6PS9y5/lJ
VviqPzKXNCqXArvfBYKQZNh2A75YddPabnCzEsSkMtYq0KUAo0+mxUq/vsZ5U0ILJ0ibJkWH1F9O
WrkcCTczG0DEC0Q1RHSha2A/qIOUXZwCY9RYZreUHkWcIy/NcEJ0077gdQCnavz4hvg6Jn0rw8eR
NABTSbv0U+qKbhJ3XMC0S4sadMj+6cU8VO1Y0RrBwEDCBtUfTEIRrh6a88iSfFpIyGjq9jEQm80N
Jsc8UXW2uKHi2KLQ7g83fYgnoVnXQJSlTe4QdSWLTAJ6+F5BwTg0JjSnRXLivGjC2p70sfUPvTxG
ar7yrFMINoAMAffTMiO0pCGOqQCHUoJPjt5EdSKvB4JlKothgXWxaMjbfm7N0gxPyGaa2i1Sa7eg
BJC/wn96AtnPO6Ar/W0g13j8utdSfBSJKs+Qh0v2kOU9iU7d/OLGTmlzwgLNwurHOjzKEmtKATdr
gMF3+GA96NG+Ap4oWFZsCE7KYOEemSxwd01S1YD7TH4x7gDMeNxxxWzpsODYN7SoQgOVW7sv74CF
ircLyLsO3du99toV0mQ4TNF3qeGvG5z1UZANvw8U0+lHuWeVdKDb3c3ZlDKaqUtoG35LkQpNohdr
x9W8i1ONqotYghvvaOQ+/kdlw98DU+r1jbfEtXU9HXjdVyfInqC4sYJQs3UjX1HXtDhU5cpbx1TO
yoVRCUu7EhG7ls1dlJfLaPliTrM89l+/LzOXwpxYEtsupcWf68Wd1YYChr6trpn5Pa678SfjsCWb
U7hZKM7E1QrzqYDB467jyJ3vBlXhB/Hf1RTe7LVNVX19STNCkCZd05MGB//metzxdxRsTZhcybdo
dQDwwMpR7zbjfs96EbQ/mdAxRu3j3/RE5zpLc/dMsSzE8HsK6qwqJoU6q0UzMcG1kPQbaIT1YuoA
7fV+g/aazkpoSbk2Dq7JTs51DBZbJrlB0huSbTBoJmuuLA+VVTwh7uyqwVtgfmIxsrlF15yVm7uF
xg1uaU2w5SEtESYrAfnBL/IAnkBWcPv2YD2i8SexY3Truk4wfFR1mbmwExgPEbtLl9TlE9ukORwM
athTd/i9LouE342ca/24/KG+HTJ5FhibuN6meb0FFi+Bj6ftgIrTSClXBYt9Bw9S9k5pqqZrcDB1
Ed+4tYuIt1pN/11wURZBXSmOBlSV2QpkAQb9vWBDC6AwAI9YZCVWhXYw3VXtAeN6+xXerqoGXVbf
Axy3ztnuQ2BxfaLrgUgH6njJKKngJv+QrQbDAB1HPGvwJjb5vVlpeV2NG6JkFSjrLa3CG+GhjkpA
AKNIWnnE99KCv5pY1UYvMfwMVavTSpEGhpcOjOEDmlblAnWF2TiAfNUR05VUj1RgsHJ9/PLtLVbG
ZFKUb7oGw4yC/T0M+o+pM0tO0jFjUI+Mgoqu7LueiDHVVbfuOR6IMk7CtewtojYDmNK7VMikng6g
DVuY7H5AHNGxhLBQW57Wm86VTb/jg2y/vKL12pHCKjm2/JGSlE7hKT9cEob9PiBMf4wENAZ7mrZ1
PdMyd/IX0Ipn6jAV3BgjQcoGWxqBQTY+adhD08063BHrQsu02bgbIpjzonD8gC+AmDgGbHmUNYrz
189NKJ2YfeFmpU6mfwk7iaQuqyAdE+Ban/7mUqqntaT5K4MTDOK6Tbvn9xbSnDfNpkWUyPde+Xbu
SGJfCQ6vnTqFP42j6FvrAt0TuVJf6e3SGsvdl7wUYkJVNS3AMDTeFYgyP3IhUtPbH5NFcMa0isTs
mB3/yWWJxYOHzorQATlRstwhw9njkK9lG8jYxBhlMUW9Pc650XolSqZbDgAThUNvgdTStJEu7Z87
zQeJi4yyQup0SwNwBIdBrATzKJTMlqxC6AcUNas84hePsX17VDryfkstsfA4fVHG2muZUcCpMsSY
dOQ0mtImA6xOy2bcFx4YDfIiaJJ8zzMFIJiTeva7kIyz0yDwOsbzQpnOuj1O8QnfLycIutKC9LJ7
qD3b2qkrSd1o8uQ7iphXG+MS+gMaempNmQLJroXoUm8mQweZf/0jpKmRxPqYly481VEFob5ji75A
iEAwS8s3KddI5pm/maKqXvoVN8b8SJ78ZwjrMKCZVKOPinLtk2ZoMYg8574fHh3zsFbbKWL95bFi
x0C/GXaE4WwXHxGS3qUdYFF+yt2DO9lNC58nGDOP3KNFe9k21RnnAeX2z2qFNpEreSaiu+MXpXr/
Xnn49e3vWmQY3NPiSItkliRWHZo1gm/7+OJ+B2hi4INU0L5XZomdIMnKy6qLzbKRDeXl6wcFK+qC
oR9WwE1QM+67O5v00Ngg+fDh4PH0oNyj60PQ8Yrw86nvJuFgVgC8HWlIJKr/tKVPZfI5F8PpC1/z
7aAHb9BJ0s2pt/u8rB5xGZeGO3zy9euPNFZpeM4wkdTYddcNiRgAR0nbXtKVmY++hZNyW03+Egcw
AbgeEE9FR0fLkpzv1A/j4LqdxIAsL4DeItitVrZkAm/UTsoAn6N3wh5h2jkAjsxsu1knRs3gAOAf
4q0v492d0cIycLa8M4Umhc87q99jZ1FOVwyLBm9i388KXjxzuvUJMszRCUe849UWfK5K4MXCDkAa
6eggjWsFHzvRwGNQmPqUwMx28o8Undd35pbGsnwA1JeDukF6Hff+oy4ImMdMoV/+aVzAPzeQP4lb
kTq9Qfif7PgMnoD2t1pU3lm4eT4xzjVh/q2b+vtm4Ap9xHPx/A4YPIkSgbFJ6+Zg7FytWkHAsU9Z
+gL0o83gcowLJ3veBg+uD2hbfvYEgDkHb0QPzkenB+akjd/tcfEq293n+b3UET8Wq9EWGfR70dYq
EfVSCuoXbzle4ntavSzmumAn5cfhPnapLqHAXOrhvdENjZxA+rah/3qDVJolUMOMQgGjBTEQm82S
2XZw6M7wWQTl/AYpavkRNfuQiUW6Oln3OStpttS5ybShNDU2jBez5UuwaU9QHCWroJuj2a0HHUqw
rKsjoPQa9uNOAEc5IRnC+/et/3ayHhXq3BKQNQAgWdFj4GERfugWl2TyiJzfOGWGrG0nwIiFOTue
PBdh0Umpjgane7IpqIjYeMGR1fJI9SfQrrx7ii1Xmf8Icd78UGuUOfpETVpIPUJ8/Io/FfxGdPb0
vSzK0dO0SA9QcaartHWuRLqxmQha/vohE91Arkeq6LbeaEJ4dnKmsJCHzxruG2Y+bYNYX2Oau+2X
xYCr0RqQUcHm47qRSsjlw+Z0d+2y5gI00DvLNBGD0QR6tUTsSpgBsfCyba8YUNDWO5Wab45NJeA+
EMXIJTZp026LXL5zXyvbOlYfR6Dm8zaJKVRKZfyF5lgN0Iu5fRbjOebyHACXLOFCVgoQFibFwv4l
XAz7LXhkxR7s0aWW3AmJBfyBiOBZDN/0W81Tyz+GVBmG/wSIZLApUpBRAot6ebXmBmWepoorKr+j
qstK0Ksdy3fPG4Qx6RxZ+eYZFNtWiSSi4QBU3iuI44CwPpT/l/1EFO/TmmWCxMNhOuIrcX3ZxNYp
GaTpHersaJBw9BGtGnr/JSAuR+32mV0HyMmSTe1sXhWww+eQibHknjmiGWwTYErJG42pxUMNRoBr
ZCPEz441y9JQ7p3455jT/wU5nw4ofHXyCqAC2B2iRikrzq7KhFml/O6uhiE7PLQ7qk4C9dP8qqhJ
9wnukh55qmfGzX4YOSujTedolRK84b6R0eNXF6id8TjXRWzII8ncYvIVw5r23t17k/Jf1rrw20kT
rvzdLX1EB4xy7oFuCotO2bQYSnRtIIDR7RSDt2sQFX7cyr4OQ3OWJx92WsJffXN1+8XCI2hetYXO
zKWk1KUt4dTLgKf6DqC2+smytdQ+OrtEf8S0M8OA09ZR7+qKvDN/ZkBl9l9R9TNUCK6aoB29nY6h
2LO0qIuizNl4EJNuTb0O17xBssnqgWBPNYqYuk7oDiwjH1aTOASPUQXJls3q9Mn+m18pMycj0dBB
IkGp95jrBWsp++3fiIsnFmxPwtSigRgVvkGoYh9QHK9KxNqjs16oH8oOWxWoHjmo1+DsFelfaQ4y
H1BK6YKC2dIH+hz1NrOn++WCgh3Ie9Nh4xq9cyvG0jmrSV43GodSzx9+gItE//IXd3bO8UkIcjxl
cTUkzc+Jhz12OoL6VKqk7sIqtA+9zucyInoLNq/Cs0rIZdwtTWiXkoMgsOBTzUW5AQnGB3hU6nH0
6F5C+RkwY2pqoB/yiwlwcZscLpwzBf4cM3vO/TUyNfnV3sqdS+/ne9fgaWyB75/gF5bNvAOo3QuM
3R66NSHy9laRV9Uqy09rS1MuBVfQttEb/cGRbcGkDIyUmX+sTgqm8jSywyVaaIqNanfQP7VpfBQ9
WMXzdlOSmZXHYxNp4kUMPApynPWE3Djl3fH34FvWQEQMqzcGZdXOylKOFa17I2+04ArRRa2T2+OG
qz+rtKvlSyvNagvCBbX9kbpyvVx1n/3zpllFse9aM8n+tUQQPGxFp7VaT/I8huePW31LGcqGhVGU
Mj4FFRsypAjzAS56j6kdOVm8LzcRxLu5fE5Ir5CC0sVrVCdybmd7oyFJ8Q0ZHXKbPIfZAhNz9Hlh
lIG2IphMufGB1fk+FCdk/p0yY70tza8eJQwX+7KM6YwDXTd+PGUV/aldbcEz+3PZz6bDI8o2vZUI
YefHpJUQ811x3tCynTdhPasgOHGCtNc0+3kEZGkC4sIUNg8wNgV0xbYIiENYJ1VdWv/CQ2aOUphi
8416HaumJMtbMEEZcEipa3RqVr9zAYa7vAW7czWdOkvobEb3h+0HxIK27rnJii0SCZgxiEcpgbSF
xO9PMMXg1Tg4aCLLy3gXN06PDJSzZawUjjLGpPmN9xNrYF3JLyhqhJFFDr6lHQnBmvNpnEo0PFWc
Ah8P30wSnEA4bbUeh+qbdS1GK4AdYxH+lP/gmyHBpO5lfjj1sRzVkpv4qbOYmqtF0wpBPd7tBSJO
m7Xyk3WSOJ6PWecgqFXX43Ri28KMw4WJh0Yq3Vvun9DDbwff0nCxenlJ6CFfw55XF3xQ5EHNpdei
9nU5dJFmw6Ed/M9bZ5XZkJxBL/TtZPdLmX92jM+Bp8/nQSlJ1no7aN8OTqmWu179jTB+eFFRfkNk
LFGlXmYHpXFzOr9B1QPELE1VxIEouWyOpGQUk2qyi8cx8AoNUg+kvFlvjyZl7AvU4zOv933Je7RB
83f5SiMTbG8gUE7jNMN397WuWg+d1rF9xRq8gFhw4lJbS5VFapijPV1gG74MXnbh+TpLYUmk/w54
hjkxgS+LonDZ2+MT5LFZs+qVWSVrxtq83yPb7lfWCUO4cMRtMtFNX+lIgQ+11OTovebMKUogDxxs
5cV/W15SfwIebTukI3IC9xPNKBygCv88Dk+iBqWqSpYYn3ZV6T8Sc9JwzkdcfJv45gIH54P+DpH4
Ro8Z1Ck+M7t8F5jma1p5oz7EdV17dTUbq1DDoBNlveDOPFk9o+KGLqeomvRlYC9qL53t3XFaj2uP
EPHAw74hR9NS+rmgmSvtuqz40cRN4Z9Fa5SZgsLl57XT7DeicOFarCcxzGfB18UXEAaJGlilgIDr
ALDobOnUKRK2DZi3kLQLbULf8WMNahGdLzsrNxTNzvAg3s9iSNg3RSS+xOvsNkuUPrWVVl5ZUJRd
CSQvRXk8tuv0AAE/1i1YHlvUrN32cJ0kzI4CbYu+F1X8/hPX6ZeE0AaQFo5ylwzSRb4gUbSHyClP
1ecxRj95CfZ7vSpTjxCdDBylgKhcyPSTXHcyiTefUMZui0PmkCiyihy0mlafGGeUoks0tOFmEJ6w
Gx50vcDotNEtcF4W2WI/RdEPqyAPWsmX0PfTXw2LhCT9hS97Q78Yr/zhdyqgwtp+WvnoAmRXVPvj
Aq1hWnuxPcpwPkKpU9Is7YkjcTeDJHz8OUQnL70gnaweZhr6+xo4uu5u9dsQE3nP/uVvikAWqCto
m1XDpMOZM0UCrFEX5jqudGLGgSWCk1unAm4mFINpJ6od5lQMbQtGL9koDcuF5hc0xKQQakxPSYpZ
RLEkssUi6KNeQd5qWJ7FYcJDlq5wUNMA5aCxBFQX3SJ2ELXBq0EX40YV4K6llU7hGG6imrjCMH+I
JJm7TJftDiEJ0pvkogs86AvKzcQsZAvMAInCOuvDlIrqY5BvkfyXmH2aslYKoR+LL2jKpQUpVQjo
peX7xUhe1P0Fbij/08fKe94YnDL+eRvbyw35lS015BSeL49XNiTUQG4WL1+tD1V2Yib0So/1xah9
9axcUrxMN69uewFf89IHoifJ/0lMzsePHBVRoOZvWQpYuPHOV/L8Ec5vwixYG8gyymiXehAGMAnh
QGCdzF1hb4UT/uB7X0hyV+IfQvqzrRdP4F0OyfkWvA0qNDWF6cLq3Vr9U4LEunzrbJIWJlJc7eUE
1+H0h1xXfOjgET22qXGhjHhKgNaUlwxPoDLxQVFLcEZVUc4S3NoTlonI7k/CNV6AInSOGx96zaQK
t/PeSszmDa0WscC6PQhrLhauU1/CpXpnOP6/6eHtTieGvaaoYSebg0/PNvAvJh27JXrzKnqtla/M
tDVThAD+3qeHL+O99sVTnvzb1jz+LzEv2EBZsbTHciDRNCzjBXuAHvUni4SRnY3JVR8RD/R5krVQ
wdvLtpARlUjAFxftBC5QQZDJig3wSsF+O82RVlb/Li+MrZME9DRqsvAR3Kqcj/v8hwPxQTRavzuy
G0JfpeTGpB7Kig03rGTL+D5jyp2ZnxYDRr7Mz5y5FGoWcep3ky5jb0ZyqALDyuOzxU9UaYmKd2s0
rA4jgdpsLpoI5h8yHJWygdr8ELZOOTi28rEP5NJMDg4uUACNpHEU9X8I0jifibqH2eZT0QwFlv60
J1amizFi+nlQYs7ahyO3G7M61av1JxPRXD5C25hYTz2Dpd6sVVUJnS/b9jf1pP49yxtcxuV0lJKD
S46rYZZ1rm5UV7xlTqmbrVItyhfzGrz9YRnkRiZIhHdkecGPTPdC2NcgdQFIarVw5ny+ZvgE8OYi
kbqGSTg/LoIdldLbYMXu8mW2Br7csa6KsAumY+GXvPAbARQH0LWeLcVHkFPl1+1MchHJiedOGhof
hEcMWzKQun3ea6hnHR1tFal88m3l2XVLSLwtmI/rnic82gCLF4M3XM0bcsUZ9oDQXWXILbr38RsS
3g/zhhc5azE1XQ9CmzVzKAO0Tkl/zY+wczeeP//OwsICpmg6Tw9jSoy9sIu+wu4RD9MlyYTxhWZE
QVIhK7yWGbmiMsI2W9SJ8nQc+TOAo1lTF2zWznCbY5JyumQ/41udRcKnHEI39syqUYtqTH/CGB67
7HkRFQcEvqoQZ9GkDadvlZb7vqxf21t95TpFYmtkQpR+P6resawek9T5eV4fp1TyX4K7NR+j7UBX
QDgzBE5altjF6xgKA6u3OgAhQ556zt66tzXgoMckZjyu8U9sU4X3medVV7AR8G/TJKIOEB8FzO92
092HwnHNISavqYcrjHtrzsFRMhbrT1I5u8H2Wn4LIKfk4VrNRdliOFdbOVR5IFeE9cSS+TlSJ76h
nvQ1swxjljVgS8gipt1wA6GZCeHPE2fRU+t02IUVXh4pdGW/8x78ac4kx8440khUhtUDtyj+t31t
qxn3wFQRfy27HytNejb6SnR7Xxr1ik9WzYebUJAZuYnYOhiIQvAb02f34wcReVjOcLAQiQsjRnWK
XZspJ9mkNwpgRQzTrOBpm5vDktMEf3fIZdxZyRf5Ym9b9sky7yvdxQbMZSuQsxGQ01t3+UouxYYc
NmrOmW4NVvqeFoAgLuG39LzCub87iHfPKhXMo3rXV5/3hF5/ivnOSb7QFI1a7ewkMiEk9AG0/PVq
KaAyfphnT7clttekyBncPfnigk76rZBUgQigLbk5gwt+WI2uwAVjMMPmjWV/DjHF/sJ3zDDxtQUT
8dxusr0lK7Cxnioa9YC4bOiMN1jw9B53K7Vx80JPT1Do8RBjM7XZcqGnJvd4vGUs6Zn6VTOJyjK0
nYiEQfQXMq2k3dISWtLA0LMeBxQBYDB7LF8zjtGs5pcFEh/nlJ0itL+FDPMHj34E26oj01kvOzwO
eDuqRUJrg5/U9ZmIqiG2q1dZYP27R9NlMDrQ/iPr0pPUBakHdFZMQba9yY3zUmyDWVVADDiIxtt1
Mb5ImRRDsiV0yyIpjLpNNZoCcNWWVSVFAIvPgE5FGfrAwyhYoymS9XEG9F9MyVWhfbm32/bslHNo
8cj3hmqaJPw/qvwZWMIuTqWvJD4bc1Lba1W/EfA+y1q/HMAh8iJwZC0Mo/zRh3GoYbfw+iBUFAlp
VRoAL2YlnOhOeM95rE2Vxm79pJAahkqOq5s/wVunVG4T8l1xKMTkiadO2wXk0TT1B1guOWPh/hCV
pOpX+11hgZQQxbtWLG6fH9RnL7iCRbJrtDrjoXzGcs3I5XP77lNQyxFshpNfnbXyRQdMUUiHC8rE
HoyF2wzj/jD1GX+V4YEZn2B2IK2j61hAc2ZWvZCu1bVlmLDYR6f+RxQAbq/GVA6eJncVjFsKevTM
wEP0uyPlTjrlXPHr2UQ9hXau/in2upel2xmNj1eM440IfQpcOU+xBSnl3gY7ylyMa64n4J9qM4Tf
776m4hWR4IY8XoCYFH4p6W45+kqugulXPD24z3SUExpA4P9kjA9B/b5R+XDIGqU1083EaoJJidXt
+qk0Lr7v48gAvjcWOGK80FmEZsVCUNFstQtG8YNmilo+vo+7wB5wiLW5b6j70see9h9ZPlUYAEma
zTMJrkWhMcjbs79Nb0wtexwtnsbqfeFLIh2crs21iN2rZNBvt7aCq7gAcOnoGI6/KtzOoZL/TOR6
hicSZzJQZVhL0UhhkwQvwOVuBWLMkJ8OwfOxoINiz/cuMD0v8ibxkXkU4FrTIfsSeh2qY+9Fyo8E
RoS4BOgzhpMONH/WxGpxsitEMZD5tYacUVd6R+erJDe1sSJkrwsm4GmG1sccx44LsJBWxRjr2Zy9
mmY7oa2BB0Hsap5Ob12WfpKN076ltwhwwYyZadBh59WCCbIdADYm8fdLUn4bfuMz05g8CTeAhZKV
ePD3EGGszASKEim6IzBmaZj5efmjG7lcpFCZOqldpvYB7ol03pqlvRWd7inbH05wlX6KToOMfOAu
QObcScsQI7IahwcYoBHVJZW1YmrUU7XTxKPzA6uDs7vkh2scpGVG6jvcGiG13kviwdOx2AKIZz4P
oeAKJeYGF6ga/5KdVPApeSx6mJX8uu6e9j0b+EQOXhJHW1jyK5PDaXZyJg7clgzA3hTbH6FTSb+l
XRy1sfGbx6jt6Ai8I5k6y00kJqcmuDj1yW7vHeDGA9NHBYdRf62xA3WFLq8tEXw4RiLkbVXRH5+/
hhz+6cDuy7LjTlhMItKJ1a2J6D/GiI673yHLjq2ES+ITTOVeQuZ4Obw23fkjKKXE9Aptv3enZaM6
RNhzUwDtYwd1ZOMJkqoWlfwIVCH4ckN/xlk0hE20rDtVauk+isteVs948l0fzePnJ6qPjUdse7Eh
Prv6ya9YdZ5z5KrZ6tpMwzzlDmbuDYh9k6lxtEGlOdEKSM2artiVmmvwsT7qYdkvaTHEiYjIwNpv
EeuIVTSHx2dBUQJwxPLemyRog4DopuJ687HlfjOLyBfheZvb3pZ0M541u2w3lhCXLbanX4E/MdKI
GtGTkV4OHqpVR0iMue3tAAjOLQZwWD6J7kFq0Bp42FBHRg9Kx2TVOBx67qQ/WjDL4XK9o92jNxiy
wPALqYL8CipiwzSxBNoJITOZOjnRePjz0MPzI2eYW3v4J9GskYoSO166sGJXQ4SnbOe/nb1mY3Dh
egYQD0aMj8RAs6Q1zQece4p1e1lvuBvGL1ytlGFWUiVroM5tz54kQnqfWBOcC0pP9w1OX3OFga0P
xgBlWoZsbihE4uhgzAQIf1i++r+6kav4cYwDxhR+VKSdZ1ot1anlUStSMugH4sjqMhaYxa1Eafoq
tj2CKZ4iWcmsCYpK4qjbq3Fky4Y4GOf3ASu4kYy+CBLCzB6PS/Fwz+eeFc/M0en4NEeSWWCLV/BU
VRVKFCTENpl2xLKAbqPp9v7Sw164DaczRsmIJu1PiHpq2gnEtoGwm79mcvRetzcqTHRExuZJLUrq
B/ONcKTyJ26q4gVxbIwBL0Do/fHD7leVVVoa+gcHDTagZo8jd7vynO6n5XKKWj4xxnM3dgqUPqgc
/ggPqufcB99jG4nM62xDejE5r/ZZ1B3gvjtF9l2t1TzVorqmlHGcLuuRJmf2LOev4FWptZgpbO/b
2WVJ8jXhG1ifoWoAjcP1i4SbLHr+snOQMIoHoI6Y2uBAu7WtP2YQKUvu7YAUBlA3hIqZ3mYf4Dzb
ezKooNg23PlUDkyforyIY0qFj2CwGbQyC7ExMQt8iEBbuUhQeEdwBSYSfra5GWDqrDX0w+Yvbi+k
/a86DlvZUScQtd7nTiVLSOrSfNWTIk3pV8BFI/qpCMGyPDi06YtC604x7W7srXPWgHlQKfX8UU4u
OD4p5a73SOhi/hV2+tkPY3SfGOEsY4y1tzN0wiCVatjOhc+1zSNGpCTem28pcnxmovGbhmFJFvks
ps6c2jwdsPYUXjyUuNDJpyVnionv6bSBLSP008YIe1laed8NAq6k+iqRMxndvhB7xaoLscatPXZI
C7p3ncyx8636fGTa66iayrNIFBIlTEpTCRM1DHJ4HtpdscQACUEKhdQurghXOQYAqazKw9ckM5fg
4seOxXFEHZ2WJ6lEYLAEWW2BeSs+nKVHiNRzzCDIATg0mOTu3jl+RtIHtIlbKAfYftAzjYoanLP3
+fyaIsuOsxo0S0TzEvk5gTR8jsEJSriWiYx5MbIjFPxyTUwexVS4RJEiSXnEK8jufxxPBWiWOk2a
Zqx4OoI1EKVuW/uThPJ1kz+P9lW1YRTDXuYcv1oxm3V9zi7CUhtf/7RgKMWGrUkX2qER2Xr+fnnO
NfBHoYJQqZze/WT6eMaIfbYtmdqKN4rufi5aNMRsGwLwRtj9upIvrHLKNpqOiDy2czwFX8PpyXVe
RVH/u45IZTF94o8bTx+vEPelzypdDUcexrkfo1YYIxGM1O8MeZoV4j7jCPRsf+PyXPVCS0UAhW0f
0oyPPuapb6T548uxXFw1m+4vuYbgRVHREA38RBiwQO/WTWJ8AS23D/Rpz3TIBxGk+MyxRckmJJ/n
4qdazS/NJedNRzaRUtuowh9OLhdBek4z/iMH1gY9jvYagqQlZIcgzmLyT2tyMhacVTw9D4780Xz8
e2+2Ews2X8NZtL2Wm3SGo0pN3/vuk0xvRvhs85D05+/CucgXsxb94BGg6E3/BCllqvKzC9ADrnOP
AdCLV/BIEFr/c9A3k/CpPhL1gTFta3ZrX9X1e0aVO1fk9Ypk+4KQm3GOK1l4YfVdx/Ew5Y3190CP
aiK/wLYq64j4WrhjJi1xdfQB1wn1s7p0dZgXJX7c9sIYYGOTmy+D+1fFQzz2zTCx9E1AeZ64e6dN
2xkS2Kt7+IyqwIbNr7A0iyT9utQhqM9Us2k6JaPCNgFR/WmToBY9+ssxTqB0SwNThJ1TncC+YrXJ
Tu4nz9mBS4a1MjaPygR0HHFBb+OrXUfwl0svyHoTVP4Y2Oo53w+nWGLpLbbnTRXLMagYy6mmt1n7
SgTo8SJ2GVGWK2fTMxlFTPzXlTi+ake//hcPfOkQsPkqzFlASqQMD4GJU7QhMd+WG8czpyisIhpA
S3Gw1Svt7YHg7/WIb/Kd61W4WqVO4jwFgaGAgNhO4pCquv7MO1P3WDkVcyrJNowm/XBnCI95AW9t
pzVHvZVosmlSAQE1gx8VFG+kLXJN4OOMzJsyRQVxvze6JPcWTubQ3l8L+IO6YieTEdg43+3deScq
r1RfbOhfRcGsHx4pZENFKyBJriuwhgbUc1hOF5fy/Z/SEMUocZzLTcAIs7PXVdQTiLOdrfsIXlVv
j/p4WuU8q/mTvODKvH56jp0UgxyfaRIyHZiKZD7/Si2Wj7LJYib4mRctL7ofvLos+6GrcY0YEAf2
a5jzKTjqedH7CoKVspfB8xUW99WvaWqGgD/X7MDxCVv/mQl3+uVAU1sODValSGq2UDLgZxrjUg4A
ydnAl2mLyaHjh3HJcjA+IxaOxiX5ThaUa9AaJltPxv+lu6iQb+rBLEbxuzb7ZeJWsBcg2hAE/j9J
z0wHAIjT6h/XTazAR+ZHSO9zIC+e3Jx93Nhj0u9Hnfw2hsIPa3l8+Yych8Q0mAF3pZjnfIdvAyoS
L4IYqSC1VCev5oWnwnoIgQmzx95GwA1teRf62pTLMuvILtGdhCVt6a3VYfqP+HkmNqH6EnzBvpCj
EkG4vpL21fd00bJNxFbHLTbDto9YOi+Q34+d0atshfwyUHFIRKHMzfbxgaxQte/ycdypirStjAaG
AH7FNub8ypn7zqNiEW09ytv1Vncd9uF1lFR95VrSklvzqM6wUBIfjqyze/KU2ZenWlrp1gBPy1CF
Ef3rWbfkWVlq0g/y4u4rioqlRsZw+DdX6ZE62Jdg+3InwnS/uBnIZs8odxuEO3TJJXdrKFK0Gb7W
+WjjsoXjU+5mDyLFj/Z8ddR6Siv5k9hPLAU00uuCiDJovyaz+WbfG3R4pBhgueNcHwtgzBR6cYPd
PgisLglRfCmNRwY3ECmgNG5mLs2u8THgvjRWO/B4TrKaVLJ/ja6D/odfZ+uMqx44da0Dmj3OH65X
mUnjIve52pFlg8KWiWjacuNt6FEeGqa4OCh7QEiE0PMgBlKUZ+z0UdLnd484YlqhTImQrq+kvQjy
PComjovhUZqhrfLDf9szolnrQtQx8jDllNU+RMMsWCzOzqHxSsBJ1QoISEQko5DdVonzUwntcs2y
nW4KpnMviE8Iq16bDp49Su8cBD5uZjy7Jy8PmIp2M9qfjBAUJ7s7YKih5vag4kb3o7q/L3dODeor
Ob5IO8jp/+DV2RUuQ2AyE1oqgj6u6kFlXmaqlGlB/fEWqfGhSkhql/z5ncweUgk7rbv1kLxNlyDb
Y9BL1eke5jA4q2SjKCiySDV2sfXxwbCQD+ApxMxByY5J+qsvLcajwotaekS5Nr/juTbwDZH9t1bL
FBx7VnG7wSRlZ3YEyPRF0YWcfJeAJRa7ev8ch0mbvAGhvsD15O6366Ld1y1ZHg1z5UdGq/zbz9FN
IvgXeow9a9zMTAq/srYESA6e3NaMTG+WJ7liHUzaauEjojWoRWSPocuz4ZdDDzWWBOgHMnbmQn+B
VAkeYaqACiePYAF38geRo0QOGCXjebZ6XBRrUlugh2Y3YIlQp2dP7HWlQKQt/91b3VYoQ6HF0BLA
kjoHseGS7HexCXNFCGBwvnrGLsj89W14+SQS4ygW8nSNPlNGNuuVVQSXUDq1dE9DZ7SCXMYLfODW
Ibvu4t4KKdkrLhLd9eLXwa+/Bjd9CM7BiINbMSF26k2qBZJkOO3iZ5T9CSqxExh3T9s2pp/rj0AD
QHXL/b7lS/v9aj8Ijay1nkilzqMtjiIkn47gBMNd40CLX0LK537YRNHn/ypycdCGa/alTGb5mKIo
bGckq0y8gj9ZCbQTBcUlyWCky7hzzYcwe9hfbJbPgsU3vlfmnQR1LoYR9NjTELBgqULdM5r65T7o
SLAzk7tDo3qWEG5cv7XD7BZlVqyth5R/mX5h2SzJV1gWJ454kzDJ56jXl2Am55pb+Pj5IMycdgln
1P2wfufLsYlDIjfhb0kTSCeaRTC7dPzZz5no1dFUo+cSnCMLxbaYDsaax7gT4gNcHU54QWTUXrt6
peYqtIGXzt1Jyl4TEbc6Z1XmEIkKqrP3OeD0rCGemYW8KLFL/f+Rxo+rYm3PQk7HbAy+zP7ENbV/
8oqglN68Nx+WPsy9O01/GiBu2r441XdUtfOxDm+NfUBueywIsLCqAwoMrieh7EhmOflN8na9nbu1
g44EBFwlaitEwNSbljBRn0NqSyF1ZpB+ySaeZnMRsG0ZmoKFYo4LpC0oQznwX3HRopiaee0bGTgl
Cu6/US1P1Bnc6hxfX1BOXpX3vCI5njKbrW7c7nahttMDQuWkQY5N/6bOadXERVp2Wq1xxzalhiTG
0jmz9owRqnBlHuknehQSGy+JVmKGXClLwnqXMwjNjLd7kfjc1g1Xo7nAYH8FFUKyWlRJHZDj/jH8
U40fust3H1CVIKPE6ANxwRwHexYI48+f/CEdBOVWk4ikaXEFjRJhKXVotjVcr9SXLkb2JRMtgxAk
DmB3mG8E3H+xHGN0RuT2IABoh7wTNzCMM7vEfENCE1+ZEaxGS+BIe1m7LkO1FHexJMfKxUcB1nWK
fVjw5wOM9VzFzXbArB2zpqI/smi/tlg/X/6gxvb9tEv/ruBRLxNlw2mrXbyr2YmS13WFbO3/mftV
daunie3Ok3hhLbwLVT9U/uewqcjPQjBfD1wSTfspb4MYei7OMu3fnZ8hDVQIfIyuVFSvDUrKpS1O
u+/j0gn8j2aMNeyFYc8Qo9cRg469D/SamlUwSPaLGM5PD5HUEuXVuH4Bumqjv2xuSqSD6sUld5/h
GU5wSzZupvV7K4tr5PGEuA8H+yHugYKR1KOII0y9daYfM4ZH9eJdH2ZJ4XcfHLFqq8giqtnPX9Xd
ZAzh3/sguy1d52w4uj9h9NLWFYJe8ETsq3ogaH8UtPrngrjPoIxL/AzQgHBtiJApQnIvS3O06c34
6+Qp88Gnmg8PqJDLcxR7cgvDSriN4BjJbLNd9u9EOwgEvdSe26iSaFEqXBfB4fruQZaotyVOHJ/l
ESuJu4vcdwVJB4fVl+etS2TrUXuP+izTuqf/Zprzulxgl9T/dBRplB5+BuqdIxxGqAt1gMeMa8+4
3OzgWYYejpvbCryahUUMELpHSzxPHrLcNtBlRgEVi+VOVza+aYJxmw9ot4UtYZ+c/LVtgILrKYuN
w0Hpa1CZe71Ft8CWD8IvOplmxNfGPTxRmcCDFU9bgV00Hxb4H8MlklGU3t0FSaH7kYPZpZmqS5Nt
DCntaJggrouwuk5HAj5yedfH7bo0tEXfNVx6VlWZZ7UkY/lyj25ZJolQiUJ/gl1l9+zTUu5Hx6KA
fXo5IxJSv2p7gJV3b0U5fOsRrZTnDxAZLoWhZrd98m0bfKSkpmrxYRIS7qQzPwLZ+Ah0fvZtTEK5
V3wMN8OPyQbfl94+eCzTNYBOGo1A5x5do7wKfaYSsHcSyBBfV+1cngF24ntHY48MieIq3ufc1Tnh
p69Noa0sF7maa6aM3uZzxrohf5u9CZCjDe7aCX8LtMFYIZKysIO2ClbSTJsILelpIxqkXa2UCBPY
W9mS8GRnYuQfRAnKBe3eD185S1Dj2dMQk4acynXGftD1fbGJtiwBjuuDr9simi6MuplJM2qINZjE
NtZLsK5qb81Vt5IjroHMAGYviqXprilA22zERQFVuStgKa0ZhEouq9jCOP8TW8iCPyKiaTck/2uj
IElXRydHumftRKj2XFHj3aD6+35CrSkDgXCNrPKM4zYtOMebodQQFAdbqFyYOXBbbiy4GUvHWrna
dtyRYbS3ShbFIDX+UxowMksTWLmy/nz5bOkdCCZpRg5azDf//9KLJf5IXxJKIXc1/sKqCcN9QAWg
klEmLds4/aHBcDnQ+pkgzU3eqKdklxkBDTwJG2Q9eBQU32Zv+0fW/QG7SGRI/4uBJpDOunu8OQ0s
QjZo79VvsXkCcGowG5rxWIklCpkZkcKzrRXIkkrZLSQZQ5bDLCdXppyZeI2+TTK9+LJg5vF5/hw/
Ju8ajWq10rdlHimUQSO0mHKTc7hD4LvMDY+U+5XkxjEpaPbeert26Xq2BiD2rLe4os/uL2bTr4ke
eRhseTQL0K6O5GMg5vVU6YqWWG4J23bTCV63mO4GOQPhR1IxYNABd2WIofvcWWKwpOkpOyMjFzLk
rtq5MnztDIMdzt+De6x8btDf7blpQBFSgBjq959G+Nm03dINUMGg1hqhb3K1/0ALeuTWkV0SKc9J
rZjS8aorBj0UIdzRrYFI7Iw/VrlJT+JSZMhlX37k08W12RQIVACSpaI72nXdssPuonrPxx+EcCes
c6W7mZd6KnKZTUHUI8KeHnnHeOj+ajQuDk9/I/qUHlX4zfCY6Hf/GOJsFgncyE/0I2o6W7+hSNhV
d6870BavSPFrh6ncXxcpcbamSO+uTNHxalzjeu6kMuspPgdREaOwcAQR9rXC2iLcEWDfh5F+WAks
Dj6Ak0SAH5ZcFu5SHiv0f36s/Jsc+49GrrhHPSFtMoUGdbH6yj8NV1XNG3oI3Rz1mY4LBwzGiHtk
x9NXy0g6wxddGqeZRNKoKrkcIkvX5VaXmM47aFO4ovVruayqFOfrKf1QOSDsmgbFLJKfDITZOA4u
eTDkYSvhlOWAdAueSIG5z8+ncBjsZRM3hzYTg7qsNIc/PVH1pvHEfp9Liq1mHtLTmEZs1VSiG3fU
xauJ0DvLoqAPYrdJIAYZkvY9Yk8YrsT454wMvONg7yiORGK/hUv10pRHTyauDPDcDWaBwaPmNVDg
tYoJ+2metmiyGQcAWsRKmbkw1P6eHYWenjdjCpXaQ7/t5O1Ju7KEdfAoclMhx+yVbI9fqS4j5Z54
onXmVO5v0m/RlmDOuYYXrr+X9fRjpNavoj3ueBqG2755SwwwWhSw1QBUsbGc+FkUGl4j9HR6TXX/
52MsqEKFQUJc1p87gFvUwZWux1LrFrRCY0FqvtttiXf1DG+U0DacZY8Q40v8JWu7akTkFX5SmJf6
SnYUcl+7lT3eTbUVRoVi76pZSZcfQ1zDKrRF1yrAEBR9l59wYu70eRtbQ8HC0xaP6aog65QiDfWh
I8RAWf7fGe4SuooutPuVMdZOgdeJj0OUnJYKDkmU9K+YugPqi8qqcjHkMtxHtsGTCqP/G8F/eMKW
KWcfDUpmp1Z2mpG5CqJ+BHhqS6nhUp8QNjUcCQhh6L77/sXs0pyDNZD6rDOsZA1p8FwZPL5K3h14
tpBYFwUdvcecVjRloW4BBrHmE4cJL0yw6r4HDtgnhKd2nVXunXi3MuaX8qtyXZBJFWR5H5KIQULj
rjs6pPUnFaA1YjhTj+O7Y0t25HdYwVwXBqAaXEbAvQh87l6J9/upDf7zNpEEODiqVAOMyTCgCgRm
O1i74wIMnJmduaRiw1eIgifKFkePb7rhLmQuyPzonYxXSITW9Ye9p7FzLXEbAlPibo+Ze8w6tR0k
8+/FLr5zwNmas3AJ9n+jamURCWNqm3o9Bfx0ctV9Zrv5rqkck6XYMjQxOljEYaelxIFsurHuhJ9i
cFqZoqSzJc8Gi/+U2IdBbIYaYAK2iBwtMIivO3fjvfhazrSdp7NGIZiUNSTdJ6HPr0pjY3A1TwqB
neKkDSHVHUAo+BzQsb6C6UEELrzk4l0E5gDsLVFSnwVWno/GH7OcoXyC/Eji9ICYPhZ7jUzFOcwF
75Ehc3EyGd0KqYK04uoeAwSRcdJv/9nLDPtB0o6On+lIoQV9T+QzZK6y/JLELGxg7kILGAHqGsb1
UWhpfSBo7X+dPTJuXnW0SgCW0GyHbDkhKBzPD4wMhjzKvRcmteaFv3qbFqYnMExk+4WfUq1fSQY8
EcmLdbFJXkHM0XObTkbZ+CK4+kmOSZqwhtnqRCh279Me1YAVPyYZ6rDbF+DxEF9sbeQENssuonNc
a4AmC6vHofLj5RI8Cw5uoffNfiLYEsyLQCozHCYRppkThcH987ocRFxCkA0cmbSn6NKNuC62mjB/
iEpxQ9CzCdGxNbsID7a6fU3wnGSKyw7PRUqKtSB53En+opzVZUQ8YndupmxQkqSUqCwyZRsPfxGI
Tqx0l7qZsnFE/uNsd/qJ6eWk71QGPNJpjPzhPJGEgwodegZt8Y0e1msjqbUfgGRaYG+v06pFliT7
RdxY/CNgXTCiuXyfxu+XGdWA4DfxvplXvCbkMYWmDkbKx/PP0ckJkXJ7ZDwOfOd9IQm/74tvZegK
z3jIGQc+rmU2I/CjJyReTcCMyjuOsb0zQ+Un9jdyThsOcdMJOT78Vib6XXI7kEbI0WtDKuQfX9yk
4BwskRAaS9aQs9Hg19RglUP74W0cZTuON4SdDNJoGxRmm9mVJgBak9tf72+Auxv6aBoJe5Z+jYYf
EOZkYRnwKHuAzUh2kQPlUS2zLshS1xDoUy4+WksWodeRP2AEf4GcTnFFZwAktSnFOU7cGvU77BSV
GgCt7HnSZY3Dz2fJSFCapk+FgpEeXueSsIVS4Ldndwq7urI0DB+wnToFq/pn7AFx1fYtXegpDDsY
ggfLAwePx1amFJt/jvu9I5RH6rPqQTvVW617FyonL53dR+leTyx2TMUckpZn+hduaX1aVBzpAY3k
qc1apwH6Du8FmKajeiA415gcQdk00JgwppTrYN4nAsi9eVErFnFBH6ItaMcs2MZpLmzYNzJerDo8
RVH8C8G6FL68dhOvDuupvB+fODxt9HG4uEVjM7QqRd24naK/N+c6TZvCdHQc/GT6j9h2eG01ym8t
8J0rt6cLsHSPbyvH2pXyGaZ+4heSDgRT/gSqG/AXEFOQ58pnVLFFnGbGdavzwHALPHZvRXUSheps
Bm+ulqbP0FHXIu8+JeCk+zQZypjn3VnUeoYw/Z8oXjqtBiMEFslvyVgsb40A+uL2dqzRMoYb1NQn
dCzKBKj0gDG5FFMtTNMnIds84JAA/usJiuFLboK/CCztnXyEFIZpKu/eqX/UrLuNR8h9/K+Zjy2Q
hQdkzgTia7kfzK5s3sUT61+Cik8SzgNba71wU8xaFY8peddz0FFvO9WigsITcm7VjUB7HcI7l9a2
49if2eXxTpcvmAsuPfZtS5KfqL668uIgi1E6OFK8IP2voQmw6vyrosjIgGZerQ44ul7W3BMyXwtR
3sneIHW73/YzIqsYa4PP4qc33tkvRuP8d25OMQ81GFZvV+dPlQBFLIcgBEctN33dn/lhDvPpDb0n
o15TZYdS+Y1TRwzq1CSDVPUZto4KCOH7Z4LoXTuJxrYfM8eRYv8ccxksN3dUDaOWflqGaWDye/Jt
jCGe36kHwvXzKf1g9Ar1v1AulkCOWBiowz0JahPs4kIy4kPGx8ny5RxXKLosPIPPqpko4xq9gKOY
LC/HRiq8hwTUoM3h2dAqwqQg79eSnkIFwjoHhidn7VQqPRYxsJ9JplE30dELnuVB05MafZpwElIb
RxnDK3Ff81BByzcvGiHB/sw6KkON3EOsJDoQPihFPc4WuwArVPOaXPE193zgw5Mrj37TNWAs0Pdk
xYB7+vs1qh2GclIpTQprRMTpmUjtSBQXVj9msQ4nwvXsaAIRqQY6OaQXaEdMYNGrgYx1VbnUQ+ry
TvfNVMBsuFqvFv+p9yDQW5+2iSg0jcpGo1/54reBBg6jyTXhgI6/m3BDFI84dlxN9lI2N339ckeq
Ci/QwqVMrZVB7vnOC7ATqkp1PCS2iQrRvZvG1IC5/sERzsr2A1aCk0C7MzcEiPY/Pbc8srgxbmiz
4iEsIZcX2IG7ob+L/aFb2HK36Uv+3QuyZZC6IEPHXTzQxhHJGiZrI45KgdbsCyi61z6aL7dleRr1
6De9hAYiknapwVCsSBSQkUZ8+wy+w9isIFj7IdLvgc50geSzUaS7fqRMlUvS27QZbF9DoI45afE8
ogrf/KQxaaOlfXNefG6yZEuKToEJVMF3r/v9ebWee4+ljpP09GrrgOEeamstoduNN9bPBCvtcW58
eIvA4vnnBBybGglgKn1Ic1SFtCh2X0s2Y4NAB+Y1ZxQ4VktnRRTun1F9f+0iHd7vZtBt7p51wGQh
JhVo+OPsXnGdYbNl+bU6EozpXJ3LxuyxoMNZqGrxTegQDpzKuzSe3h97l9gRUU75gY4wN+ojMTDa
OR2J/KfMc0PPUifa1dOM//S9JN4wdEZMNjHTDgmOLfSpR2j8Q6VLi8uDqXHn6SYN7TRYXzzJjUYJ
Y/XM+WETGbq/Dkzz2sRcwMhCHq//vycC/HwZDz39UjTxEHn6YuMSFXFj6sduwFEqQjLmXI+6kcR/
15qt0ycXCqunwhVbbDZAU0jS3JYiBVdJwL1/NXHs7SXjYo+sSgDVCch3B8FkcoLQ6IQtelR3jZ9d
AR6T5LrjCiH6YyIKcWj8K9UZ6SWU0sqqxCHWcnnlT+KNUJdKLqdfbU2E4fD22GKzlHXIwV2TswS1
lZRewnpwY6Dp/JkupxG0vweh0Fxi9Hj2pzcUHhXubSi89OFxRSCBZ8qti9aBKF0DXx4APfuZKan2
g1WsCTYtLIV5nyjPffEi9qqxCR1p8AE+8D9qYopCpOe6z3S4mNAHGxlnmu633ubrZaLRaAPVZ4Pm
Yq+DuoROjXhAjeJDcBOi5pAuNxdYYfkX8DfZzBdI3xK0rFCXcTOD7qxn5GVzVKO2V/gpA6w6VQsz
AJzjZhQwXQ0ilue421N0zo7flTPEkk3W6F9po1AfJfl7f/2L0XN3mH1GRRx3jN0xW0clC3TAPI+D
lsgq90Qwqaj+7kp1FSgwHH16F310LvcNFsnq25OA8fsjJrqBE+2DTkDZ83xWTkDl73C69DZwNyld
tJGbaDRzBfHR2uoZ+rSv8y95xSd3nTWg0i4uOJdcr1wrbqa8QfEskURGgthYGHluoRqIEjPyM82f
rwNkV3Xd65uxiz+AsnsZvKFU2jGbzF3AArG0v5MNZ4DVFLloXxCzLt0za8AcikC/7Pc0+dsZVDiG
BCbWOrYzgP6MBQ/iXGNulXJ6d3hQZGWhxjZPMQFZhK0IeL067J+drMKqHbmIuNx5hzG04cf8n6Ff
zUDbsOSqK1J7Zr4jMg02u8tMyUMhQpR5jjTC51YO612tOmeFllJbFESRsrWlFXq6tqhCesDPH9G7
DAetCKM9zUGqWsi1jZtHiNaM09bW8q/Mybg4m1LpEiORJUQfZeS6hXWb/Sq57h+t7B/5Ae83hf2s
4NcpEg4ZDLHxJ5iYEMN/rlRKNyV6/24SGl3+ke12p+9SHn9Uuy2FWraJ9nQ5DsvPGCUt4pY60kvi
t3AAxXTNpY/ZHwOdTd7zPQ9cDKy01BZ9iDmWPKMW8MGLtqPCAEg3u+zo4ywgXcNBSqzpqUWvXrQX
CQ9zJAWaTNdMu3a5HavpCkzf8MFulW2zS2BTjQ0CON+kn2i8orKZK/VxkITNZtRrReL8KSTmg2fE
p3ZSGgX1Gm4G1EFH8a7+YDAdHJHGOrLZ4icyJh9sNzmDDRr4mjfCRlQBNCHSFJ0qmWbIOTAr5DfF
mIl8DLrSMbJWfZg07Zu8Nlr7dJI2ladBEsypJq8Gbs2vm7NM/Rpu6Y1ZXxNwU5Xpr1WTXNPLfo/D
ljqHvVqFZyMhilDb6U3tftsx+D8P8n08mc06dcuWYVcdm1nGCS7gnk++wLsM8VWyZR+n+SJt7Ytj
ZoepA6f3R/Qox7Ylcfy4TKkOuC5QZtRH4MxK1oVfUsXq6peH0lAXyic56shoSvgT69dNScTHJiuq
oLj5Vmm1dq9hdgrxJMJSsCMNnbCFP6/EeF0OL8GQ4KvOygHQqKWcZVb2cG9AadwQMRayfeZlLJnx
o1kBMGKG9PnT7ZLJny/HIOHvWQdSQGh36AtIJG/DJ/jBoMspjj0xRUlUoEdZqxbANZyYQKzSOaGq
86iVScc+o2Zjacv5C0NC7TXfdN6DPKCSg6aTpmjTt/kNKQ3I9Sh0d3bdEi6LEVW+H7zRURFXMc9R
b1AdFsIB81WwIWuOPHi4P2t/dv7mz7wk09EdcAHvUcKXMw5B2ll5hdiQBrdjYoF2s6m3rsBk5H/8
ujPEvWlDJPBhfRT100Ry/8gyKy+i0qx5QzvRYk5vKKA8w6+MOe3WQJE3X/NEJRngwAPxS8/KZzzP
J7C2I8yAXq6gJiGUNh04DeY3qqRpDNloIjcCBnblMVFYg9rwKXm42fU7Wu3AOk+vrWOyFDgZMU1Q
bbTA51HCswHfOD/+Gxnz5A8UxO0XArIPr25T6ELpMZ5Yz1sg5tP5tAVhznO+GB11r0RGjBAnd6e7
oYPmpVQBYDLAGsRvura+L8sfJBngy4/DgS+qr/10wzWkhf3perHa1WdZMrEx5HAAES0oRXiW+KgP
wy0oNzvnenFJuE31jC5JQM1Gx48t+cwYUNU4jvXTKFksTCwGkUu2FZvvQ6EjrNWs9Tqm7t98K53L
orrvdZjnGtzTpBJaU9QZWonvmqbqckNTHxlkxKQXGq5/WCuSmOvGz2UpUwTtQknFitlzLazKCYIo
zQdoceqKMUk+Wlm4bBKGty0T5R81va3VgefWbeDr1PqZ/pjIP3b7KFoGFRSXS1p1IYUb/qHwxKfI
e3oD4g3rYM9pjO6sxYEAqo0Lysym49/rExHXU12Mb1GMO/OL6LZ0reaBU3V/B2bP9aznJZ36cKW+
tq03xk+Tnb1qSTGR1qqiskFk2oWvpHYUQvORFqb03yShM4SpEePMzCF0+D6BDNJKMS8Ol+ZQd9Fl
Gggy5u5Zva2huoHr131nAw+vLumDe8USAbb16AV94SyNDsBzPNU3FnYxNaLsyxizcb5IyJf3fdUp
cn/02I2h1L8/gHw/o9oQl/H7fmzAvGX50FTD9wBJ9wf8fRKRK/en0D+o+d/oi/a0OnEcArs/aOer
/qSZ943oDkzC/t2H4Nvi5GYJ/KE2rJOGL21ECVQEB9xTnPJOyxuWIEVdpfXsRvW9rO8N0eamYXYh
Hu2BN9K5PUNgI5q56/5I57iXBvtyhVBsw5B5ThrAqvoNMHM/2MEKzlju0jVm8pqTGp7roUIBvW6u
D8iXNmWaYAhw0eUJKXLYIVrRyu96MVBxJohJ0zkuW/NRdzpyeA9uFI6F2GMfMnVODTIHQ2X5vm1+
UHDotnIMo0+KlRt9A5X9svoj2giEAYUNIwCfzRLa1BBVuLnJd7fr0pDiNbn9sF87e8NGjT+OCrX2
43GeYw4VWmTPbJMxi/N3bNNhT7ThZIazONjvUL96KZzNHqq3tdsrDMFOpQWsnXHz6ezVzzILsoEw
A2c61Q70Y3pGTUkyM+u7KMfFf7ZNgqO66PWi3xAq1ZRAxN/qOOMmduOdi3ObhAGBVhx9Bz1X9Z8L
e3TjrJFvjgevIfpeStxfRFs5PdS47V30KIwxvXFNdd7wN5+miMvKd0Ci76ZhGq2AADAHq18Mj7ti
M79T49GvYP41be4fy0TZFBP+3HxI+s1ol5HUnQwJ+xjGXRwkfdxwDZYrV4SwTeHHjLuhRtLHmgjI
8TkKDGz+XwY80t3xn0v6HmIlVUe19V6wRqLPFJiZXmsax/M7ynJjvHdy7PlB3OfXyLsIfKKhCHaa
rAADOfk8YmpteUa98dGKiP7Odq0U6T87k3E1goXTjB8s3rXWhYDD3sfMQDrTr3XgQ0tSZq7STP7y
bXvXtlrtU70R9gFPJZpPSLxWYNbenFiEHYjqTGteKHSlDwaqjnKuB+rN+Bm32rvH1hm0n1fPg+3N
OypdK5ScwCaYJXIglcwKeeU1sf6yIXgc5iO8zbLPUZBuM9iJGKwSB1bDdvzxkNzH3KjoKvw4EX8K
f+F0meVYbN/uJEss/AhakmDMOZmo0vMR6hxH5lA/zb+94p8U2G9wBh4MJ6YHPR2Vj6iyR7DuSoFP
Zbalz3HcsBe4lLpxeP+uYr5rH5Td/8LW528xyLiGwiyFLt66CafgBYisLQkpzvkf33ykBj36zjnq
9OIJMsWFyT49YcsYNlJc/2VxDXklz7Pag3J2AaLEu1LADUWXJoN+3yTRvIWAHTiEdU1NN7o/h4UW
LZtLDJzI46Z/BwvKuRNhwXUntBfhoOsNzNNxSDifh4zfOCr3jV7ztzKumNPNUHo/DhMIakR0XfzL
A2WZqEf8PvaxX4YfzIwhkamJQ0vX8+SfR1DSwOZy6vhArOVw73F8Kj8Baac4AkV6LCunX6b/vfvy
xGap4An7vVuaqG2uB7s9c4gSWEMqDceRvUGFnldtyopse7H+ui9smj6U502wZJ/DWy/J3qhrJBbl
XPO56UApt7RQa0vluL3xu8jPqqBYj6SO68/OYKSggMh2tK1J0Pvh2ZeXZchkwootBYhzYPFoSHvY
p9WzPfPfXwYSjuFTDzB6c/QkwqAbUcC9PsV3V0vIA5oyCc8PMFGniA61Cbhmg9OR/E6UDHLwdLvO
DPMbmLg4XnAgCtI1/3pefTle+1VWbID0MZCZ9DXAGm8Zxa2iDYOb2KD6hmDx3hUOuuYJNeXOTL6i
1UgpRHzkwrOZrAmfCWdyk7kW5Co2oVGrAtjP8tb7YTXD6lDiK6//jzuzvSc8cl5t5LtpAeD7PK4u
MDIudte0Mqbsj2dR9df1iUiYUpMPGS7tFPsvYv2lMAXz8oEaN0ldOQ1gqeNqcZnbjWosxXSKOCsW
QfPGadNq+OeM494kP/knHKV6v3OLvLBbXy+tUJhqBppYhTJTZweCpsBA5zhYCXcmEVdX1Z6i6tlh
GhfWpmb/lGKNKE42XVv8m9HKNxbH5vZTUGCw443pYHSFMB2vqZDREJdvz9UU6migzWO0sz7r5yWK
8wjOTG4tEzhDSX8giwxQwNDE9L9gH3xDKPVjOgb/DL82OoAynH+rpllqWQyJ9xALL5YAWGjJCRdY
U66TmimwUtwkHQpuRuUAashrS18lAN9W3vGQJw5QWA5OSwb2ykSlO89hZc3CIJ9uvgiuUizAI2/R
Mf81dJckmYva0vZioNIKThItjUGffp7788kqqBbaGYkkBs83pDgtmH4UUJreIWniMSdkpvR4uulX
OKUxWGlCDjqnU31Hfb24rh4t+gYRQYEddLXzQgIHlYgyCnCpo5RLdzrkvUSMTVT4zyCYtLLsC3UO
GCQDR1cGuf5TUMo7w8cwFv+Jq1HZGClg8GJJ17QfKcmA9X8iwTGvpSxrmp82Nkam2BMwQF0cViJg
HXEuwafwme9A1wd8yvLVnLPqfA7yRICbbe7Q+/21P7JnBy/APLcg6WbxAXeBLamWRc6AwSolMj8z
U/Ihmvu9MOz9eqt3PDNkpIwXmmDY8Syev2qh8TWoWW8EYeUfxl1O0ULL5AyvlHLJ+pPH8n3mS9SL
0SqNS0y4manKk3Gnwu4NE0vGm0ZhzDd4YM4gLPaqakuXfSzmZkDhnRJ7Vv+tPmyWv0+N2l+QmrEV
zfsYmnqb2jEf/5JcuSP1P2v2C0yVrKBNMa02z1TlNwNJwLl7hRP+czmOPTwRw4dlw7GKs1YwC2hs
FtnJ5NwV6+fkgWQQJ/2d+jVG8xpUXNKyIiUmjmbXfStcpSjcHq/52UdP72w1nJ5edISOoRqtISB1
PWPoz1DKh5f1Ewyaj3JJ7c9ufLdyorEU4NpMvw3SuLiQFJZa7yERK49DnxniIkAPw9qkrNspOUGt
2QYFcy9VbBR6i3cDGmMajov2dJ03oXeMAPVD75acnz/e4W/ihSsx7Kx4v+H+5FzarEPLj6dXO6CH
ie/9ONxzy38yTvMG0J651rl/SyqjOxlXIqHUQ6YfkTyzpSiBTx5CaBw4P/Edsn4Q+doY9KWNZUFO
40En8r1Ib8Lze6PaAK/7/prDx1aIL6tZa1mjCOEZZgfENrOadQhK8+YiJR3veG2/754RhN1YFvwu
1FOFt4hZHGlinwOn0R5RaLVIW+HwtEStnMqOcBYRmKNQJaRwCLJKamS9l1FoXAhambroVX9yrekn
GPyIqEep2OMjtkeVBD65SRTpL5yMNB/nmHof8OvGX3P5Svlk5SQcA6ndwNNNAVkuZntK2FZA8cSv
4bKaK7sr566F/JdRmZEVM+5rjyoiisJeJ+BmKt+AKB6Ld5Hq+qjAB1mLlZO3JdqaLVIkRlFA3XoA
J5pWL3K5Bfch6BDUA2qISMcud3Mu3Xdq3sNEs2lxjel/BodWJSIckPRVOC90o1D0jh9Kwk+fKDjB
aoyeQUKGFWsXUzDR2ZrGEBCdxNOkhc9DkOKQFbZLUVYXM1L4bJUz5AOaCfsj6Q2orAmreUJxgwX8
MKhODZ6UwFV7D9NxR3uII3URfi5w8jK6sJj9rJgaPZNZa/skK/cF186mVHeiEPddv0AkvORxf0Md
CiRw4Mw/7gn66CR+Z4wW17HPkcZNk2kKt3PzHEiNRwjwz5WRcrPrPOk+fK+GX/bWkEHIE6tmxOds
9wY6Ts3TJ2l83QQYWdjKMyVvx+UUBkqxqpxZnIjzIrLp00OCbBM1tlL4K7KEKM/wAokvybXTt2EU
49jQlSS6PBENYHwNfBSLTb5AqaPMOLBFWcdCHz4qCAajY2eOUG9+wOrPInsjDG9PILUFFjMOb82z
XLgs30jwvjN66U+YjDsiIRMXzwtLClrmSgfMlx0hqE70WfWzIfDA+E4Rcas3eVVChiMtNp0rMuCY
2prE7Cin3VlH9ARXbrK0e44OJX7Rcg2dSZfrdynh7/x64woRF0qbWyq0i89zyG84FdKxwsoiag90
e6r79dUFFDRPxw1rdHP5DHsjTJn4O78rhpy3mmERwx8xPx7CwKNS+NtalAAp+9SX7o3yJ44euPnb
6FjQVXqt+EKVbrAgfQkzq/uvlMJfN/Wrfpdc/kCciN/iw7pYWjlxKIu4XmkzPTl3n4k9fPjZG3vx
WDPh8ZoAPtiOVTSXQnm1Pf7h3taFLkaHcq9ymK5HiGoz4lhyL4f9AlOGYKSKLAU6jWkJczLuhl57
iyPxINNjG4nJ2AAtYDHqYiiHm8k+1Y1s+lT8uWH4CP+LNYzwkvSYt1nVpP3lpPE5bgaNWun6Wr83
HUFM3/P+UtHWwzwCFq42Xtu7Jwk3M5pzOdy7fJ/aOBBrKwhDRlS2PJVD+f2cAqgosp/oB5tNqlVn
iQ61+tb7Y9inwaRj8qAIRWuqf68qjGoQLgRdTX+lvlfxpBs5qmYHxOzzDp+8jxfsn8/7yd5HhzHa
9TlLxOeVOBZMrA4RwT9b0Q9DYELWahsTaOzv44ubUpIFVP1uUsZwuesJ5Q3Bod4IZz5weIyWcVuc
mE0Pdm5QaFT20X8adwzZi85iySWm6DxIc2Ta0LrTZf9nZlFktySHIpsvGTJegq3EjGnWL/63rcnT
Ay5Bq8UriDF48yERM5uvQPzeM2Z6+wFfyfTfKWFjAwQ+KZUrggUHYuseaZ2X2mGepP9VIXD3pHXm
jdM0chA5W0nhPg8g1UkPTakXVVb9vhedG853knDijZclw95ucxEJUYxRku62xuFW+Navvcw3pNn8
+QGxjf3zNScxvtA+raajVYMUprfD3DEAj9zHlbQ+QWaF/sOv3Nr8YN+yw09ieWzqZcHKt5/uxd1h
yzjx2tLidFo+sR4NhGWogI5H2OU9avDhmIJKt4WzyXVEzpmuiywgXMR0v8B0bqc5X0I11lxUoChQ
gAFGyL+OMams8byK94AoAmR8f76Jdw/b2bcxJbefuXY4X+Eofj6PYOGy9077BfA5Yt1PYi9Od+td
SPYWakqZozWulQNuigDEPsRXsCQgqKQSZUfHG0A9GjkD93OyQpc+QtZLjw6mj6W2Gm2bDacrOvC/
5Huwosx+Bm4o2FjJCRm2qKq19bAZeFTFyqVZZpPZEkFe5EYQp/cISP+GBQPn6u7c/PEFLEzEVqyR
tz4G7M9rFkkyWA/RFkm7XBzm5zWM6zuqWrVURW+X2kRkL1smSl7DLbYU4I0lrRlNIv5bpqfChXjO
8FWNwpyzQIyFDoAwQKF39W2qabSNla6NV5k8ShfQdaotcjSnejZ8jRD7PGwSvQBCbIkAoYCma807
p78jNwgV7X36mSOe95eTZD4e9wLejev5i8+vcgZQLOeUtm5HkYyrh0hRR4G5QnpxTjadO6euw3dS
CXshXWcwulffZU/vl+bM/Q0OUItVKwYgPBPthLuhAtE7Dq0I1N50To8wGUNaSsdp/TfX9gGO1oBg
uaR1a7olscOWCxXyvswFdYxcmzpCIX43eWQP4vPMc2+uEsmStw5K1LgBWvJRP9N9fe15hNgl4EIB
/vXCjhg/9eP2sHl2dwFOmd6tk2Q/7I9lRxD4PldfgO5wbMaYx1ngp1MaTnx6Uz2MQK3VAAD+haOc
hZjvvWmLkfPrazgEXKOKNfIsqm7T3/asBAlVkrFLKX91W688qu8K0AEwXKCohe9r8Ytev9R4Nd2C
IpoqiVUKhgWMrTOTG3NpF1Yo1msWtC6Q5cY0WW4xuPBJ9/L0sbN+BREO1k6IlMFZdza6OYlTHW/R
RvMkp8KosGsfM3XI4tjYf3z+RBasg6ZcJI8VtJz8sVnwL4Cbzx7slXMe9OYrws4bdoLwxUEpqD4s
pQTUmgp7CGxQ7/Y/w/slsnTe9L34KdIiqADthE/dFhhzFHptvbdSMOriYkEGyfHABh4zNdQaGWIu
7LKBqziv+BUDhgYb5aTUnhD+2YsGOoivelaCCuQhJQaMarSYi1mozGv34kgyg08nHZ5AFnaekGUs
9ICfn7v7x7O4kyHXHOJ3wLfdl4HxJ+wLCTGqofm2qDm4XXPa69bmKVXrjwDLM1DVUZzsDtkw2Tpb
OCW0Yy6JC+8sfdkdBA9IloiwTL6+1hO0HyA5RVCEuzGohX0DzfPBkQgUIErNnA8cYIDM4gHkQZlY
Ir7+BtFuLW3uz5GlG7IfOL3tK4isIMB/6akzyQpL9Ya/+DoNOyHuWYgvExazC9ZHysxAVj0Knqvn
nvra08THSXuK1AX+Cooe83f45eUIss2HmPh4go6wZ1R5LY8oJzE4AbzmARLl9sGC7UY6UPa5vBqB
JtiE0uPOqq0PvE/RrsfhhIvNLkkWYc/RhTPNVMVEOC5XJoGtSsCLbb767tlx1nORYEcfJXYf3y8c
E982ZgNxxtwTUHGNd8+J3uBPxewjbfeUwjdD5tYe0AWdPBvpyZ/hSEjPnazurSE+7MVmu0BTXtYB
v/mLR5SqlNlaCfNzxTSjOrWTnsj67P2bsGEWWf84Iy8vGYmH/TSqx3jLKZYFnxGXBh/pm3yHhb9r
HBzGIp09feRBMifpfWEYV1dBNElKFh4a1bo6/Yy+X56xnRY+493sA10QdtmBsEeN+aOtMPjIdib6
gHhiwuUhBwDYLPlf6dDjzRrsmjvWEAWrqnTeHREKdLBkNS3fCSarNv5Slkm2nHTcowxsn9qZPaXP
3YZhUZ2BbKUQ6mqaFK3RKq+vUL8XZVZDb2eiDPdEaHAY418/g9XRcZG+JrMBsGprGcAqwjdjJ3ZH
Pdzz3Iq3OQLi1oZVsmgs0JKcTYOLsOQWeFfMCE0vC/eGonRNX1eeX7ZMFfQejHGAXTpnYaJ2Of6F
3/uS+zzocXHd4qOOu0K815n51x09zL5SnAzbzR/AeXfbPosSfoYC523FPQONmFstBQVDdMKnhcWq
/hW1MRUX5aKmoPmxpLBAGhf3eSSAaj0PKxWkU7pczhksulwuotmqTSEV7J2nqwsUCYul30DQLzNM
HCeh63LUwMXc5nZ1R4JACknsLCarFOBh7qntWfGzSE5AgWf+rx8lCWADoIEuBjKUL21EvtyhBYUj
pvUMdg7aK2SMCThSMe6EUqg5/5hJyUE8Ps9pGrZbEc2+V9+pV4cEwZOmcMTaKcvYS/x3Gs4bXiGL
J3LmN8nwqtkOEPvcPSHPu81jpa4sluFDi6C1WQL9qWSFOMDslV4ffMP8mkGSDnAEqe6pdxerTMXk
IYdI5pgkL5x/h4kh6QpzQD9YZ+ofScGZpKIFnAxO9iR1PLPu6DnMTU81x0oqz0xCmnPVxyzk9ESH
MU8iAWl+W29K/7l5d9aufZ6JkpSMXEtptvYlO4n8HnlMuR4uhyZ0Ha9ZSf31XyONPi7i/iAseEoF
qtb1HeW4FE+u1btV2QFpyB/ejPzxaTMAUIF4T92Liixf9YCE2NlT0OKEqUk61qe4JTuu4WU5ko/O
12w7H0DxJVIHZYH+/Nqcr33OOLqQBgWLEgLik31p59ZspBNLqXOybUlCp+Gv7gsksiGgDJZ/VOE/
2f6+ao9kw6fZKY/Ff7IVtmpgb3Kv8yO9862JRJ8HIm40SkB4APJcyXDSHP9WbfENy7ipjbaCsNy3
Qs7fjWYavzTmNNAucRLPnoqlkccZJxhkN+yBJmAUTM/aonDRMJC2xd6gL7u9rLTu0+kTHIZr5i3T
mTPYZOCBRGoByQyLpn5H3JUvfvMRai1Zu5he7SwLi258JTzkRBqnMIPKGesrCcHomYo4tgPzoGfL
s+8SFfFatVvGr4U33G4+GkmBN0MReEDY7M2NiundBhRMuCQuVDMwtA8GyjPFEkPtkLCBsp/4GLbP
YK9VhzQPQ40kMZDG06iM8wjciuRe8aj38Lplrb6E2dETxIx4niCAvUGWkOQ16myoErQRzGVfldR7
Kx8YRPJje0cn/8gMm5vwSOKUq7Lfv77VzUJrt8FSJBSJeqXAh7eqVGnm8sB7jbQ1x7xHqB0d8XFa
G3T9YPIIVs2uwOk4yrAcTQ1cx3KosMKgAon8sabP53pnCmWnNPec217wTrbjaWmJ98mWYLdM/KZt
T3CxjyghiQ0NtbJfRtZxDEiPqdHajoZlkWjEwRjqIc1QWLxc/CgOtQtnwib3iJCxfkRkXM+CDvbk
6KzgN8Hmqs4p+txvasgqZzbKaoea9C1512c24MJ1ezpR4STmWnz+KHdaKKNt6LWl180TsISXlP7y
EUolmCCeaD0F3M2cryF8HcA1TEozqzEOFPSM0Yt/IjwzHUx1pM50BOan7QJdIlf95caPT/db5ijS
3vchbKPkTpfTW5Kg2RfM/f1N3Dhvjvh6llJ5Kd+b5Zuh+e6Y4y54eLnxIycEnPiFA/gOLZce5XUI
k9gKJ3BZ/qJlxnC4HbJlf6LP8zBzP4TxUxEpLWU70xT/wPK9Da8OhzXASI8PZz6sxbOpFlX55cau
41YvtSLhAiiMX4f8G6DoPa3x2vZU0U5D4QINwN6KVTjFskWZygxaT6JbcbS47foKhuYE7ha96Tjq
oV08RdVHMVzGvhkxMHZyELXIDPEi8KQacYIYlfUaiXY7uE6oS9DU0LScFWnkUNiuQnvKyvm2+chu
AI+8GmxQS5r+UX8vPvQZIV7eTVXF+7HgdYp3NdVS20bEtF6/v2d2wHIO6kfPwJJf4yj3ApbnQVtU
3VHHOMY9aiH5OGcpQCSwvUXI3EJ9RSS1ODiqAxupYwGGDNsxskHoHcrSO2dSMpPi/0OiG7S0qrsh
pzn0Eo39KK8J5j1eloupt2/zkoODEFrCB747PHT2UEYul9Qk+bsNOSXlY6Zf7IwWjfRb2aPM3D5M
bKKv7EBSGqUJqZLzPeDPettEPzDutfTEAaRigTVnmBGb7rWShW96u/KSoPOwr/jUiu+zNHYfYfjl
y9mbQVJZ+X0miyldRiqwPu6LCqA6kIbrpEcNd5SHEjZaCjc4SyLJHXj1K3GHmtci3DDaumU0xoGd
nHhM7vwMdmqJDLPRs3J5j80/Hagz0TUqcDQsgdIzC3fif2CHSY2yf7qUVx4ytfUak25+WXERpuJ7
yhbQOscKyrNlylqGT9TYn6FxXLjcsFD0SDP80jwzgCQxGT6lr/aR7lrQ0dNrtBc9RTPGLrqI6Pbc
jjxxqNpr+TxWp8ZdD76qrNwj/XP7reOFOk2tpfiYVs0sMQIakEqwk8Wh/9yqGz57Q0NYyBhwCKh7
+TDwwKNccqvL1VFbZe9ZYR6z64juLCvOZDDsLev5VSU0IUBunvpnAS/1QMcJh9YQCMBffu7+vpyg
wGzPCncxrQhUg7dsS3ragvkR90vstOqDYV3Idwkx0nWk5nCWJbsMtdIxrdaIVm0FU0FwSWdvbrxT
tJXkkC+Bv3Xv6sQuU1z5n4MUeULYxZzHln0ZzKBl/Wx2oqy0Vu6S1E4zjEU0zTD8WVD6w574/ih9
7rnh4HIDFH5F7N3nMvxOQu6n49tS+DOEIO29iOKvFEBVIN5F4TdI26qmW1IqhuXoj/ATFrEJcp3n
cWQrA62zoWVVx+nlOxvHiPbrXO5RwPrkRhJEgmGsjlKOZ1a13JDx99Nj4o6Npg9jmEIOS0Q2iGf7
wZHMH/dendheh+L+NljDat0eKs9Z6c0DWajma/dM+c3CMYg9djjTzkL3vI7Zfalwox1dRt7vKVXx
mJEy7sVXEcnXwYrpxqCaQ4Ua2G2AGt57+/7tW5KSdfZ5sjUXVvf3C54XXXgfxbFZ3Os1ywFr4Nyi
pVOgNxaNgEimUIAbeiynA4SQOvzvHp/LRmdSo9A7z8KMaqTPVbHK22fl8lNiTW87Q/hdjPSh6Axh
ITTMcEAo6cdIlkj67SmnPPQQ9WlN0fsylcjDhyqswM2vlbCkBt9qDQXXRNxVpkdmUI3Bpz4VknX5
tCv3IYPeOIOivsUbv2zu6AUqvvgo5wLqy5aKKQsd+AQ068tdQWB3y0d5babmWFSLPrXmXDz6H8GP
u9GRH6fcuJYVCpA/lLCgT1sDBK2EA0CKnwBuSwqoEoY0m3lnyjrg60YFmDqWIep9BaQ6xVaYdcz0
O6MvHryezELMxPxkDjnO2iXcbuO3XupIn23KfFdd4F+TB3mu3XbeCPZYo6kY8w+o4geqVM/mrshZ
1R7DzXHdDagaJneonHsEkhFNR9ROasWksmEstEAGflWKfoxvJ1Nu4f1KuNZBhPa2ZuPWpU7e5l+l
C+4m8z8dF3HrVHuhEWOfr7kuZpS8Oazy3E7VKX8WONw7+eSMGFhy0HUl2bqKFWSbjKG8shXJApXI
4vpqfkyK4TfgE8CzzFGZbg00++do/Hr9towDKj9+I4skjwIHXyRlvs7y6oFoMmr9X8Pw5nQmICPe
n+d6DkK6+52WKT7K2MugvMKoZySDxpKUV/fdUNT7pvZaR2xZy1CfMVr6rExD2ZAreDgfSNodZwiL
aGc/ISL7BJTmEVaxfLKtsKYaYU1THp9s+SYrbunGkClMv0CgAt1y7k+cEA95QZ9SevxVB+VNzXqy
YbK+VmpBIHjzk+M6dMmQorCnAbiR0mQB/mkueUoB9yehHN8Wi+kjk1c4tWWqFyelhEn0iYTzrICK
6IP6iWQpOT+t/HCVuyBh1FdhC1/k9q/rR39ICnTlcjtte6yPqQjUzJHM6SmenJj1tgvzrKyAD9CH
gjfni9pPS/XBTcpDjhp1Ean+qtfXAb5lNkSLyCxe4OrMvZiAmXGQcvIlatIkBuWQu95ey0W/cyga
boTjDsS19Kc3XmQ7MIxDkPiC77QGfOb1883Og3XAm0Cr8Rf5GyUHj+kP0LhRqD6HmU7fhtgDXc8B
suhPDVUc8NbSsJ2Dv9Ll+egCxSV2B+1wGqpJhLGfbgyDNhS2h2GDn56+IS5jTyNpfrsFEiokGMgO
JYMwRDa7PU8dhiNbPoDJ3kRQkKc7ncs7zxEqqHBp6a0raR7sQHyzFTT4drveaRIsJS574TSUJVRK
4F5ck5GuNHShwvEhPPAvmhk7YuPD70ENfI2h7DT8S1uO3DQ92B66UqpNlbIxCRaYRLel9AOse9OP
wyHMBf+1BVecidk0Qtd5trWQqCmwHZ0UJAuzD/CWsVPzxA/hCBgK02v+Yw640nztA6SDL0Tb6mux
7LyMNGDllHozQ9XJplRL7jFpXJ1FtRa/NK96XC4aiqQbi/GRgaQUeqRmfl2JBabdx+wEhPX0/drX
V1XHwdcPvWagmU3eHljKvEt42ica31TNy13tYsXj5yt/0RNMrp3x4YjM5Ih1F0vm4wnOtqlWzHyp
SRxV5M5UBooSA9c+ez+iNHCL9g+GTiTee+A92eTqRfT/Bkijr7aeGYaz3RPmj4hZOGcAC+lAEEsg
iAkyGWzkpSs2Ti8vA3kGwL+ZQrvdovxWo1bubjnTzGyNI6oV4f6ct0iZxV7dZKTzIi8VQpszq+wC
TXtlUmfgrRuQLToVuat7r3OBPCAVDrx5dPqhvKOKwAJhLYEXONS7mELEtu7QcWVekv58jGH+kXem
sKJPrYvi6cPY6LEljc6Wy6/nbpFOsLBoPYLx06jHmUycB4o6Zdj6KEJdUAcNjpwHkWMrzNMs+XDa
u766eC+o3aaGB5GTUnRsFGtj0D/owNq8Ivg65gHGG72xh8g7Qjpih2Qeps+U+qUx+Qvi1TOUcvML
VbOmRRHfUS/CUtzQwTfUtESQ9rdt1nIj6SNoBjKc9beStZrq6pUXO6wbRhzXx4FhYpVKP5GeRX3y
lIvNYBQSnI1UjuPtLmx1YtNebh/MJaN7j1BzsW5dVF20ueruqWfb6bKvylBOCcgHTm0ZJMwDypPR
ny2Pov1EWDW/xVWgu6gGgoAfWVA8+d0XO4XPAQMm/bgSxi10ti/SvFrWUBy6IB3X+DLucAGjv/CZ
7XD0cQ42Mh66wcOtQ9BJBsruegc/vRgqZotghlvdyvxGA/Ntpt3lxa31yIdvtRmkSjg3xfOUY0oo
3A2Trk162JUfDp9U8ny9GUBoiTxIKqKom+zAn9dMtvHzMbKvn5QgDQM2C0pdcyHFEEeuXqQ/h/qB
m7khxuvfE3sjXFcVxwpTFkFVK72yq4jJ7cvJdJ+ndMLhQOPsRF54RBI8Rg/ICzXBCig6+GtLz54Q
57W+6g7X04Rp3PbUhZ1ze+r9fTKidT8TYxvsBKSVQUAC0hpwth6fQ/hmaVlCm7lQ2qBCNPQg1D8G
s3RINVFNYAAYMG5XSD1Izc1/Dqbx61MZFU9MEe7tU4G7vOAZBk/BpPO9F61yk5+7euF03N2LG/px
me3sRDoBiZImeo0nGZ3I9Ib9gTw/16IUhcz0Prb3pQyPUwwfhNNV05KKnK6Kl3/oaX2tUO5EjOkZ
t2+s2lSvrHyastHtT1/NelYv0mja5Yw95tNSb1oShAAGbvOIR2q+I0RLZIPf00piK9Kk2b9UYrFj
vKnyojYkTXjHSnQB3wbzAxXFTRubY72NriRGOjt9vSgECDoMvnD1vrDlVLNFOje/iVobiGDx9rws
HAzxBewYc/BdwW9LlsV3v0ljVgDW3MjiVM8dypNnUtwbqnQV7cDMYUm+fJUS0QMHU+8z5WU0qgGe
4JSA7REwmma8N1zirvorvWiUU0Nfq3HZLk6PUcioPLdmLwPwkTAxad9QBwfGmbRrRYNnhEHiqhkX
0jZ4TmXnEWKG2IpOHG3IJMuxM7TjI1+uzNy/oP97hgV/5icaFLr9Qv/22gSfDJrmpAn1sZo/caH/
3UHEqgCYfFlQL87cNe4F2Rwn0C5bLLeDVW3BxrHRzQotik+4xOCvgVD5jubg0J9irRE0TffOc6cg
Fc5AXl7qaSmFeY6QDS/t44UUKvh8Lj3Kp5wJr/PCO2xo0YSWDCJdIYMJrzhr+3ci4s5j5TctOywY
LqatqI1tMpFzzHkDOLoqZtRcU+bIuPTS3lVv07L+N8FHV3/lZ3dwlbRCiDGNMUNWZncjJSwfBlo9
6h0RMSe1RrIpEbX+EJzRbQZ5B2K2hZ5kiHsrp0gIW3bdyV5yKPIgg+FeCvc2k7Y6MNI9Xo/nBd8F
aL2R6Ikl2IFsXlRU1CWUmdTt5vLtIEkZNjm8+BGF3//ycigJ7kP3WqXQjS8NWX/R3dLlwh7bb3Um
e5HS5q5DqX0F3/KxiQikN0Cj/xM2ycJfaaQhjDtij0w9hhFwbSr6JdfsAwMCxt8hd8esseKBGn2P
cxSshW+WYBdvNSJCKnMn3lqb5knqj6f+u6siyh51aFx+yZH8PLsXtDwXnDZfekvJwhttMXryx9CY
xyn8M4YfSKZ+oN2ZlnVDxyRm63WUIlsHgTBfvJ/AUAgBgAY+7e7wbJgDqknp7bHVrRCf8ArBXMnt
8MsCfM92QW8gKAIz2q/Q/kU+nnH5OQETrK+5cjNGMEuVDHs0L58/HETr5MaSwCqORBz+Ml6qJYay
uMPUD5YxDVSlNdNOZ64kCJyqlo1ZMCboCSGZ884/YlBXjYVT011K9FUPX2pJTsaQ+1hYO1tTXqti
hCKxYEs5MBSrc48qZG5ooxGln9df/v0Au/56590CCailwyLD8atcZLYjC/fWQEwKqyVuuHZ6+nIi
VhF7dCC8GNwut1HnUeXtSZSZCP8P+pbXAfKw4/MscDnRmh3NM+VKdV37wRNYbmgEQdeGtA4zGKQ+
iq9j5RtWQy3ozAtSc/PjW6uzZh55sciJsaQetcxWwZv7/Vw1udKv2BBkMreQiWqe59g7Ev/tZqwy
n8J31/OMPOu8i4g0Vk76IdKSaM48aOuxA1R/h7fL7w0Q42wKnDCxSjmFPexl7JTVZv9SqQsDA6r/
b+A72xFq2xXXTlNOi77WI1+NgACPpYUT/KcS3CSTIX/I9DOxyBrlvSGj1NoFGp7jwzk2W8oZdYkz
4e6LUiHmARbjSvnPajVjg6LpHQNOIpvrcgi9COHrn5iqFsAhqDBF8fDOFU8/f3EffMp0giw0aTRh
1JFs/luNdWTn+iWfAb/YluMcpzlQSZQIkmyA3sTwFHY8k25La15FYGamHg/hTzck+Me65+hivwCr
8/VVSQ5WPFsnSMWIGlm5GFRZAlpSVLVWqRuanZomrkywGQMFTgaznKbjIp/BUtXZPnjN9IsFTFKL
IkBdRCR5MN3UPzarkVSulQhiR5Rb+gn4VrCgVcduuNQSwnLuhQcIjxgFpQHhAZDrN8OUWAFrP97k
EtTpCOT+ZLbBy2ie91k28r0fKeeEHtEiqMm1mGEenQzGZOPzpFCWCquRMO2FGtkWrYrVTPl2CSPZ
zr3T/v7VhL/+0tv2e8vg4VYxZmSUFte9zrJIx9JcI/rUGGLVIbEPisKPEeYrHtYj8YVYZ6EL0rr4
L3uYTlDJKgvgDXn6yJSd3fK0psEfr+JHvTn7AoyO7PhP8JI3XfKSCoP328ySbW+CM9djGKkWTY9H
jN5Eirw+ndcmF+mIJI7LUA4vcTN1D6NqJa/8JqbP8l/M38CxMpC0YjJXa33/TnpUzk3inTxDAfEp
Lpft4/k0izaVAScwiQyLL7nZE3UAz54PahC0YJQ9pNPnf2z+gZc1Zk7R2H7ApXlmSVMEY/Q9iyiG
tSewXtAF6rieBQnc/yJpThhO+QQG4S6bZ7gfjZwBCUkiKEE2z+z0kkrPE0C7GnM60OsjjfKF4ViJ
AATh+zWnKkgrknIKrHI65WcwnRUuz2d5a6UUggbjykE1md4doaA/CbVivgZ+GPh2EwQO0zhlU393
KRYkOaqQQ5577X1PGmdbRGMi2kXUF6jIe7aL2oBZK4hQctUT3vw0/LfWvrKD/8VKv75Y7X4v61DM
3UITfxFKsIl8pqupAr0CK1UVGLc7GUzedv5n9UpN/aunAVP+aVu/VYQ0G0dp4PEcy3VcbXf12dCr
04D0x0k/8AfaB6uCYYeimbVBJ1AruZ4Q0Xw5wE20+I5JfNbg00gFIXswIex0x2/+F/YgqP8i7R0s
kYL3r0VWx7xnjfpscQjWX6V9VUOJYVMQuRsIJY4zk8us05zuedbAKyE58olXAs32PmTRX0ldCgJ2
hV1jPwKyS2A1PPsjvVO8McFOnJ7Oo+TD8qtpwvXMjNPnBKvJM8tivE6jFC92rOZYzMCIgBF+HRow
xP+ss00rWPLjwHznEKEiTYV82Fx06TQ9orHw1A41uUkiXBVmCZ7ahchf8GIkilyurVpoEV+I0ioW
T72C3xyUE+2XQ+y8rHSDmltHYH2PSGLtn2vBlV//Q9kF5NMRRTg8WQsbW0JYDSZi6QSy5P/dNQdg
/ZZIIr3B3kFtud9xcVmdJMWpc6n+BM2wEtC+KFf2YbcAfHf8VJFs1Cl9TRtZnPzSWoA9iJp3XuJJ
hhq3COdUAa39L/n7OdbJwbbaUm/xFqYE4b8Lilt9HyxPTcmBUgaFo5gitAmho2M6asrp5ThHt965
ZuT74nA/+qrX+nlbLooowupVKQEt+6TX3rOIvb2KwjLa7RFtjS/1f5inUw8t1i048a8/aRqYZ3Ts
hlaBsdCIPAWUHf1pOJNFPUtRJbJoqgCFPp2zjeQHStEgrWwFAXmFYwOnacqkSqKcTaZq6Fp0+fkY
3mmXapiQVQIfiCcLCz4kpRB+J1fCAxmfnF0Tr3+c4ozDkNy/79+XTmv969LVw0xoZd1oeB8TnT+d
9tzk/DzdzEU8+X4fxAbGn+xtk688EhRLmBpZlihzpxUk294Y7sC4BWZipcc72MblfZVA8fHaF3dj
TsX251uSvU39RnIe4vHOBEyu63MSBYMPPuDxKvr56KEdQ+8nbA1PMjyLJN/a1BnK2Ca1hZMsxK62
VZ3ieCarbyPkE1MYtE27UC3wSLZb1jA9tvWf1XV3czhfF4NnJTfyubCR6Tk9LMf02tokDa1sdCld
7nCf9vs0ak18s/uIEwwkMpQgVpB/453HbjL0HSP6dNvjRkz8ggNu8pOF3mTO/amQGghjmGEcCV3I
Y+6ibvPzxP48U1WMQE8OAqoZIFxN3e/a9nkKS0joQmy6IA9QsSymxjCCXT4Ww28npwfcEE5en0EA
v0qxzSV5+prbAS1unsQVYmS9a+1RvkQJ2lk3nIrdljTeGT37mBwjCWkOaF06o2TubACfWh6cbGwH
NAvrd0T06/fPf/PRLKC/3CYVS15zrOdC3efZXUx3kmNA73mlenHVSqJ89tLFb2cyZcA/AnnxdxBl
0IXKpBta+JoKbFdOllVmDDigRVwSxcmj29SuaS1WfB3o5d7q8gIAYjmlL7yCHBhfN9V63VkwTBkk
qOSbeV1TRs8SDGhF71wFmfYEtUux5pPs9GIo8YIcMqeSMdPRRuxP0PFejBky1nzEyJjK6K/fGx0S
vHs7n+yRSQzsvwarYReJQApNgaZCqVi49pz3tRyXBOESqMCu17/TtcgIAvebSMuxOnUORuoILoiF
N7SXMiyUhc00mS7MUy1rCxFi4DLPtJlCt8m+6HungzaogacG0L5Kd341pQZHpysVyvn+db6ikQS4
tloM0kBj3Mez762H6vy/8cECuIOtrvR+UMDT3r+OiTk1WELsrSp944Yz2AJ6NN6Hg+BNhEfHdZ2+
qSFX99zufofXiYzYBwjp5GSoA6xt1s4QY2AsWUUfuF2PHVko7Bei+7B3kLNbMlbKat9yyK8q4hk8
bIvidnDDpoRWtHqYS6YKNXpAHL3TLzJ1w9j7A+OVcClDMUY4NxW1XENAotRpjrrQo6QBhlXmYoFg
GKY84qGQwpBzcRvMTQQDtlq+4mWnILKgDQghb01WkHaxvVgB07U+RG3Njzzpy4wzVMjUAotC2uBy
RiJ4mgh4bNyBZc0UK2kn5OZSwzA8am3u6vYMCsLz7J3GWsgW4Rwidi3a36hFF0D1JszZ3hVFmqg5
HScsl0fJky23Txl+/CwCItZQZfU0NZMkHrKCXyfRBeobY+8MNBQyCfyldp5a8p+OAJ9DQi99P6aW
9ICWTb7+KUEZnDj+A8El2Knlb/WrR6jeoP50sLaKuMtjuNW3ty1gC6xAIOoEDH7wxC04XJ2lElL/
bTqRu+ZGNy17j1LW5K/xlEpMjJiGpa+NS1UkLfbCaXOQhTXDtHz1jlW9sZgw1vaXSS1yNdzXGRbu
lY1OKHXZvlSFQYhY7bTnCaiS8phMNPz3KreXjXh20C3OgxKYDZ7uSKMxXsUBhxcAsz38lCgSLVMS
yaCm5+L1bzlSdgo7wtJLQz6RFocQiWe7xU345Pu91puKryXt9HPmmp9+RwLCzUjOQ26Z6QV+iBcZ
zJbK+Y98kba/CXpOUTTLneBrpBdHMuKOFtYtGLmeimQzZ8OQY5oGKRjur5CrOFiQJdYImFlJZoZR
DesJEaAoiTXtoeU4GICfT6iyYHu7TBoqzJ66Ic7V4zoRbx7urGHYvPUMHFgWI+9TKq35iiW9szST
36oQra142KdGd1QRG6oP9W5LN+uCGMz2tMj54cyutqS1VKEXqrcvZBbTIkBFGF2aBWMiZlr6aEaL
2hixxEtwx/yYChg+RlQ2YCijHpaqSiXK7fxIoiM7MuM/j+ItzBYf9OV8yXB9NpWrjk59fm6SkkEv
ySHv8bfMEg3En2p0+PUt7hlOBop7A4TqoMFH3t6TUtwoatDAS2bG9LUbJuiaR9ThVvzAIGbwTQBB
w8JdYw8COEBYJuMwLKq2aOMF9DyJKmOP0jBCOMe6SJbwai4baErL1CDP6jhosvOnB7lSXGiGF8HA
7sjVPzjqguQ2RR6weNzwhQcUxtGl+sQn/D29csvW2oKRVGS0IyPCinHn9w87ijCpXbi1MPX9fm1B
WUYPZoBPRanfDSP25CsYZfy6ZkFNfWOFgOsDKu8xSkktaxntwo4gnWGy1sC92e2OPUI30/qpGStr
mS+rn1JbBf15ev09bevamSL9EjFOaLK700uZWYbh+SRcCHBU2KjtWNsC1dAlDrh2SuXFiXeFL/IR
9/QSmd5Q2POrP3IE+05P0Mim5E68zMuro5L/0bNX8axbEBq33CTSpZKOm+rk7C3vexO6iwbh/vjx
aPMUqufUgdZ3EYthl+puEXPOL1jNSGzaIRTXknly0D+jlB6+UWqIjnAeI+LgrC6kSQogm7aD2zkT
VUN3CBzjahFV6wYhZxvCId2Eh2XjZrofCGIEQ3w8pMPTtZo+RJ4qEowDhKKEo5HG8v6t3LSaYIfy
cHvnVYyHQMuHccXQseWH1uPxfZy5t5U889IB1ViH3rvsNwVBVz7V8MPjA9HtQOjOQ8W/byL/oCHw
h2KzksGbjEdJvtvAp5t1nfaKSoC/lYYuXED/6mGWqiqddPk3a3wKsZjDpDOBFyhNn8GaGUa9arDh
EYPWdJz3Kv0xLQmOnCr4iJpI4dAPTgi0CD2NqRsnOJ6G9mMhd5/pGCuaDgVaW3za6Ra0px2qjwHI
XyP+vhIVBv34rf2wRRVUt1MwOgJ+rKIw+kIfNqdfYI1pbNzpaSZxaxgQpiJQvcHTnh9VfX9Zxih6
j6mxSHJWwksYgCGaX21hA23XDHDV3pTTJJfvGb+FwzL+b/2oeYGpBXzhsnkGhyhwjE9hORBYpYTf
EnStny/YyAXU64CJIzLKFeb2GZrlIjuCwRjE6uAqdXYVbdm03xPIuR9BjujifAd8VRcyP3tpYs+/
/HNvpiT0HNIdQ7CwTEEmqNdho6UGBN27F4Jl8jYvK29ksD9RNZXO5S7gfy8P0F6QE+euhnKDua2o
fYhbqrNwgSFqNOUo0K2V3o5Mf70tdpqNCbRFHxtSXKUaqTRcIuHDDyMlnToaJqWcJyPJ7O+dhf9C
bOFPLkSZV9Xb8bJsHAWA8qhpFa2swqU4C+mybVuotP4/AKbpPr3AZaCgyzUGZbjsNQpdBm476tMA
li8WkFMpzzY8jjxN4DkTKiaU8DcSgZdJIrjwx9MDj8NwnXjs43FRAPTmmrtlpKLRwEq/Z0Rztlmr
sus0Dr9pFNbN4lV0I/ZiEvnWgdQUnecfJiStLEcQXRncRtqarDl8RIQCjoncWkl8hqyT5EsRKJCv
W1vNOl70stQrXok8bfjW9Ak1ohnB1TLyzBD3Q1GUlKDjb0YVfcAlfv+acoWvLETEcSailr+3Js/F
2bQM5AKChWF618YzI0YjCrLrAtaeHeilBKBCKlL+Edaryw1eHlUle8Lyfz292pZkjP86a5Ff3Xur
uzlzlYtoza6EuAdZfGtpB6zKivCJmIIRZmzX/12PCxTWkM1l1xhDwAUcAzr9G/cktJo4bnaunqNS
OTtgKLVN/SNqj0mwMgQVTBFNp6ubwFwecGau04p8YHdNeMkQYDSAtrwjSJbFetgxzGz/mKQ87Puh
Z86utKv83jAyg76m0PooLqDpZieBm0ImLYwvHnOr9Igsu+iZsmITNsy83oW6mNy/SZzi1bFgkSTp
au5LqjAsdhRoyEIkRz7HY2f0ULxuxBy75Rbi/KG/IhC7lBQiO/m+HQRBahWbfFxkIF0TJl4w5GjW
puBiRtV0v/+rPTE96Ht4JBZPMSFKgrDVyXH/fExb2SHi75gJnBrgWgk6Q4O8vH4vrZtw/KM0ASM/
jq+NaxIRZ0jmSvBb0YIWvlN6ZzGvogwibiX9Ww0bKvtUiDON4bca1BU5cpOefrNc4EfUbO15Rgxf
TALMHvvonnPDD4rxeLzUvDqhwPq/rhKVn8eRU2BKs4NxRQeft+akIm6yeGBTiP/HEI2+giTOxd5z
waC+TZjpYRuatJUrfX5CDw2kk7fW/wqfNJzqwTs3GWoa0ltc2FySGk+ma4zhWmv9mUh3Ja6q/l7a
x/rB8qEISktVMgPUl8RRQ8kCFaB5e8PiLSvNfB6AFcZBC1MKsa6CJBT2YudQZ0lhajBtKwIiq5zQ
/DrWa1fEx6m0wVeOAG2UXUIKRrfLRZQ/5Yn3aUh25BnPS2GX/abVaJK2+jZziX5o//lfxmJeJeRy
sw/tUKWfnR6S/NOQPuaj4JLE1G8LmRheIWWwv93aWOb0IvXdndsU5DjdpIBjS1XQksLCvPCL0dcp
Db2WDZQbACOHRRtfPClWYGslX8/l3KIJl2mOfJzJ3cF6IZU2IegDmTdYx9I7PI2lEl3l68BrNcAb
LDcfTle+rldGbQPqUBuWYMsdJnhyBGX9ApLYHWBUAnI3PRLDnHqmCIVFIe/huZ0naOl9oV1nMG43
HETkP25hr9gZGdBaxGLfdB/T/ZjUrl4Fz6wwAKSy9xMEtbOYKT+IJ6VHs3c/Qi4Mkld4e6lY3Qkf
wl7sgWPAwn7jxUEtpLLyvX7r/DQ1OjFJOAIZFXHG9frgBWUm2M0Wdu5StjTdYofgvdP2Eizrbbzf
UN68M0j4wTYgI6357NwjqZs3EIp4nY2FtYVte+WcW5nV3IOyi0L0oX3mefrUI5lcu2ucje7btKx2
70Zsl88C5ErZtCgW3f+/s3uMpsiyB3f9RJy+SldFYE4AH2TyoGJQNkOMbSzJVhNjJ9XCbmNnSTEU
alg2MJPAgOt4zxC+llyd2Y0Svk8YyRFZeygj+0iBCZDQJn0MeJEOj6PzCKlnKPgMwexGIU0PjGzG
Md5Fr4YS2RG405ssZgP5WNltA4dW2Z3nXaI8tXuxFlF96F3vbUwW1A/u0AaVS8yQzBMp3TdmLSw9
Y1DS58agujgXCdbPwiZy+QAlwyiO8YJ8jbMPwBdx2l/M9L3i43tTDozFh7TMd3ZRDl2nysyIKuFN
YlZ9ZjLrlIgGeg6+TNe9Ww2D3f4ybcpFbaRF4x//CKdHGvf40LW0CWdrSv7I9qfAazotG7G22s8w
/UIfECOYwgVNxCnE7QOXQTWwGNxzFg/0Ive+VjyJNi/e9+mKV3awYzPuTYNZtcY2ETDcC0FY3a5D
ZU1SJTmb4Og/tCfne7L4oux2YslByD3GUtgVgaIHK7iWQkKryH6bJX8XA7BlWYHOLOzuDpDfHMnP
zuLB6i5t6EXzFgRXk/DNW9TQtl4qn+TwAMiZWNYBbHoNKcLNLgJcM/smayKzKLvUFOYoc9G+aThK
HDDZIRXQczb6MV4BDAOZFNz0mYRP6DS4vFhZav0zUcMBJpBqwlsRXoN3NheXPymZKqSGi+rgW1X1
EJWTcbeQVAv+5bVh1Rjn4OQZxCB6nrxHhZcKdTLnjG8K7au6IaOtn3pX1BKII8bqk3Wf/lle/FLB
hlzkOz9tdAAyFaZBCKWpF+RAzBAerA1BaJlNiAGbe47YK1FFJC1g2H/cpg1Vf0G1JVM8zmfc+WJB
bCGe2FwSqzM/IZ7DZereCJtHs8epgXEFUEyeROBWwnMNttwSm2WSIicKdUfGx+Fy4Z/D2uuM0TPF
BFFRPyM4VvxptJxWSnPFz4/NUEn+I07FPioi7i1IcFhUKTsBBHbRr02VHBJIIT/+3Q0I+vsaoLoj
XNziZskiYybsuOexGeK/4jX1q88k2xyKVgdaCVoHqCzwdn9EWaDEb8k5xuxXkVcbMaK3V2Dod1HF
el5Zss2b98Vb91GuQ2ZPY+R0hYUidPJYsau4aUE+GFiES4bRHr8TVME/QmXJBVNSlyKn74sRcxAq
PYbYWTe5/aWFQs1YDMuIa2MRRxTeb2bCizTIj9YwT3wQDJCCbR8xm9ImAaT+MGQsi7Zr87YKuyu3
ECHsWA7O8w26s5zwlsgE207JmZysqtP8tEdI9kvES1pIsBK1cBQ3k+UN8r2Yi9hKkd+VhjJA8IC0
mGFf65LzO+KoDYwmiYFZXWPX2Kde52DRd5LhRwyFGNLhFbAhoVWULr1UadY418mxTQnlI7Rfu/c/
LnYdF+sEF4ta8nWzYNf65Ry+tuSrHCDUUHZuQfhU8+QwSl7h8fRWSUeIGTkuUwMY54q/+DSqkDD/
VjHgqTMOqc1cGC7GXbVwo52zgmURvWjWEVFfJM9gh8D4r6i3nS8Lr+UWidKKl98uyvtqm8CxwpCv
CAJqJYcnkrAbfoLRbUWBuwF8EVIGhMr6dF7CCrSEYqV5jpIH0j7wYLmwvuXfteE12KO9BdbvLaPu
kWaXmUWnvls4qeNsaDbjV/TNHAUpkhEc9B7cA9S9Q+oGVTtaYyfkGwPRXIgfX+dWwO/1STIlfgTQ
RW1u59Q3KmfCRCwYAzCwc3gTVmFmfHXKXQMcRscR5uldSXpZUx+GBk2IiLLxvwcqU/OrrWREIGEt
3Hpr8CdlfH7FWFy1m7ZVYFbwnmYLFozPacwBfXiovZfXEOH4zra5k2CDox1t+/cfNNcOvfKPwfRG
htF3KQma9tR0++VZjZzy1mMFlayPZ9gHq6vlp5K/I408TIg+1R4WuwBMPrZOhGqT6fENlxPoFnCy
1X1sVSOg/d4GpKW+q7xt0eprjRKhgCe0Y6G8GPy+exOPy+Z60j9vJxz0Z8aghuOT7AEbEQeiDYIr
foNdOJdt0alWdjf3x/BKrcVGeK/3IYShl1NgnkZoVNvoxh2VRg8Eb9eLsNZPvtga8pt5UTCTgdeT
yxqqsjcL10oHPR6FhjsJR2UBodY4c5AzAkqmpsfzI2jz9rGS+hZmDa9Om24P9TvSmS7Iol6hSiNP
bShNU5L0tBMHeAQAsDjqWMuQlSt2M092PvkVXNe2o6CAjzR4TZlXwsQeLbZkhDi54XZA6jM9thvT
p7PAw6aodmO8mW9CWQ/c6SUd70EP8IwYQ6wcj7qdMAevNM4tPcIiHb/vhK+hdcFXTevgdu9gxvO2
PX2jDeST+sVzQpr1IcsrzOeOHf88Zj9joeeyGcpDIYFZPKo854CKT80vhqCSw9tU4JcdneQbq/ux
kK0k4Vreh36RN2CVlRcbmi2zt5x+kRapimKtDvmM386lDdzDaQKC/ApVyt1uBYBsG/tZkz/PSfl5
KBwKuz+950jQYTFD8qludyxmdO8NDkB0+Y7C5kaF0iyV/hDTZHMwSlKWqTexe4gduJOkyFWWMYGb
CCUAVVZmy9ZhjL61fWsbg4Dz+JQPzDfkQT5hehwxd9V9WlnNZv0b7FqH1pQCBlvnWpO0sP9UNmMw
XHrIv6/3WPu7/qFAkRSLpJKa5/TGWyzsY4Uqw9q46/ruaxhoYo4iK4aoE2LDR9WmbUT3tBM8L8IW
UfzuWG2JNrQkunof7OImnCTXKQppoT0K4DZa6xkPPDOpraKn2eCU3KVvkRpKHRyYOouxixg4fJIM
dSf58GO+3RfuJaHBEF/q5uE7XRjAC382whliegyUgdbruHOzmtNgmWgq4fOCumq7NnWQkfLUZzdH
ciqzo8yY3mnS+KYqeCDVAW6l/w5njJ/u+yj1tpl09EiqxWmgvlzw763mD5IhArJ7X7IwQsstlqH5
N6Q5P4WLLUvdiOMHLNWjuxYJzGm5Q6rdkfXMYgnOHNgiroqZTbi1dX8/tsyZl7wEwkBs8qmX41FV
sz37ee2mtPK7NUSWKoySUIHXaSDO3Cc5W2ChNaOSOnJ8zadOI8yGwdhOKYxYjN/8RJVnZ0oDTVv8
ZNnT75jd4miW5o49UF3VGWclx/YRq/Qo8lMLIJUY6u5fqqJvT8ckQIFLl4uyfV+FXTuqUsxtMrOB
BpCAr2kAblzWcV98jKxXh5gmnlgWYLiLpo3UHavnrZCroNQZ582b1DJ6BuQ8QrLlEH3DhN0GQThf
yu9urEy92rlgWBQPNaqupZda4EfjtRqexraSN4SRf9s4xo9J6OYaYveTMRnEJ/SVkEi/AEbVkU5F
KlOVf69SYkE4rFatOq8zhIwZsEct9hV8I/Qc3wCtI7qaOHTNy2UlD0QmlV69hZ/C2qq4ALqtwjhj
fDyNd0zwAGmUF1GtLlgj6LoVbnfMyVPd1zDmS/1CmXyQ8418WIc1bmBgjMjXYb7+oraGJF9rmMYs
lApmE+PA3tQ+EI5tk/2R31ZkBQAmqjZqNwpBfd1wBVBR/m54WYZdnb0RRr98GjIGmJTXd/SjEQsL
YRqSX2AYQZ/xLFOFu5zzQxfzl59EAG23Sn9y/+zMRLcJdEjBRYSCzpQzqQHEN8MAPe16WTY8EdNg
aiYml3bOENDPZOxmG5MgDrk3adxGSoWGi1TDQshhKwnmep+tI1N87ew5p7gaEsI8pR2AExQJCwtV
B+V52U1uZAcK39FlaHLeQKz4hNlfgqq054YteOKSTedrkWHp03NokJx5nmhuS3Q2rkmRWFIYxPq+
BkSo+V7McU7ar9yOxKgZXpgpKscm4XRMyxgegxePlUSjIEoEaXat14M7HUwXp6t/zXpNeUPC+192
J/AH+d11aZHUMilgV3C0CBWIFy4EzILillLriN8k3il0TqGaiSA9rus3AtjgO7YZULXK+29YlUgO
HNbbmr6vQjeb+tSmyeUVyz5oq5wdIiEINY5N/4mB1RM0dlqJB+1WfzfKaOIyBWIOHQS7ZReltoo7
nKa5fb17qEMXrYj2WEfSIbIHNJIRO92VBLnlkzivPuZ0tpchODkpy8iOfHZNK5id4Ob1bKJAi5ju
XUpvSg2l+ekD/kyuY8q2TVv7YPLP89eRcCPf/n8n6VrHpwVgK4IR2mCYEQf1Old/jr8K9XBNyxxp
2xzImAZcr8Go4dXD06dpwP0Cn2TdTeiAukkWz8zwlU4/DgLemTFw+OANLnJdf6UK3lzVuBs+opqp
aSoi9o2O1g+gF+nG8lBCJd+SraXvSz42wMWXU22TfMWdUIwyN8x+j9EmYc6aWULIBxg5rka7jXbu
59Cu0T8RQYb/NeCMsgqTV1795qDXT6ePnf4jN2UbDEEAXTulvKJAlLD287OwFgciFOY8Lksswq/2
bq02FWL94RHRc5BxzUJv+neWAahCkujKVaatevXr3yY0GxJRqhT9UHNqTrzkdgf6hQCXSxce6iJ/
BdiXBlD0Mwc8WFXPO9ZKP/orPZSZbX3tSyqNhoqiewsl0FrXxemN8+IGL7n68JSRpZdediPF2Xbj
Bqw7NjsCk7Ay+yJiS/Qqn3aKL1t50tKyNue78S0Lii2b3MzlOKx563uUOXMwwW+t6Li0fMcH8YAg
b7LgtS2qNw6GEE5aNklk/Qcf39qksGZTTOsQIc3Lcvj2ooIVq41OWv51SmHwJ5GiJWowjkY6FpLn
bHh0g8dvORxGQLiZ5lkWVFC0n6h1XJPpJDpXzo35IHqEP+lx7yelTTXlZr6lTIFMbrDX9IwWKvII
DDeJE6AY/5f/Szui3G1tym+in5u0WrtSMHovQ/Spl+cnwyS1QsPYEaCesgPHZHRW0KwLU2aRp+pF
gAJQUqeTtqrtOO7aSYESI8w9rNKXcVbxh5HtWNj2to8CDt0sXqtJX8HVFlb2PodcOqtBCaJxOg8K
j9VwcCiVWTosRqUFZVpxlHazSC2JctfFxlqBdAIjPi735qgOAvkzQwnN9d6gln3CAPDVaRvU6IDz
GPL/1HsF+RSAsm13ZQto+6Jv/WqFYwQ99StzFiZyDuEhbRyoO1k57wAJJfvZGIQyEVl/Y/lljkvZ
hVp9m6vggaH5OuADnTEe/XrHjyj7VvXtAr9k/DR1dJ/tcy5h3s98L6+SmskXMUF0Kbp646mN2Ukn
kADcHF+vfOMg+vSdjnDpiQX8bm4+tdwRoO5oN0L1lcNEGToRBRVkErAQTGqZKd37naSdOhX2j4KS
xbX0hSgjYd7QA3+ft1EABOEbHXQsZcOGyLGy6seMZA44GPWtgBLEPskWD1lw5/gI1oW+DrfwaL/r
HTfdHSjy8DKfWFnmhRwYouSfIeWKnysieRW07Igrf+69+rh/4Sb2sROCy2fHuII9FIcfjyfx7gNv
zDcgCHqQJZZ0rfebjMOTfz8caXNxyWkO9zKXWtg5p+9mzBM02EvRtz17P63LWdvhaJavorgubqp6
r/bkBFKz1AWlZBvi3LdYKuliP1Z13BfRMxNdmY2ZQjo1QSurkbgwVDpg1tS5AGmBnqIHYs4gqUe/
a9OYx9jvlwu5B8yTVU7h+AsjzvEam4GhwO4MDWXxZubpwBMlQwlzqA4GfSlVIJMi5XuwEMEtuW4X
pv4Zrxa3bf7cwZoihlJNXiPZ1YQTmbDaXXU+eNXYhbPDPdJ3Br/zhR2waQ02ujC/T8Bb0btgeo8l
VO0LP/IvMaSyjpBkN/5cOe0E/RLIKQIePZOXWr3uIQF0LK/sz5Nh217E/0cj1tsNwN7Gym3RmIQU
JSS+6ZTje5G6tCs+CfGu6Jy3ePyZY7q425VBvEyL2j12pPm4f4NIAAT6ovkQbisl2erH5rYuvbKk
N1HSliJ4L+7saq2/FqiAgse8iWCz8TD45EMnhMvTrtBZ3B8m5XMzR+vTCveFdFFY5YzqAQ1MrsDf
TtuDXmJYx2n/RWlt4QDuSit1ZHh4PdbVlaLA7FtLg4fzieVZfJPav0Vw4p4P5bUTw//msUA3hOL2
PsNr0VAJ34a5uBAOMs8ZakkoBZjxtQta662sOqUFLSlwU9JHRcP/AO2LzNz/mdRQ5H7lpRxzzA2c
yImZ7C8J6pykO6l3NQLvIQq2AoG3B8mwBhnPQUWnj79zKHHSrQTkbfDd5o5WK0186K7Qd7Jfn6IP
KYNq/PkckkYDwd2xwQjJzyLNUwvKjj5UVAUYJ2hIJLVEJAzhLKXLo+Gwuq9Ok2NkdCWG9O2oMFxM
KJnPQQVB8JEyam00ASZlDI5+gwpG75LoMFSOaXYQNlIDnLz7sL7gDVqQGPn0z+hEFULLECobkpEt
ffbdqxb3VB9Hz4FY7MjfVn+J5IT/6fitJIKVLJZJ38o8ploXwtLQVsErGqYqSwxtA5JGGdPLAANW
2uqQTM1SKtXIO/jzAuCD7Wvv28dlgPIAtMGWVSYaWfvXf6jhyUFBUngnU7ZBaWAg6j0AGaGNkEJM
88ggtJnNZ55DYvU/RhHw2rsICjXv6e3yMgggWT2mQK2q7We75DJc+CrmPQFfw9XLf5+iZZjGckv9
DmYyC0iuFBRH00vvjHES9bXL2QJ9HO+8wcWx8sPr4UuttZZnRDCWNbiyXmQ7ER9zzfog40EtCDfR
Y1JYkC0Uzw/x/E8XMfzYP5XFYzDOq6J7AtC+NMCqGX+DTjURRmcseF4bYXe+xKUmysg4qmNk4JkD
75Izu0HLdRvG870SrB+TfHrTtMvyszFM48kVN/hGfHpDck5W2ewR/OFw7gMBuxt365hpP/Rw+f6T
2VoSSXPE23ZDX7ZVZ7qgckaG15fUNf1ti3tMWhxVY3WqAq28++MX50tGn+dRFvd+m8w3a3FUJ4Fl
+P+MRZZ9WtUkOcfeA2QUuvbP5duuj+DhxPurtEqMUXJg23KK18/TuoDX0mkRxcJgUqMjt0wl4OQ8
EtNolAEeqS8sg2/v2IWITk0hDNW0m0WaK55ml+pXFTnqZrHEZE87Q7dRHwEdvqabWYqeStFztJk0
uw1hlneZcnnNen/mOAAnqLcb369mYpgNtr4NKhtHVGNzJZs/fHtWvFFVP3iE2O7GhxDk0RLq8dB7
Fnsko+5JHk5caU5jZRmMaBtN6iBYtgSCSh1tdTKajt2AoUsXEZbj37SQA2zqVMRt+4ZHOWG/35NI
2jiFp7IxAf48trQKZ1yUa3H32RilsE9dIMomv5uBvXNW9aN2skvewkGMFJuR8KJcyZQk0mJ40nhu
rXkuztJC+v9YcXXrRiuxfi6wmbaUjYgAuIf40bsd7rZM6X3BOSU6lUqJJQ1hLQ3DD5XPuigT4gMw
C6wESikn0wEiAC9k59K4fbyAL8yJ+YGSBFGEaYekViN3hCyKZ+FwtwRpfs/qudxAzQ0Ke5hYPhiO
Ra0l1WcMRbziWPhcuZiXL/w33xuekeWb2vhWDeGYYGYzAj+tFZAXfNva7W/OvdbuPpHRXulgYpu6
a+y2BDpgEQpYpzSbb8zTczZIgshdaW7D7uJV5fD+cfIVKPwJ2RYJMkzubwycmmbrUlR36F8B2EPW
myl2MdesWbNGPgHSU92fa1AfeUUcbafikcXzDA4AaUe+kKJcqMu5KNZVAG1rkjzvdq4secL6Z/JK
tG2kGa1n1FsDUInk3MntmxvTDEShVbFfjkbej6jv3zjRAY6r5kCeeWXeK8K611W+ptPkyjMKBdiT
mUz94WM0uaEvB3l8LA3iXKgtPI1CamnkdL3QMlJzzkVDm3jhVxVtFLsOS3W9ikeq3t8V4bKIgRu3
pK697zQK9GfbTsEQ9VXAYoRvDNXmckrSomsDLxlpWVEybkRWeUs+5cNPL4MscbdB/XJb/L24lxxe
iErbhT4t/94CI0eBW1c9xwIFEaubZdy8wcq2YtIjVFRS6U+5kH9VjkJQ8WCYOw3Fp6h8ET8XE5kK
WP05uQnWc/98yUqfiq+tgzWXxoCMpc2qb+Kr76aI0pGq6xyWAXZjJ/+EGn1eQfhEw859e7LVH6Rs
avGQrguXCi1QBbSu/eN6nY58NDAQop/xJ0Yn9uwZkOEthm8ewps1LiJQV5xR76iJQFDroQIlHZK+
N1Uob5NFeoMrUEtYwhOwInbmUY5+IsfUHL3WdZ9Yuz6Ks14yw2sXMuMg1puy+zPDLkwHJ6sVxP66
9sCgR2FOdU5aA33KMTruozf4L51tWrWQbLlSGrjDpP1ieAubyuofhDOxinJHeMg4j2qnMZmyGPV6
60WCd/Ly2riIUAZCXwhFqKFdczp2anpJIeWOmQqqLfhDjydnkI/2g3MCou+BaxnqA7ISb2LhnNqn
/u4Q6DJ7Gc+CitifM58dGB8ZtqRkNdMkeWJEGxb21AkEQv2j18SM/6/CFqnZdRnfmUbiyoD0kGbi
V0P2zTsJbbooAzs54YOksQiKiADTKQRuA4QXxOndCHdZ3H2yH2dfBLR2G51siWMeRD+RVyBjmOBm
IZxWlhEjBmccq1tGdNVBMwfNHBkqoZ0ZOWTni/ZspbgI3U84jDPXBH/o7wi/yFMfhwKGe5BzJ3vf
rphADWCsq/tuyyeNJwp2Ca3LLKJzOwKO0Yd3k8vjrGthkJkSHGz4XFtXOVl13RkMD3zaIlJ+23sv
D0L5yawGbdzx2BGBB3m/4BkSz4Hjo1oQmw1ZGEmVw/nMGRjAcG2ybJr4AXJ1PirDZSyPyzYI2OEh
jPTj8INTLJJ7UW4kNKDKeNvSKmNx+ELXBfSbWVMl7Hkx3g6a7RYd8cVZjZnDjZ16+6aEzauenW2K
i/wkcW1NeJIxlIfz1lRh9Aad5SzMFv+obw6GrYNZGxA612d9JL65te1zqj9Bd1CLO3FVI2TKuekM
QLMn4D+u6jz7Xl7hjYW/CfvWjv2yF1x8YPMthyZhuWnJrwhTkLo/293+kF+tjRbGxONueigEz8gp
CFkBJo4917MFPIQrxuOl9oOAg9HBxCWFHv3SmZJukYa5ktrG6n8L/115n2dUrwJ4MuIjb+DKVVeh
C+AbakG1U36T9tLdqtQrtCE0DIlGaxTAeHUuK8NmeBuZXQgX+Ly6ge57z/rmd23iN8gP5dbLN7/Y
gyB68EY9DeqZGp1NYfkGg9YDhdtlUsQnypH0G80fRQ3otmV/9+yFZ33JK01Uo0WJVTFCLyZUuT4T
gduGRr5Zf81GChgI9P9MhtJfH2yUjBnueHMyQrbwzSGIvANbJUvpg7tnI/UlPW4IHsAf+kX9quuS
EzGwiXyWxpp64hlsw6QXUy9MvjMjvHE65LWmlXA0EbZfkpdAVWckvAuf7AX0TCXxL4+S5MMJzHtV
Y17THLRCFiaSJtIgxM5LsAzwWQTxzdLVSYQ9xeuXSwmLr50883oYY5XnKf1Y3gepkv6mfZHy/f3L
BePoXT4zGeTqWTKgNE75cQolmPHwlAQFK03R9JW0moWLUJCcydqOk5NOS/RM805ET4WswT6hHzea
oFU3EUnHCSHUfCWZeeGh66zpizA1AVc4l8o1ozabD0iRK5TURI9KKooVSNUtIi+PD4G41RMriTfT
RZf7vNI5038JenlTjhQlKDBeyCbmwrqBXP3rS9YFbqrjRsLK3JLo0eRFqKnl6/vVgE0kKG4tV/HM
tEyCqBItGVAsrbbM4DDWkvVNPLEmlgKfa6LMvKDUw9+FpHNb7EH5+3HKrIGYCdcQ9dfyonFAE8NY
zPttK1fymItdCWQvLoOntMu8vJgIjYQ/SRvzHXVpPk9+E08R17myQJ4fMGheL2t1dx77qHBoDj3R
PrqJDlsLKZUahlE4ptnCLDZHzP4kPTcpwxFLwPjhu5oNzq0u6i5nPEHjOhVlBSmf/fg13DgWh1gA
UfxBJxTe3x2XPQNaH345Y+KgYLpp6Z58kNAtjPqfbRsgSvr7R3uu9f08ef4RTaQaVC/TwmWbLUDJ
DN/STit7wPAcKXcIxHBk+butP/3Y2EgbxLgW/oB9lVd/TmOBpcotS5d4I0Fd/Pmnzf2zF1l0rwhH
fMEkvKWHa/4S1fMUCObCOkBkGCVhQprlDw36bfeg9HSdan7GSDXDcrGy6CoP991d1d0VDruX0GYO
Rj4IEdSvoHJpwI8jXaO9h+RJQtNjHKDtVGwl5igM2vaYhlEX8aEjgTxy2QZArlQj+tuF/uBTXMOG
RfKfsm3bfRVrW5yXbs3pZbCu7dMQS3d8vaP/eOSc/Um8FJntKeNsNKcZ6P9AHaAvIw1udIFNJoDm
HlZjKS13ZgZxGmNVPrVoinlzmxduoV3fac04nLltcSzmkA8t2S8NpnvVm4b0jqXFVTjLfP1wu/g2
JAQVQBiDlRMHiNmfh/KpuhBzMTrqbsi8zNZ6n/mc/RGRPWPieaGA12cutR7JxNR5JQUBVy4P/ESM
sW+MeOSPbpHaCIh/KS8NfBS7i19K3pXKas/ep6/hNFN6aOStT6IedGDSgXgGmWV3t/jYBN8Azkc6
/v0biER8o+AYt6eorU800jpHoPJVr7xyZ/OwAOhZ/sXAMwA5pMxiSbg6fFyHiLpiBtopdS0+Qn34
Jco+L2BF0AS6PNzzjL+EeEc6z+qWRNhNKPrIi9P6b0r/Y6b4r6as1X0P1pac/GucpqHVbr30v8yL
fVL1l4qgoQCsvfoG09pz1DIuw4w6uD4qszzJGbphFHnbvGU9EnYBlgLHWaaXsGxXC1+q7H7FuLwA
DWbuqxk38Dr4x9sMSazc3SVuDVdkIyQJ/bC6qC0jTQSfai3UstudDy5CH/9T+dsk/XY2rwoQoFo8
WRo78aePKDIj5zKI8BBxWoOe/mMw+bJTF2zZYiFEZY2YhnuzirdfAupHxcZj+ffjkhpZm59MspWS
BxUpUDDe/7Gx/KUSzSQ1M7xi2CkxMiFIqYqQtGVnJpxXZZZbV/OGJBIzWDHUnIhv2ZugDkTNLMO9
MKDMaXrCyNfazxIDRfqYWVwjg6kZ9tWuAud8+5OipVgoP9L5luVGMFBKr5mZ4rhJrAK+8OlyNANv
aF9Now4gAP+iT+Lg2pfAeSHtTjGKdTiwygya6lqTyejaYd6E/h9VsGUlzPsG87TSosORlOZmo/xn
lMGXyXJ8DLyjc1k85vAyoOPW4MXENxOnZRPxSdvVBUGr5ugkX6kOr3oHePo3Lq8zuTAZVwbx/ZuQ
G8PZBOIz98VZ0I5fsU4J+W9FoAX5pnqaLNsGi8U9HNxCL2Ca2OQzKDaKop0Xo5LG6PirR7S3dUv1
pZLxRJJhDU+LAbOsq2SQWtk466feGFdGiKR9T6KQqRnWEzSd09jWL5EjDPMcbrdfvqEekJAj1ySE
D3yzaCScHQi6/H/QhFYB5qzs0eCZy6My8B1y14LXbldp18JOxMRh0br4ZNjY41nknVF5stRj64I0
kU32Rn9VMMJQcYhmTUKh9+3Z1SRHjUZWlPsRhCkrSl/InMW0532otEU2TqHOfZWZotY6cEVqJ4eO
IMBZKI8gFxNgTR/KwLYNJLJzmYI/aRktj9FU95/aIGwpGeRR2tfWVrqkiUou4epLkoDyVMVGYnkG
8M6z7lFZ0NhxS65oLRQdLt0dHk/NJty/iZSF/2Thn7JREAsXiWlBOGkvvddlsZB/kFSZ7SlslIq+
35Ry0D3c4BiBdRTrj+0/XowPNULWN5w2ofbGg8xTywI6myyieLavH98ByuogHhW8/W7M3fCAvTVs
aj8tnd6C8RqlXQXGmKKUwTL/0m87PaO0qlcX8/BoZkRnZWUVLnpUDbRv5o8CV79iv5xRL/C1HzI4
F6ykh1Bk/Y7K7MLs6/hg1wSLIipZgnFcFW0yYY8dfGSNlAE+VCfpBgsFEKxfVZWzoMdQt+D1GV8H
CJDKnzib6B9Jlswe3Drei5AEDF5nn2QAJ5pxY/Af5+M4rvsIKJBvYPvrh+NOTb0rWHIeAt3ioc1i
BVpGASaYmY2qRNLpdzbszgTZhtqWNt+piCsxTHdwrtgxlwodrk1ambIXGA/xsBHF3u/G1mAdme3h
y3DVNWQyAUvBdmTfXJqamXARlrVM5IazU2GoVSOk7i3dhoGGM3ZahCdQiz+eKROFOAmqhmj3gLzi
WaF8zi57OXO3K67U2TCuPNQ0gAHVCmUimu6v+hqcNxbLq606BLcEOZp788rYlKjbKR/ZgpQRlmhX
nmAl6GdwTZEDG1aHtKc44ExEDmJjkUB/T6huSKjbXMX6VJgPa6zcVe2tXENmn3TShjz6ks4aWtWr
2Bmw2VEWGczdrkZZ1D/41809YWyxzUW8JlA/IrUH27AND8uc0K5w5ykEkCDGwZmZTYb7M7cEl2CT
8ON2ZxhoBAWUXrF0EoLngVPgm3GmvoPQJMYdqM8LhQzLunYT1aiQNWUZ3OKoYTnbws14v/69iRSL
wBzRxPpGqoqzuyYvAi6R3wTH20rWUwtzLj6WVvVkEWKdJWqwSt8+7a22hUnUFpZlw+WUnICOPqKb
tHAkYXQYwA+cpxU/uGgW2zU3Sih2ldY8A8QLADUygvztJii0im+u1Fl5/J1AV1g+W38udODe0N7L
c+DKg8nM4ljVef5SvLAeYznAMpyois3s3AKWE+jKpHh2LlqX1nhPMJQm+8/Tsw5KKjLMBmJKKcyt
TyLhBpTD09mFf6B2hoy8yf2XzQijkj9nCxlYnPKIYg/STIAGzSRl1cBC4Q4AdMH34lyXp9PcdvdG
VAIgl3TrgPzU9+KLIME2NorkJiU4++gL4DSY1hJRMcLk0DOA5wHLHi139MnVHoWPzqNz8IpTXxbo
ENbfZWOmtligOQUy7quEDLcNevNxxAXbtjuxirgISsxhjhQ5Md8Qe63k1lX6g7r+Z4XRJzgK74zM
cN1GCHEBcV5rpi6bFXCL/9aoMYnRY9EATJ32qhfITfgIqH4Y47ajj6G97IGCJ8vlY0Yzhl7E26FL
7HjsLudpY4cz9MC4ObeD6i6KPHxKns1PA0+gF4giaYY8+gC0W3GNjQoDFU0TQ2/EWNARqprRgMbr
SCpcoE0iEHVfBejvhj/vAF2ExrLDRIvNj5dsatCl8S9QSdURCTRfApNjc7gjamyeP/Bob4Nk5ip/
6S+e9e6vFNL+YHHbe0sc57ep4EW1mr9eCxts+JZ8+xp1UFQuPyL2KR2kClNq30M6j/O6pZ397ZFZ
lWOtgHp06C2lkcaM/nUrJKnd4OvM/A83lvfEI5u01hhkITGGxTb9ED+AIuiC8cx+1Lcvr41Q+KOn
vjsrZv8UCluTysNN3kC+9ZQjqv4o9S/lL5GYf0vTwgM9o7B7FNIQaooM0mHeW024jGh80ErTF8f2
OzH/sZhFeIqYi999Hy1b3fsFPDt0wFnb2wXq7b0c+Z5SQjcUi0mSVGFJf2EcxfRjZNQLfrqvJcYi
+xQQ9yX3fh9HN65atH5dxXQlTq6xNrLBWA9uzYUwXugZkEBtP1ewCuFsMM0uNsreWj6y6HcwA0up
A3jMLXbIIycQRZ0QntQDDaP0ms+I1Fr58zPSFCdkfHqdSAAhvnMu3SXycojlHRajmQxWo8eNj1Qb
stdPmHOsL6Yi/3wnTrYewIYlfJwzu2Ixj6vhdMWqC2mT3qMdmP7NhTo06LDIH+N1MK3qHYA3FI4t
k+oIyCsM8f3ity+Jn3NIdwDqvyYoias8Aasq0EOdpur5cu9cmXKtX+0JPyolo+CjBuhQTQwjix99
cgK/FHWWt32NbzRgsuF+VPXqamhGa3GR88m7CyPW0/osX5fHINy+8sx2cgxQgybYxEPMO2KAsi1b
eJkSWK6+KhL/7Wq/GnAmXHZXQUEvAKLTiLvVudAINaRa7jDmaf9F/akFxAkxlN5GcdL6OH7gJ/Gg
Csm4ZEPfGmq48rZsULXicynZYX4Uc5v0xTG59C0VIbBuRvqLMAqAPYRX30AnO4Lu1P0+mVDQG6XG
ZSuBfbFpQFjcgtebHmiCSseRAg76vmVxAAtQ0tinJmLZ5692COv4CondeRaoInqiq+s7xraFhYyA
r99noXLZAR+40UFQrTw3NyqBmww6tmm2kd1HwCoVYcvvSR1+KfspM0GR6idXCZ5JNFbiP4vqwy0J
qEmAIXuYpSmkCk0O/pd+nvNwoQOqLkZcQ/9Wcbb7ObySzQMRkGVj+dnEYKXkcb0mKBhtrdmpsllV
10fvTE4DL4Kwi+AakjzWm8y/08Kk1Ff4HOci05OdVCj/iG1nZOft1z4j6i6nDJeZzU9ir9zJL8Ex
RmRkHQ1FqRJUMPMSv7zfi1CxmvdLtV0uwIEOHP8uAQbVCZQDtaioXbFWlfvN4UQoh5nXFBJOhSB8
Lo6RJaYX67UT/OC4G69VuSDEazjl2YfdrLrYGwutktLQzyWt/nZRjSZYE6oH4LYpWPRJ8SyPiKKQ
ouQhcyDqwavN0q8uo+460i5YGamPrBclHEEKCbqX8oWkHFKByJ8iRksPqZpyYbiUjmrN+p0nG4Ur
CAY4h+sqqCYujFU0IWPqFPYhOy0mLOK39QJzu2SEwNJhBf9wclEa+HHeeigBgxtqg/rP/OSJPkf8
RW1Z5friWmwqCeo5BjLwL9aeHmQKTYfIxPIkwcUOK09W3VKak7qhNStTOS6dMyJzcEdkfci28roe
NEWgJU796Q1QK/F6h+FZRgT5nAyrHX3wXEyKk3J/VYdBXrPD64pGUxS3n3Zxdq4/5SFPrv/4BnFf
wxtKHkC67E3SPaLfkntYQwtAcPODjphz5yEYCCbWdzJ0RVDBpULfB74Aq+BDZ66n0C9hihsyqe8z
zzLRSyt8xVodjx/BBlEQelj//ZWAVC6JMYK+xvOgeZ6zl6GkGMbShyK4JCgzzm4Jjwxr4I+kowDH
QD+dR6TzPweNVxBKZOIDaDS1dUf3l3oTnX04eq34VGTF9FxlRMry+wPE8UHINz9diLtqqFxbSnGC
3gjalwvIwJFMmwX+nhRQ+eE2NMsyLvZQZbDlk+k/1rwvqHkG4TRPlBu92i5QG3R8l2Tgy8caDPj7
TagdWgq7h8z6hyz/T92NSGB0eAyPdC/+yAJrKhBNR7BgQLBqmMjieBEoHKrFJeFVfPGynZWp2vwV
rkQwtzTnUwX1goDJL/B2dr1++QhI9uFETkgl+L9WcPTEWMFMm4f/VGpqjJyytMybP0YX/ufr0nvZ
oN9PBgyz9wcJ+o0auzIyR+5y/bKs86ywegiy6Q16BmckHK2X6RnKemSm+isVDHR4cvkbGU9l6Ci0
ldE93mlGwe5SsXWOlM03EBnWiikL4G0qrRqBrYZk57RDMAlxQoiPnN1cFRODzvzbLU3Ct16Ht1ys
1JVWxIGVuoJc50bpoDER+CKXUncns8tu+zbIcgVvJOVPYTCYOxfh1gONPynF6+27iCG82bgjBmaN
AseriyfZyuGboe2jRQcR+g3mE6KlG5ze0aj924lP8wSFM8ORzC1zJDS8JY6Au142mxVcpGYBj+9R
iRBTTtekONELFwhPXfD+bDq+MvAxlNCOWmiwzyOMMwzk3wyz99fCYzQGTrF7RB3nGTygZFwGkQHy
10JnnQdyI9IHUjemSPe3paW1GwuaaVs4GSkeWNf1SxApDcbqYKq6BOcOQ3ayYwanDlNeU9w56cE8
5n4gl4oNvGVkZyzce+NgVhaY/FbwiMcAa5Yt5wIs7G3AdRitGCWDy7t5Mlm0xPYeHz8+jn16Tmuu
P6aBAMkOKPWnvWzdqcDtZwgMFC/qJHw+KVjEi0OJr47s7FHksywfMZMbwcrj3VLb7sawRW4Pt+VK
fbOTdENXWr2voDwIlRm9Wqu6tkp8wvlwkRbpOZXFIwtSeYHUkJ/FygOOwvU2yd3c+j19pvowShIx
PUUBVkOs0gfBFw+Z0aaGQfBUXNAW4M1+2qHZBvYh3mG4Blik9fGfzWpfSc3dGvk1VlzwIf9Si4rQ
oia1gcVl/T4bihB+I+qJxkFF+4WWYZR9UK2/p81G3wwQLBvI44VpIBW3+ZaVPVsVYEjbCBqq0S+/
u8vIX+Z6fblht9NifVMLGVBrzUt8Kcx8qI5cVGJ2ItYRGVWN0b/GBFHl8dqrDut4ZbCdrgCvTWt6
BHeBByhNljXiw1FFltComU6iAiMd0DIekWl1Hs3nJgWWzybw0ZIMbMYsIV1uNgdnRmxlGD5rIYae
dd/4qpXH2BOuS8u3k4dn9KQQomFgJgUppD+w6fwzlMg3Us0ooTuqvJb/vh3V3j9mh58YxhwBq0wz
qkJVt/8B+W3rr6C2E9jOaUTVN7cmEpHgErplewbH2aWkRroqoFyu25l5fvrltuisngZmt7NqnpQB
uewH0vLC8bAahI8wKowWr9aajFM4KYGiCHu1j9wTR3EiJHa/QZaOrf1392XrSg/4n0jyVNmpSta2
EVW9rk4MRl8alwNWRVxbMBKN7HkudViPa1rjVnVl0y4xk49hPLIY8j3xqK7AqR4zlib5C6woB0cl
JJbhq5qzG8i310yIkKivTDwFjiVuoTp/iZj1wq07Hy4LImLrVs8t5wcKa60h5Pr3ZEpKdr6Btmtm
dD64BoUI9DJylt+w7OZvWmsbicOckoNfdpzAPW6Vl+rEqnfCsKfemzTR4+6dkEawlO3VgNNLld/v
odhwrttRf0wH4LdmZdlAQ/qmKCink2Oe6EY53wJoIVX+3Q1th8Rp9vAPt//FT90gZfuZHfzff7ww
o9qxWc3GnDuDukEt5OzIztSDn30bQJPlhyP4uxMS0h0A40lYuI5R6RP1o4wmgncg4qBeClKQF6C0
hxChAfOIPWYBwzuhJ9zVZmwlI2J4fMqiUH6MMYtywIGgx3kk2AEwkqO5fuXfnTRnv3QNj5g6aOFh
qqNYS+opG+iExZpJdv7RF5sSrcQwLUigHja7wIaAmO0gxVDGDXlnHJkoCpgQW2BiK0k6rBDb4X4d
FwheM3nMlGfbVbX8B5OScwLUO2ovhua0gYUC6PxBZihbikWqPaJ7NJREziLpaVYURbNIabFpXyKz
IybUtnM9ayE1JpSmUpw7JoCBm+H8jv4cgPjtuHYmMgWheWokHUR2niFkU/2LC98dPXWydm31nCFf
+EAOz+ckztV+Py9aYRnwnVJJK4sSwvmxARhok5/n9VtLHWvKATW46IWeSO0a/eBro17uJx69w6Sm
vakHmf2RKtZES+wCPXXh2iyw5mB8FDKmj6Q/XXCSzKwOUAimIgB7mrWkmRjrX/hugm14rYLOZllQ
9Ruo8caxvKjK2mtlFiMeGY0tBuyPlmvbsw0gM335Ab0zlu9F8qQJTzad/dG39WF3mNqcbo66ZEtQ
Jl577IO3Eqs16Kgjs2l0ImdRsytCzIhGJF3FqwZO5U36TS10CVCkvf0Vp9LIOcju+nAUbXRbySw6
28EfPToE8cZVC+ySuq5VSS0MvLdfAkvcEz9rBw/wx9zfrwWTn2p1Dn0+JFsiY5bO7limpDnky6jY
SpJry7FC9dPi6GD5w1341jyU8tNu/On/44u08ZcfR/xcQIOhRwiPB+xKCDaIGCZ+C++3D9leR/uH
37x4bPTz9d/aqDISpve+njfdXjbCCk5DdxnsY2GzwSBQCCl4IpYp0Ip51uc9YfQ26CkBnh4d6ez+
GYtpi0XzdzNWTXZmX5zDaZL1ap/ejFeKz+zt76e8zybsy2atp1gIa+a77flHJFUo9dRf7ge3kCNq
CrwPHclfHOISEema+KbeFeOAYISg5N1RD/Us06iHVg7TUe/c3pCozclPWKkDJEFziKPGJdm90QIT
/Ik1M9acDUKhQi75HJhcfrLyPQMDUcBMilTz7aKRa4RhhchbItfyWZ9MRXXFIa4WQIyu2ba4di28
C2ICy7E4ERYHre90viXWY7JRuC7xt/iNKB3cluNcQZWW0hPDMcsK1kp33Zi9J7TXh6n0XI0fMA9P
7o7BZT8/FB46/2Y8V1hRjOsb025KCkUJ7OO6vP2RmhLsTiEBvxbTiAkxZGDuh2Ocilt4zK9f+d1S
uZvQL+Z6TumnJjw7j2uMUxKeGaANk4t0co7hPoQX+VLYKGtMrNmwhWiQscjBh71sP0ZgE7LV/Czl
sBYARcvHlXtniSK6v1f4VnR+1IIpZr+Fs709dTuvP6dZjngT5FgHFOYW8B3JSR8WwaoS+KgSnepJ
1hMkfQ6cly9Eh3n1MmHSF9mYyQmCxddEh+kt98hRAlu4g5MbIjgHtSt4z/TTxpt0hqufBuxf+1Hj
teBr1tNBxtp3RKtoXd9ODJA4zYO5jXo8ZfKjdABK8pIywB5vx/KP22PybJzPpNVBMYW3G/neXw5G
jtgHwpBXj/vom+uvq0rJ9sLGwJ+OBQy1EkwZD/HilFZrsLCvXFxETKurMz9Olptc52WFfWbPJc6V
mPe7paTtKjEanCBgRLDraiKi7cfaNhWRlm/zQUj5XYUrDyM1Bk8qzx4deGBAFY1LMglhdhs7RAZN
ipAngd6HlCaMsMTQ4qVkRjPQ7jH3DNFT8Vz+rYwJE5YYgB3ywCUdPkEfHsI7S/xY4Jv0csnMLo/8
HIULprVQRgQGT9/4Tbza8fRQynq0NIjzTwUPVO/vgt7+q0pV7ApMdeLlT3uFX4E0TNvC2COkZ4SU
aNAFLzQqcV9qWHa1A0mXBLZWppMJtac/RCb9k/f7FHGB66YRBuXLhphOUUJl8pB8uFXi2Z81z6Je
yHRK/etf+5Q3KVn8byTtF4awy2XX5Ik1KL2o4i0RFZaVodU0VH/bjwamlSgqHEHkMURLGloCmIWJ
lBHAv9a9Gpbgre+V5rAUAsQxrVjiXu0A11BEnRQuTopd8+RwPd76XiO9vdHXzpF44XrUuPDjw+ye
BmqtLvtB0CwTm5VuzZwNhiqCXvzSSAhiUn80hrCtllOu7o60wYVVc7WH28Cp+kc2LL9JWF85S11q
HJMJN72YjpNwBU6i8lJcoIA7QmbORvfsU28dvJmOXWsevqYei/aWmj5f+speT/AfbgUzGlbplxJR
hLftpfguzUX8frxJ+qQAq1XCTtPH2A9s2Z37GxaTSH7E9GiJaWwA0eMkHXJZ5L5brDAf5XbovOvh
BlQpqxsTFGx539l+yDW78r1rAyaBApnf8VqfJCNU/nvsgj5SnGi6kkXGMaHjcpIqWkRb/NOwsWtl
UqE5yOCcgGo+0zsBLNWMOLtK8DGOdzY9KNkFLkLL8zGrDjbEj4Vd2mxh/h5i/bHsBCf17atTf5ci
WkVcVE81aI0RFQhbpdewcjK/EOQVNHLTgsQa4EPg6+32dkNqCleJuu3YdDwli1vpyopRnWc04uK1
XUXFFvPSpSrtjs0b+hejDTXI4jQvEc3rstKIeuJpq0rN9tAwUfZqtmy1H1dFDYz6ItsJjx/Rtcwj
roo9EKchLsRgCfXNzBKTOJ8/OurzV9Vch6cUbXPa/PTFAFe8og2X0n/GY/j8yGmsxNfkoATK+Ity
6mg+SXlMGvZ0UCnP31X94Su1xgoGFovwkt5UmmyqkyCsZ3Ge/5mEJhZTAcTl2Y6zUe7sPLJ0K7Id
F4iX3OeFhglgbKlwHoSJtfiCttmHscj2YK7RmMzu/MYpGpsF2Fh84jeKrkd9b7aF9lEZfMFeCiSU
NJ1OkCdba5ca6BPDkadjfNxBEPBFDgdidhcqwQ7y6rZfaDcSfyXlzXz5Q1JWRA6I3m5+NcLRVbFm
XFhsvC9ixU3ULPZIiEfWRCaCoCXea4iwiRt2KsjBjzRpKOnmliIrG5PDuwnPpd/3Kq1EI3jCAevh
zWyxLYGAE34Z34RvfiGqvZRbkc4dkl/pC0g7T5kF5PUmhltegvKCSwOpZWR+LDi/gaSBB0OVxiTE
XoYCrFUGpMau0m7KNdIaDdsY+lHV8CsMmTKimCaIRzC/HBYHcIpXZb9ZoURXfWjUtEsEGvqi8fl/
iPiXPOkm3YX9BKikEWNugGDACme78gB1yTs1yxuU+SYKPRMtUC4SmvXKcy9ti6W2I6ruSxpagdQN
L5/z0Z1eFm734WPJcxBq0Ef1JsTztC2RXBFK/hfmAoqa1yrrOk4sW1D3agiECeTbpoJkBB9d0zxA
eDD5k3yB9X0GNlLGq9rqqEnSEbwewS2Vhi0hKLD1/a0Opope69eGJ7EfAHKFRdklmEJLwcnvX62t
f7QQ6s2E8wO588OqxsaOV3F1j+Z2n8UVL0BMOc4JL8qUovJJaWmGoDQW3VUw90Ov8ERkbaLgLPpF
cA8fjacMnmIYVm45syvrvE2f/Jcx7KQDqr4NWHyaoaT7piBGMF+v5MzPwoqLch3VP3YuqozMT3Qu
H0i3mj6sKEQPQGSv7BUTymx32XxM7SrmycUfk9YiipKK94OyAS90Pp2pf3CkZjFY45dYa/66Ufly
azKBeghbMUq1D1l8SBaHwFmyvUeMXOPDrndSkc+KZqyUYHX/zgylCAK/ujO9wkhidWQrSm/xTcl+
dltxTzpqzcCGzBubf7ow+RCrN/ho2LIxqcmxAnj3D2zNdv0IS57FLW7jLvA1emN18Ll29Szs00ff
ZyQNW23WAv1aFHJREW3bSCeZC5UWdvizKyzbw6Z0nJlxtMF1fcXoCbEyRfVLwde6yWw4QMLOOZP/
QgIbBAfIl7iPG77/K2Yw244vKPd7HL2topJPH64XNWmX/zFLHbEKyqVYICkHdihCpJ944LuYUuzt
pqBRcl50IduLfsFN85ODOxNoNqKqo2+fwJQSyB3Z8k33PI5hFr6CStJWlp2p6HBJbb03vulsC3Nd
428KyqFYyQ4jgPEaNNwZWhP3QdecoeGs/oQBycdNWjZU5cj4p7spJVFSc+K+CYssJORgdwT6SB+8
aqRNG7AZQct3ce3JakUWArkXKhNYcOB++Ut5pCu/sUzn9LiFc3h2BlWce1+KPDTb4VdjOkiOybJE
kkR6r0nAs2Qjir1tezC9xUUT/iSKvN0VkzCBpHcU3lwsD4tQZSWDXOIg/MM1bUAuoFXw7hu3atTO
teq2yOvk/l9K5PIFJWVrcUBAU9YurFuvcmo+cF9VWrs8mX7T7EyqhyOWCpZAaneisQQ61YhJoPrY
HVNozgr3fMMd8GfEFzlAMpFQHs5tnydYpJWCjRj0vEeR1h2Br0P+HekFBbacZrp0OggMgr3d2s6B
GC2d53B4kHsKzgU/pQvoRr0wOXRsq91UqLJ379jjJFQO3iXwQ9WPNo+nEEWpfwbbS/NyogRmI+2u
NPpFRMeWDWNuD31Y3RccjgsmHTy9tbYAjkSNZxVY6aG+npVupmbSMwPbcfnXJmYdcKQCjEdugpAO
1BakriPz5V622C5U/0JgMknpyRbnhG0/qfad/fYh8tUEGnwCphtvwAklQK64uWMuNt0dszXhU6gi
eEEEVlXli+d7fhCuKpdv7njk3H4pJ6f2KCKtNaYlEWeLu1UY6TjwfLooKX4i15qaNloz29csw6mn
Ym0LuXnWheIXe+NmlVm3y+KH1f+DCoAv7+1ecOO0TJjXjVpQGNTaQxpOTV5FLxbXA2so3C1pTsRA
NFoqYwRKopV22Y9Xcihb0mA9yLcxtho1Aty6kjk22CC8O1NTT8oy39KOSVEbW19VW1Ffp6w8A25n
AMu0xvFP+j2Y5RdNtlk1ROsaW530E1ZXp5WZRu0qqYNpn2cWKFkTdojJg/Co7iqsK4p0tjDACEul
336ZTFxVkc5kEBOXUZxE6SSQ3DX1Dc6zAWoRNrfoi5GxgbsmzdDb7nttlwQK4oXjidWrmrLrnASo
PTQzCEFVdmEZCf2iE+wFpBMudeHGwZDsxPJZWNmhLLbDH/sGEvv01fCXFBwTkF+wVumTOcu0ZYBJ
oJRJMJdG7KuK78ZHaq63tC1wgvyWMfzDgQgEiNpVbf5ldNrGarR1uF1NuBNtL5QGGlnpjcT5vU3k
oYb3EGMzTO2f5jVDn78NOkNcOr25UIZbrxU0dZkv8M562Ba/mxFVgEpE4IMdFABhF9KhXr8MCyGP
M3vjegYbEVmmsREgkP1LppVPGhvkQc4mFZJh7sqK70VzeSa07Fyvz7qhCaoBKRhyE7dCFKCzW1cq
RvGTqm0l7AbJAya6dOAhw80vgWO4EqfyrTBC5t8KbJVtJeBgEX53d0KtE+Wx+Htqyyf8VU/XZrWK
s9lBqXLKKMBiRCFj4MaEVYXG2TtHk8ZQP7QZgOYUT+xW69BijC18Ba/pkehqHv7SGnAvdA8X2g6a
l8NdrheJBx6szuGj2CoCGOH2cAXPnSS43EGrZF/c5S8E0qYy1WPNqyuFsuoayN6uyF5iBYEiMa/e
r+Kl/gmtN/ZOxM6eYB+TeFlDq3+cmWPP+DhmenODg9CMy+geETlIrkzsec5GPU9B78iZocA8JV+I
Wss+QoRZelwqPoNpHNATeGThLTpuTyWfv//a/39N5X6S6pvRwqf6PCg/c3hMxihrXw9IS60bthYU
IEX8Kk9bfjSXwP39Imq9XJj1s4OTG14f5BE56hqQgtkXtJMJlBZ/uvzaqxE+Sfov0jqDdYGnqkCt
P0rZlLxInyG06WOS/nKFw9G2wMrB5H0ycRpocJAXcsxh87WMFdNDPob9mqCZk8r+eBIo6egcsIEN
Are/2KgMVwRwKqLlXjlE5SM7NCGrQx9cv7F899eOYoKJCCq9Fux83yxz43wnwiVaAy1XqWIP20fk
2Eu63uuFhQrFl8D4JZv2PaI9acTL8PGSklLu4bcZeqBfk7boppvut+TvJ5+118pR+HBfUX5Qt3Ey
Jg4aFv1aVVmN7iLxfvt8SNYBRbHMOGWXUYxPhk4fLyisr6szcgubfDNZLw5QviKtcic7XV9RxwwI
feAE5LDXgJGsuUCVNnMubUWiGj58PYt0xvbzID7eEvwSryiXWrZphpXPSevb8waNj6aQLzhunOF0
2UjRLkyp2o2DxXtjtLWyAA55c+l8uQhCWvw+5N5GGJu8J8GGZ+9FFpT6DbeuX53zJka2v5EHFqeW
RuQ7VmYbc/K7p2IgliB4SHTV34JJDqtOm+6OzAcbU03OwUu4Ynk6kj/Gu6O2h0gRRzmJnCVVmu9J
iCmOmY63UN/hlNVT+sC8o3Ml+UZulrT34x6b16mFJYnW6FvCkl5ZKaZrWGKLaeFTh5QXydPGoz1S
HrlxAcr3IEAE/2DzjYlcBEMW4pSNJEmrrKnw+q+F+xok89JfeiRn88HEDGxUUWamaIzOcF4zHsSZ
AtBqyRAgZRnT7GcaazmXrz6NRGgKmP96i7wC8crR1uM+U+bBKvLGWAjGtTia5mDN2kEEIvkJVse7
ifxsONVAb4GYKeODLQBeOdnbTzTPG9CPpVR55oBpyrHO4BZ/aJ7a7p1/Ly0jBLIo+x3B3fAJ+Jzf
bqNkbo4NSAAQDg436gMeTVuFbAjxINHt9TtujCF5VWyDzwTAEj/5mD5XrCwT7E9vX06soUpqeLSS
SR8XDobF1uF8dQdFRucLkOdvKnkM0WEBCaBbmHrp2tYRL5AUStsP4Wfl4x8LMSCVVrQFVOvJem/I
UbQaae5t78Y5zB/i1JEMijlEI5IMVPhgQi4oy9yAFcaK4NH7CMBKEnrYrVuJ8DdKUGc2+RKfsTih
lIfUxI1Tl3r7JEgk76obdcbES+iO4ZLfc4wzI/XfzlqXhnS1N9gcNTACN/p4eY0Wzzspi0IT2Qzz
JIdRJ9C7BMdLqKx7syagkI1zP5nSXuPNj1UkN110u5ekex7R2SLCbNWeX7gOrXXmVCetPzhKHOsP
H0krqfxy7rv7AnH+0WCjSVhcgBNPSaWFa8lXa3nbQPyjvGtE70ALVtjh17RWsGMEbR5q6Sud9RjW
FQLUgvxt95/9252uDyrVcyHx5rhmHlAokTMifKPSSxLlpNDE4tS54ZtDxWXguDTGDs64ydKH6hAb
C8DQ3pzbTbMAVcpdKnLMMcvYmjfylrHmQDyNiLvJY1t4K4WHhNG/CTPYqNrF4SDXEfjs7aVYvRsR
ZD+fjCpTWfoTFdvkRPO66RoyLqnP6DIJcnR4IvgMtIAP9piWIk4HhmgDUo7x+gICgx56MsxeUtXC
QVgXLDlkNRdQEHrDY+gbHDDNA99BmcgNRcDvJdP3Z7KPX/0AwKdah+Saelnc3A3CqmGHttGyaVwc
2HiQHt0wL9k1wX4Ll4YSp8GXa0ctxe81hyxf3N3aiPMfeVicqDxl0sLWQAor+1gIEa0lpcJCI8Ft
lqsfkVxfEQo1t7Hbnt6IsJfmYTHFaz9iGGqDKqNK8+h2Z3bEZgT3NCoqDkJ0G6GoZp4XSZVAtv1F
KA0SjQC0rTlaHp0DqoSUoXq86tU+2CJ+s2sknjYOSduMv5o4jDRexSdQ3mm6VLFvhXIrtESWyeQD
E1ARVLq7wJkFE44tVAOBz1M3eV2Cmy1xisH3jrBoLtWIfS8RX8uDkvVgz2hvsEi5BNPctJ59BGu2
elXgC51jJ1cNWoHqResyUHh/CX3H+1qnZhppjA3t52SLKG8YqBJzA7c6TlLu3xuCOVQNOUN9H3+x
pJc39bLlRv0Ib7CrV2aNAOTzv/wQGoMHczarLkdu0BnjDPZ8xUeivaetmmkbCLdt1MNrvroCI2ks
pF2xsUmNgGCitombAJPxQXilfZ4wiW6ACT0bT3RvuB1EZTv9StJgkCuGVsTrj42wOOirANa6QJAl
1EQ63qcsFvUyB9NhfQ2UMJJ/S94KxVDP2DwDH6XxRadDnBpMREMDc9PNzTdftbMk4zmw5P2Fr5bD
RInxz6Kjakk+r11y6AaEAmDg4LotT1E+1ykxeYv7bbXH4bs/S4coGzcnFKrBNS3huHvEp+wNERBn
Gxll9Qlqc+ezxpXetr1LACtpmXKl6LcUSTZvHwctEJX7EFHSlGF9JwYy8wkG6A357altx72GMLcY
Oow+dwhpWYYL880rUs69evi4J1W2GsuKK6n2rSXNYUa8G4Gxp1r6mF75MsBDJj1V6IXkomA/mrQj
eXsPnj4bJ1eaf5g120iJEnaG5E7KXyFuPWFCJ82ahSaEQX8NtEWprcB7EYCBJZH2MdSPPT5pAMN4
DQjrrzZMTbd/YoTv+vp++wmags6fDBP85+xqImdNDtLhvgR7TG20pSCWmknjc+UmsMR3B0hElb1g
9qRcLGMeJakb/Qn4/smE2+Rch4MVi0tBR1AZt/u2c/EUpbmUA9+Cn+kiJ5IaDj+Ve47s3ksrfztO
j6+Pzrin8VGUO/3slfkoD9PrUm93RYYW79rjqbR1ftKxcI8sDieXBvul1OntKdr4zgkLp4zTJ9Jl
SrIVggbo73eQ7azO9wCPPox85mvs/5fNJZiPqoQeAGye77TBdsiEtNifpK2HKaEbFfte2a6QzAaS
uhkJVZExQjrF/PwH3u8ZjU3iNwC7YEF1hNyfpWQ75JCdjAd3HfJGEuEFl5kNyi1uXUx0N9k3pfaa
TUCNrlR1/ds3bP3e63cV++nGvkvMFMHL+UiTXQd2j7k9nlZ/UP9L6SrpZnhFoxJpAYQsdwhaBRuv
btxAvVIaHBYFdi6KVh1IdzPcsnuoi8Q0bhSMHFpW+jX4pgFUjliMDDfxX/PPYpVMDKF6CP+XNboY
QpILinIUGMTVNE71iu8D2LuJva/gQ70lPLaTvj3R40sHd2AEoVyDyx02v2xheFj+vx0w1l5dNnuF
IWMo7dlcCND4yAoIy8FO/p/6OG7bjVzcroywHc7+V0MPk9T0U0+X7EMPLsB/gRVId6Ed16RPD596
Shgpat7Y4V8Ytf2ym0YpShtP/7d9C8YQnrBGb9VaqCcAx7an+pe0XJgR7rNcBXbf8UUNcO/pFfQg
BAt3Z8QsqZ5Zh4ZaPwCe67lTfY5XOLhL/0kmPebU2JaZOa34gt4ZSqxlNoWjUoL774Cz7roap8ci
iqf9LVLJaTnzF3xgNszwyIyOgK0dlijRXdWsitI2sbosJCBuoB/sjcEsazY2egsZjMmyBYM+nAX4
X/cnstKA0OTa2f2MFa+wTQoH4Y9b1z9CRKpvVyzfcfnHfRi9MZ0JyI9+TJ30hSscxOeiy26levyv
YWJkAeeeHu2bGqtluiNGZ5hj0i8f02g0jYqN3PeXDMAYU7cavYjfw6v+Rh9tRdMylZRjOS8/TwwS
H0Fh9vEo80q2UwX36RRPGJh+diEa3U+Cm944oZvzvTkkI4Ses2zDwiAJu/qpmm+8P/53s6Xp7SCX
YhJrpB12PNteq9DT7cGvd+12O0Q/4zib6WJkATEchIS2NL7JsSYLC0VBlToEhzSVPRIqiwb9eh1s
UZx4ncMSf+hZJnOEmS4EC98Q1lM+nrylHdPi50mRxfyLCFcXBL29BzQ+0iRZIKj+XlEOXKPu7cb2
84b2I0vrd8K6cHJWeBWBrhVakTeYLv6C12LWK0Bnmn1Us9N5ftk5YMXbuRsRp7XJ0pmpds0gFVzC
ytFrVXUw16S3m3Iz6ExqeQ2u67Je9XUMfPfKkefgRrxt4SHcMHudkmeTyMpemEUhIqmmUZkfxuoc
3sH9oNBkTp56sz8G7tZufcu45w/TBjyFM7B6TVsTg/XM1ZrnNvsaULYFDXBfQeWHRlfLZm4AgEVS
+GogBU3ctXVBwcUZc8UjWWqbW9sAQPxx93WKbCOxFld2H8OmA3fnuSQ8XSbfX4KMR4uGspXjAHak
hghPvLlS8Z//0H1CLRVW6xhFBwz/VWjxAVEZqhRszZS2+Kv4ABVPKAbMSBtpTLpz4/MT/P5GGnIo
4LPsX0VI/SVyvXHiGdLdhATgqDIIvD9x7LFqTsFifcBHHh4AA9meLiSmojkR7Fba3UtclQ/XAXm2
yMCFxEOmxaQ07Yzl8o3oZNppi/6zVsBczKFUQ5qBrobDA+ZlwFfeKXgyJevcTPnqaeON1cEc/tzU
BfSNXUbVz8ffyQ1ouucYf04SUUvD0C/HQ4rkRgA/yF5guOKNbCfxe6BPCo7CIc3zhytoDo3HIZTS
ktSwl9euuCtDr2UGQWt7Nkm+OBN+l4wOWCbv3iNx57VF94g/qyxJ5XgXZs1fyvb41vIFF6TUrw0a
JYuhzTw6g670J1uI8NywtQuP4w0V9leLnEmB/F8VwN0WvJ2cGv4CicFhzQpUMqTtb0Rp8lxC/NTt
3kFKbnZT4OiEgtMzWZF/NxGnlmDQ+y9Fp9o6fe+usIfxeXg0Wu770GckrSUGZiy1d0WeWYRGJ6cU
qYGPEa9veh2FUgRAY6LvEUPwsk+e753pC4yTh/D+DEDaotgA2wRqCMI9ZsufO/ta7DzUP6+klt9O
Fx13krCPvFAjW1A2px+hbHiax8ohUlT49CbSzWeV0ODHzQyiQq1IzqnJo4oiVbgTrm4SGGWzivgZ
I924f5KRQva5Olp4Zu5FVDr0a4N1sUBP4yW7RKLNbYbaYCVYEBuacxeN6UhLZ26inBzXhXTGWd1m
xJ6KVqQp2CE6VDZEt7zjHpEtIwvQJXsINRmOBdWlcUgEN7PhSFz00NOHGq++je0ukht+6o2a0wlX
9NTEi85tUrc7JFdfDpydncXbAsk3osgHpC3AgzGxO8GPzjiLjxiNvrMYDDvgVQaZ64wxIexF59MD
cgD+QFmw5lk9xv2EOvyAnYKkBQ7mZ0YMjxoBAoTpCyT6E2O1LVhwArfrqnvGDpyLqdvuV0XxAk/Z
XHtMiHKIs9DBBKGOXwxUCx5VZQx0r2XhTdefr97j5StLArY9DDhL26SA1h8JKiFiZ2npO1FoGKXk
Gj6yVFwjZ3/U6v2IO3dVBWAayiuIBj3JB8IAboEfY9R+BZD2UImQaAHLRJwAC23yuYKn759Fe2Cl
b0i1aH1fRCf3Iv9nfXHmAeQ68lMxcpKqFlmM6qPbu1M4CqffLGkX41B7INI+GclCYKSQln0E2Hcb
fNo97EfPEpXZdxoiZY5dUATUfd9SbgDxfPYM2rcINwcjV/27GIgekkyD6ho4R1q7vX0c3uhWt7Dv
cBMwSwdvPQDrL4Ly4s6E9Qp5mRCV8HuVLvyA/uJmGK7Z5NqWinahr0GcpzDN5LxSyXlIyC6pCtQi
tGYky1agvj2WAufUBlymxLHQAp+jKaKkWpasnPyxe5jAyvvSoi84pwaDybYT5LOGJFpEyNrha2Cc
RAlqAqBWlhovXKyHVxeF+K4AvH+cPVOW+rX/sEUyLV2VP3aah106fMWE4LM0ZBxfSWlxERnHU9pN
ABLdKReZfeyzJYiOrcbJ/AiLQVMVc+cCAEY1Yp3/O5SxjG8ts+vVhlaOwkCSJs0in16f/LI7RBLl
+FBvlI8xwWqNMzUUu7YhCIxMnFZcZG56kOKphXNbSe15xp4t6TD5YPdPi9J6g25fk+q/Gfz3DcbI
Bqg8GdxxvyZb2K9oD+DoFZiSgwC2B8MwbvzzZpULIZPcLLpoTxaJTDCjMwjzNE5NrN1qyiTaD4id
0dpZROn14XPriFd/HnQqSsMvYr/EpjzFmdW9OwAlC8u8vZhdVHN8Z866XwqDQe4/R6OoEl19jh+Z
cythVHsbGYEjpyJM9MH8UHtFODVmbNTU7bDNoF55wylRb/1bai3AFY+PA6hKvPhlsCfAO1+TVLxR
jvk5MqDj+wBK7pVHZouoUxT+uRRxZ0HG+IG4Si8yAUSW9Uh39/D7XX0Vcqpcdk0Kaj6E1YO3F4jq
oA/b+CHFO/BQ2c+8nsheB71CZIv+MOIB1l4isWMvOtm48yf8ZTHoRkTb9E8Lt+L4ew2kQkVRwxBr
+Js93id/qG4psp6uXAf6JRqv9RJ5fx+lQQwUPpSwI4PO9fgYWCD2NrddwLf3vt/tuJxFd3E78ACz
LsqDJ50zhk1yjy+wb0UD45FdW6uDKwr8YHOURvnP6JMENTqtspQUURD6oQOg3Ad9YuEqsGRR9D1r
ZL/Tv0qIC+6Pm8EVl0wmcSBQMNc9BKoOSx3PF5++B22+LpSZo2XnFvW2CA+8hu9XUM9y20c1DEKW
Ts6hCgn8lBjEzVbHrdosqOZp2UuWcaRQhiptSQMiEha1HH3S+bNapw7Edm3HA6V8npycPjwRSIwd
YtmP4ZwJEytS774rLXOqZ6fbW0DdiPATN+vsmItee0y5aNPYjIKTswy1+m6QZVYivLwqS1QEqDi6
TBOBu0QFv2SdTF9MBxqZw3utGSgowWpHdPGS5Q+5kCzdSYk4/ttZaKZ3N6xnJm5q8jW9BaMi8NOu
CWCx0C2d0UDdr9cSQqCXPMRQEvfHvmt16R1YJGLluaqejwkVdXizD6TT0UE+j/Clf3v0qTl+5Z/o
O10I4OsxSyMWq36qRKEyHFQYcOvz3tr5eAt/Tm0rltmIMWHMpYY9I2cN/YjbJQCUGkzySZO157Fw
IobLUXdyaSjdmIjcLEA7pA3IIPkCHRSb/kCE0x20U+7/a7Iy+a3Ek/ruF7xCaHbrEft+DD4rFN7C
X87xjMWvSwZ/EL9y+VpDDbMsTLIEccc5ZtUCiEBv55+8ru4ApjZDwJqvtTm+rpv7kTyPxcjSQt/u
I+X1d2g3oRV76FIZseS5MbDIEWdB/tKKaJ6rUHTgAOOAOqGvmlIVvut4ud2Wq0iJVCyNiqOE91lL
+dQgmKtttCwpLXRTzFbU7GLh/D4F+YrSyb7dZHxsFDW9O/n3uvzac2QTY3UUJQwSF+WEhsqOHLeI
E9rtiCYqVOOWoYQ4T+Pk9aCDtR8MfqAuyLVttbgs4sinpWRJDtMJM+ZVmZ3iFDuOoX7wP7IWD8xV
xMH1y+kJbZ4Ph9vMNd08BjycZB8g0BxfEjnoNn5ll4PSd2wku8Zof/LxkoAJlBPgssAAJA9T4B60
qZWO8mh2nWRyfZfkZlRhI+Wvkt9U/Jj0nAHzsVkoYZUAHS2JY19XmBlNsigAlzdo3LLe/poddC6Q
u6rVKCOf0BR/0e64ZAWmj+Bk12VKbhr3qSDPg+ikLdzD7TP1G+OiRQ3497/Mtu9qJq2PdIdzCBjL
k1vtd55YC2J/ptTYjeOFhCz0i32fvu4/pzuF/ddiH/lh6DOBUWxN6TFuIhs4KA/lL42C8ft8w5m+
qK986D3FfG8JdvBR+80j66jzdQ0tbWhOsiAbMLngJBLdhzwsUebNv6hBN/IoWuPIzIAYfcJzLo9U
9e1hiPapx2cdm+aaUsAha35Vj6q72mpyTC7aaiGT1KlpEfLS0CK4KBN/uj4zMJeUKi0y+wrcoXwz
GOwwUbvbu2oz17m8tXcK/0TN5++TU+v8WF8JzZhLfYNv5UGJUM/QNJ22aGOX9uD+X8PeAJ2nO9oc
/I2FVQYCNnr6P08xti1M7Gguy1F9fvx8oSdOLDBjm3yoQkYL2LNjdI6QZ5oSPJYQxPDsP2APWE6P
yEPef/S0txbaVQ/JHjPrfraXjJ31cPoav41uGuOhMSM10FYAnQYPv241ifxppnPM2FoxE2LiTMUH
eA2MN95eZcsAEpEADZ+fFPnM6WDiqhM8zNlNY9AyBkRdb1SreNtgsb/tSTMn5XBzH6CHA9Gp34GG
RtRVzgiSvFUYe+6polAfvVcaEHE9doXkDESdV2y85pO3+6q2VmKbTYzezt0d4KvjbAFMGY3YU6B+
FJUmn2orHJDJGFIe44aJ2pp51Kf4VPo1y4XUyLGXyau1NV8q8lU9VwnM+B/ZcgSjcGbIzB9xTr/1
6n5877hWj6dbRct9AKj/0n8TNBTluku985+jOqad8xd/CWuTIup3lgHH1FvaWHg4QgZYq2zHPKJo
Mp3xtvNDGM3/rXLh8mh+vpYXCih9a7RegWQSKakV7XgAelkHlPypCXmPGLW+WhPR7NsoMbLUIrWL
N3PNCevJEIP0IdQlFgP5HDdsfRyw38mGkdBZBHbMhP7WdxemXHteEhVJWhrHlF8lxmNo0oMxfKTk
uE/3d+S1oEtqzV7dBV4ZXbJDl+FaLPnec35SCafGLdCbaGv74El6L2hJ23G6DrELHCjzQ2AAS6C8
KGs6bO+soFJ3vHF/yLCjLtOauRtvio5TCgNR8gpl4RS2jK/PuFdxMTsCG7fECgoo/cyaa95H8Vm5
FDplZW59Tfu28DlHZD78s7cn381tE3Y+bZFM9+ZOJT/TJtFgQiIl30KIS1he2iry3yWh34XcAN0A
LUamfReZxgMWfMBPOVvFGkeF/qpkTXZG7qSsEyBxGkKbYUobDUmfLE6K7XguZPRNpjlUfqSnAk5z
l70LxI/7Xpt1Jkr3JavY5vusdkt6If7u6wxrhPL+ax+1I0u7lEdMTYiVlAwfOLL+Ni3ZQfbkYuwM
mwzY1ZdrHCyA+zvldsLDqdninfwwcznK24Avy2GUXXeKovZoQG00MGbpkpKo9wU+0705rDrYULPz
Gap/3rA44NhW/Liw3/tNaKSdOe80PuPcj7FxB21y7SNM6Wnp7OeMKW/96RzlTzXnfGgiFZXz+eoG
7yUmKi5psMIp7EtXN0u3pkgQLkTMGeh/C0T8tfUzwULWxbnbpp/EoSLSBoTWuA3yb2QXxHyb3WqS
vYO3kB2CveCiURPGr2vpMdVqDN3qqBNq91okvTFykvRz1PU3tdBVBcxT/KuUneF56IQyKJ5GXBxa
HFV4bMsHevRACMpArfIKiM3ek2TYjXdkXaqnIu97XtuLSs7epzkfkoRlZTy8gPYCayrelCUZ8vMW
eVXdg+6vugbap8DYEFjSWNCl4BSWDOhOtZxfNNbtZxGvAYKz6ZefLEgBfc49RmdTlJKHaB+R6WZl
5DCusbV3QgFA691dXYhAc8TaopRtQdnITmR8tHJeuJ85Xa/AuJTVOzC0LweTbAcPntPopVyfvb3m
YvFPXNt9MPwR+vZqDnCSTNItVwtn9i9wFEk90gs6NA+Wy3Ila2xpR7xlmSd3QTLKxm50UgdnzxRV
H0hFngwZEigu/jiJGyM1X7kON4Si59YTX/29fB3Mn8WNeJpMO2pTE7PgZqEb3J6B0LZV8hTWf+Wm
cumLtJbZXJy951EbuRqaV3DupYdnAOz4gIyhPqGwSQEDjd8M5lE6kiq0Abmm47NEIwL9yVsEiSTD
dGcgLzpMpgUw9gL9rdRb/1ZGEVAyOcf97rsF9iueCzSzxHM1hjxO6A+LtZ7dEwAzvb5TUXrQKOzL
ai4WIBR5XEtoqeCeHYQn9jq2QAkkdjjjswi+mbCZ91IcWXCTebVn3jeARoWVExY3J8tPGkv36vpb
i4EPwT4en3czfEw9lsO2Av1nmPrFXiPRBWi/JKkmqeuck9BLWVuRE2CoFdBFAOJ1Hj1ogeEnlO48
ue1qFGQtbn0q/WW7jA76BgSfUA0TBxsBGvuXGCJCsLccsqZv+pMX9FN4kMdhjm32sG/oVgw2H7Ft
6bB863nLuTMyNfQjwyxpjxWMQJj1VYvSgT8FZl1+QgR6zIq5HXxKUE50ZQjh0uSY01Z51vnlzaWh
RpXsEij79Wyy1Cmn2GWek77ZjomETua6O4McWjkY/gcznOttjymV+A/MNkTqU/FILdjW8tnrYUAA
mtz33ar6DxL+ORMwFAiVX9tHmBvmDCOiDrkOaftTOjuwIaO1nYcHc1C0JzRR9S7eGc1eTbz+tKgP
6ZwssiUb90t87bRwlGYv6Gb+ikQ1jalVOiI2lfCRUrkU4a2Aw60rz1EInNMGGqAY3Y/IBKTlX6ED
hSDSqLveZiGm+JmHuYRk3AiYDymXH/xXd73Y15PB7uBIm6NyZRe9sim3QQ0cb2/vSVQVXjIZ/P5w
h4Ky0nIhRpX99Qq2QggEtB9wRgcmTGEOqGSSqI5DE6hgF0CJ1GhvYW1KjHopTZ4pc1LQuRia01bh
GbVwb1isclhkpN1o68X1pQXd7ercVlVaimrIDfh4Hgo2+WfpCAYnrG3X6aSbNf2TxRyuRac65X/o
ko/1LOMbVUsFMK9fqBhcGIHQZmb/7CPeTxGYshICU/9cgA2mlD/GRMm8rZwIBbVwzyhEkcxhTHXO
ckAhf1nvYTuAZxWYfOM4gbAUhDXjZ0aWFhXZLvQNXAza/yxE4Pj18FITUkPaPaPo3PF9NKO9C3UX
Dl23/ttyywE0EXx4IaX3qaHsiP0LVbdPkNL3KgOa19BHakth3aYH9XDGoIAWS3YTn0QQRkCZlAAd
tpDGyi7cwjKNup+eMTP00+8gudWFADwYPLoXy+hlFwxmyALEIQ4t4PIJCtNDjh+hNIORIjOIxeyp
rFx99ey7B5llQeG8lMrrlZqjzbBmOUEEO9ztEAEexYqlNZAc8f/d1tH+6EuOgBVETGcCf6UrMttH
xCYy4dN8GixTki/UETQkz5R1Nly3Cm2Z1+8pwNETaclt9UgRpZdZW1rWMGrFpyUdOiovMlhwrxlx
c6dr4jLYSiW+e0TSJNrp7rkBGo4j4KDh58WnHGh6ItEFw04I+CGfj1Y8zBt63xxSRgepsD1qsakz
FUN8ZebC2hNGUQ8p//pjjFu5f6r7iV7zR44gfyLdUY6Dc84QFvmzXtVb8TXwaQAAhzr6uY9kCEVS
rwJ7MyU63E6EcVmH87s9l7v1H589o0W1Ju3K2e71aSesISiZrrhRM2SqdDVoO/gw4Fe7orPAvMH+
xcQffhdUWdjSaTMqN9jVg/ad4pTtujMWQ4I4zoB95iZO7R7rM3O/oC1874r9bltrNmLKfqeV0Aw4
O1SqaFIcPeKpYI934vMpyNvkMnb3qjTjbvl5LGVKyOkuFD4EpjDbbFBD3s6sf71WF+lS3cq0+Z5/
AaUaBNFsQf1HblljbZ/ZEqkuY1vbJkL/RMhZnRLh/a9/edL1Eixz+QuXYef+xTn7UwVnOkpFAlzE
A/+DNVK3d+4FiDWRpWJ4WBMT7AeLwse2yulvxjDvMdrHk9xBJS/1djNxRU2caZwfZEihBg2E2tP5
5N8ex28IG/Z8x05/EZqold4Lc779z0cbNtY7WW47rDMIm5UOWXa8Z9FX3PrRYMxzqTllGNGAjw+h
zYinzqfXKSuIZyLD9iRQL4Bxwf+PlyRkwwnIr95Dfhj9L8i2HMnCRTPYyol4J22wusAQWUrngSVV
urWPQj/VKDrRG4shJ86ZKnRnDbo3620KctifX6M8OC3qKl8kSk2jR9vXdCN34ndfbMQv+BVbUmzA
NIPwM+Xr+kuEyFaKJC/xX8TQ0kljjUTuYu69IcBwmbDa9RQFEVlQMpVTq53shtP8Zj/a8Cf3O0qZ
Wef9EeuVAg/rmkYQSycW0R4wN9SRI8ro6RWNK2ugb2CZBo71Q5y89wkue+fAXlf2cUiYywZNpN8g
73CbBmrAKBZH92gXIYslONMeudxDqxUM9ysRHFA7RRP4P7AbvLV0m+you9n9yenoecIIluaFcpni
DlCxGYx1fWHm1825el/FyA0txHZ8amgtM2tS0Gdxfo/6Ofo8kc80DqCxc4t5PWaWpsu1TD7iETh5
IvzohO9D0zNYaSXabKNcLIGKE6ftdis0rUvAz7AZ+e5X/8a99JZC6+ed0Z7ADJJC/2UT5DaK/hYz
tfttsT7lZnEPhCExs2nsebqaX/w9qK3T9/Ys1kxnAmtpexgbn7XiY8teCBVnAza3nLu2/6EONntT
6r5wFZCcvUwVevccgGyoVWlk84DLFP1HxHF8l7bLaLyNcp6Gu03eV4hhY9qclXIfJnf5t0wz/lP/
GygsBkZ8HaMAgGXaz9VQ/Xjn7z6OLEcmIpyHtNQSjQ3jjiAd2yD7VtG0hIkFY87mBsKKV7kzylzI
9kdo3ukzb228T5KpOt8hRlUwaM2Y5bU3YXs+u7RIMDNUByH4oUM1v9chHczYPUiQfcyqBdgKN7AO
9gOwVf56anLyPCMleUDbY5tCXsMzoTTavh3qpR6QWVUtX3XbPd9kW7jX+snAU2Tr9ym2heaMEEc3
aDwHwfXjJvbtCDWpT15U2LgCLKX5ikIRYUpXn9rdeLEAIaavf6C8OlufT1GyM64lyu7FU7Sf/HhT
ipWgaSrrWjt03z41PcJE34eP2u99tRWQxzLv4ENTQEuswYQFbl9RllkFAInrepqwOhvqQQf7glz8
LvcL55nEDlk/qEAjFLZDmZLpOtT2R7zZoCYwunRTRNLUSFO0PiDtfeeIdpBHkeWPMaERLTC9u4Iz
S+1vYd5oF4SdVt5YegNyl9MTmrH/ATr+DiVVcCSa/dR7aJLK8bl45G/E3W7r0vZ4rzMonRn5utIF
sqenEm6SSh+N+GOWlVvMEnlAsmDk4w7UlrsQ9wh2OA5MMDgclDfkUWVUCIXuFCLyym64cK5jKaCY
0ZbTqgDVdlAJC0a8vDDm/3iyLAJL2KaSbZEmcSryBTtSd2OSCvE6XW2npDmvH4OJbn4c/Jlz0wBn
RQKFlU0s/W6ejanq+Xvn5wmYnwjR+4CsBguRyROkRWLKkqz4JoVPsrCfiLGuSBfO99QorWWkEqkW
D+Nx7i+ThLykbJurDYb5jEUZxF26nR3qqt7kjIKOABkm8y+YVgtYQcKxdIHq+YVPuArRSTpO0kg/
MhBZzYReAbm4NKjT4uVRNdLQiNASmoMUjqOnKpA8myWGP69GYt+Ueh58jmr1fXKZ1pI6XpCKot5F
n25SIbeViUcbog1r59PSXey5CMniwVXziPxHFjNekWr42rNgRGvkHQqG8pqZsmsyoLrFgs2vMzdW
VVYx5aHalWZ45LiGlJm4B1WnmzZ8NkuUCxqlsRy9biPW8bUf+nBCnFPscUW0Wqp5W3Gf968dN/bm
iNbuQbd83GqXZxAZtrsvpXB+M6o5BiwmEJkekpSrt2dM2PbFu48GeP8F85mN0GkNu0YccKJdeeaV
Sz9jXK9OqZ0FWUf+E5IeVuBkHVn1+5yyGsvKNCjHqF783oBfLL32YAzK3M+ykucWFrfmC2/ts8aG
DIN03O+uYsV5A9p8TXMTKEQbrpRpuxZS/ZaAMI936s1W8d4j+Y93Ad1qyhw3QsJBGZHPFKrSuzBM
0wdMbiXQbkklJ6cTJsAMPIJRDLO3KBGezka4UPomVRiFWPA+wu+0JNc1BdkFYbljrCzoXLLvUivo
jpmZ5YGTx2DSiJEvr39EofpFdH9loq+4OdFZ4O/N9l1IXJtCCzd/weyQMcS257KWEJRZlEduVJWK
v6kFKjp0S39woqdtpKFVdgFuOU3nidyYYkBNe8nhHAYhrJpye7Niss0rwzolIUMkgfuY8B5JZPd5
G0fLHgF2n+MuJn90BnmI15cjeN1gcaWPhU+jkABgoK5h8wAQhoGwuEmC7WZaDJugDZIgsNDvX0cy
yKD0eHcNeJ2VE6u5AqWpoY2s7FSpeYMTFAKXlixqYDfkz+nHWTiuS83wOby4uy/NHHUnGg5DvmbK
j9wKd1a5SW595gFbYwb2IZIuAixa1c3ryTeaLGXzXUfyW+gy/HDq1GXMNWomUthKkOogZNk3Shws
O/yqehz5J+3H/6BLiW7cateKAZYYmR7yyjwdVZze4OsMslhOM2yIhDtrdg5DvL2VGNrq+J0mWRZE
TdLyQ0VxYk5/uyMYvpZGy/UASDBmWH5zg2mvN4qsCwEa9Mz/6PCxGq2/fljeoPNyVacGj4K7bHnt
tJlQW6zPsDADhCKsXgMeaSGedEbfxY25F8U98LI70Js+2wqTWSGdiP97OQU6cn9InLaKfZ+/Enql
jifAxLrS/gtKM+ZR0hgHZff16dr+UCB8T917wyyvVMpb7zlIrZF/naUnF0BVCi3miYvFMCXwE76Y
G/bMmMzSUNgP//4vZ24rwQLtDBzvRa+cNmpCi+kac1FgeYZ+vcerh2VPr3GOm1BU6RlGFLEZB7x0
YwJP/5hWcSqFM9G2drDMr2bUnL5gW1H35wCRtT+WfjrywQzEC8U8Cw0uoMOCVw23+BR4jrwMuWrd
PlnjTLK4gURN5htZbXoPK2ECHUYn7pwMKF2Pqn0+603O/WjESlvw82net1KNqWSjSStEdjXWPtJG
4mvXn787LJPZa2Z/wCdI6cQAovfZptpb3KQKHm7RshCSZepxPgw2vpBeQXTrcc0yUoKEyvSIg84H
huxvLZiT1E75fBYRZiiqJLnwkM40ytBCqnNia0cWibt5cpjyb/m9gYNteqaRfyoQs8GyVEX4hiQD
AHSPY0sZ02TZR7TvN2zVyem74F6JuKdiWzZs791Eoerp8EiMbCwmGk2AIxsM2MjusWDUplEGtsfR
Rhd6GXxpdGi6d/lWf+gpa01hF8n3gQsZ7NWt6O/TmFeMF53657Tj7huj1yGuZHo0OMh5NQICLpza
K05g3Wf3jo9NNy5HEWTs7ZJfYHRJTAFjobi+Aa3dnb0rUwu4F4Qev5jC0R5Q4XB+TpDy1J65mkwY
NxIcnTxBSEbWWg4o+vBFZF90XH9AaDBG9hwaZl9SqZ3Ifx+QtdMmli1Ioo5tpO3gjYjFBCs9nN4O
uXHgaOO+lmychk4X/SEiMcvh+Yk8LbbKOkGMmbPErlC/caf42FwNT4rjjBWPRkNyjHZPkt+587n8
PLr/U+dh3YHDb1mdYHz/XQnneRvQrwWBLAygOGVszwXyVDqsq4OlD2J3MHTYuomNebZa0Jbg1qq1
7VXDAs0l059TGj9T738jpavM59IM410WBxL7/31Kb5dbDhZbwGj76qHLdimaqPMRkM5A7vNtuza2
GiB5PdPZzs8zRjSqgl+3rE9KqqEI4cSsR2RANC5jjgsfnaiouPnddGih+EPgf7AeWKAgaxwN8R13
efDyXaGQ+BhWV3R4NlAhbft3EfBoH/fGbUDzKaYF/FNpcGc3fX2Z9u/Y7W9VSojfFyKnCPwHyScC
a9k2NwP3muLGkePPjwZdI4v42Cwl23G49ik2cg/4c0xPVGaUI3+WEh/P7EwZ83RHaxj1xEHWGTLY
vffjDFs508cAVOljDMJDJGcloaOOwjVwPqxAvFkM04iS0N5YcN5SctMNieNUMxetcKJM54LPz0eU
vEuRL6H65t6f+4xvKQAdBX8Is+qeMgHaYP43WwUl6IRMSO9KMbpTkKv5alFIb3kduFqdK+EkRcWo
vNEwG7HGIPoej2ZGQzyrVWFJpx8m3Fkoa6eRdhBA2z5XmNQHXEZVpeW9yh+F8DQuIcVcIgZ8hhLa
MOPJsZwE6PjnPAyezBqYZtVzsW26/FsDJ44CvcC++N9FgA52JyDMXMBes4f2hW5CrwTWfOtvQ+1L
sg0MlGt22s/b3/LiGxUm3MsoeWCUJG3gh/eIZuUwr4L93DLlFZaDjYmuXGBcrD4GZpSiQNrdalqx
XTBzEJlutD93a8UU9oumLJniz9WjCTfjUF4HXzPJN0PJbZHChkY+X3F5tnsKr1ywV2JXKy9v0PTN
JkanbcuD31isc924ASRk0ntnUjjABuNBzaXSbVjhCU0utNmsjg+U02dR5zIvTQwaoRW5314JSOjM
tiN2m1TDTixmff/PMu4evQK/wuToCWloUHRw3arfaOfEOXTPNUyfQom4tZSMAM4pHg4Im9IYU3Jj
rm0MxrI+j4Boh9P4gmPaWOqi3m32W9mS/KgkGxWjvD41XMRzO1t1YzHqJBpmUQNZklmHTIN/332K
PKNH/8iggOJgoiNr4Ds43chzE3d3qUwMnUnH2DumMzdDoBTgpj1fejpD2G5WZUjqyEyEoliDUrbq
51IaMBeRCWkdGrhlFfZPEwWI7/i0BdvS4hUOnCWqx7fXGg2BdNNvo4XVRQ9VYvqeBm2l3s3wyza1
Yid8w4lbB9i2dX/MUZiSaFw8vtHkeaoO1QncWVuz54IUPky7iqyFHZ6SEAS11Ftlm5snz8jpsAxK
Qj/gcXCwUlJ9TFnzdgLS7GzWaLO61NwnMSM81FIkSllqgXhdlRehQtemoqqonDjvk4R8QQBq2lB2
Jd3+SLLfs92fZfZ6A5PxbH8VppY9548Aao8ibppN/mi2lfu/WAK5Jl+Fjk+U4UL8fAqfGXUDd+35
sZuebqOmaYktlfH+EabEC8p5RWzr2BHsTUPuxVDba9+4AqUeMPh7pAOzr8SHSOZj8bI/6VJm/xBz
cbVyMB2N13sjMUqXC2PW4LXgG71iFAq1t5gLs0RCOIsJ0AwEcGn16uOxQpJurZfaXqupCsx1+UDI
uMRGcSqayZImg3UjEMk4achndlpBEXKJW/dL4TIrN+osim6trlx+GoPeJKmQ7isiWwMc+ASXl5CT
YEVetEAfWoyWH3iYfBwVUIpqnBslGCHrC9QBE528iX9tPnI2EtyCpJuM7KpYvKQ7uK4KUdUxVJA0
0RK2l4DW9OBjRSb/ujVc+JqMyPLUZqNYEi4HKimajros6o4RpgcYpQy9Hv+P41LARY6FvowGefXL
IC3Th3nk6pkqphy+msXjEeAIB0RUHceZEbg0RW+HLbWmzwOjgEBrRoBef7vnhUhh9BUrZEUBTYsK
cCsYWWsrGaky0oS1SLNznv4jqV2jyZXIshJ8kxDdFEs6fuicMzavdJvjhpqyUUYW5knO7/mlwG7X
rq/uHzdv1NSxW9j0y0zGft1+dm2OTO5Dxxr82BX11F5Ls6bMsbtoVeqoUF7K3bOytmP+pNLbu8Ky
GkofNfpLGk25kOtrpQD8YkKnTEn2pLanVovo4WeJJ1MP7CvuhWtjTB1sDQCvMjCMZASMrWSCr4ja
ut19Xgkhfqf1DmM3rHbDNFBvNKpMj8GP+b/xdcvMJtBA5HWP3svtCqEfSxRr6VP61obERZFlWzwB
sbvjkizKcomrDLKT38E+2pdw8rk+yKpfo9dkzTeQdM/BmIX/W931U2tJalUVU9zT64upunhNLBgb
oZ85d/HymC94+mgLl9eT8BH2IrQe1F2QWEnXN4IMWsSdMQs46kuFF7FzKhVp9pyLRLytBUkDNqpc
6h2gYbz+vpaavmLLcdC8/RHYoEm9NpKcfjvYPfpcS5M4kg6IkM0/wKR8GhPzv9XC33HmdYrRTzXV
TZGqfypDaX/mkw2QtgDLVygvQUXtmJ/64OjLDhNhAnzVrD2DZPpBE/Z4RVXqIIqsy/yZ8N/RxDYL
peOR+Nad1n2NGySEvmYpcdrqC/9JgEr1KJWksqEdc2P7LjEjUYnJDF50vOyIu6jQbyaKo1v3IB/a
m8r6o+3EGPVrxydtHqvuTE5DsSNIml6mfunI22kj9UkP5lBKkZeJrsWj7794Vmq+wDQB/eB03Lc0
d1fbCuULPJ0ArrYw5d37Rf/3LMAoPC+XCyDoJIe9zYAM1ckjicX4ii3+ba1XWgvIs4hchDkgwYrw
gHTzBTWNU5fHdxnrr9XM71OvTJvHNH33ykAnNbnWPdbRnEyBZ0uFo5SosyqKAalRFHEU5IV1Lx2S
gJoZXXb7SRSDWqHb3VjyKPi2GYw8vgN1V/x9jBGewIYSL9EPdN3KWHK1Dq6EWYZxhGE21C5TPn8E
TiWPY71PcdAWNlvEgeKdceJEv2Qe+IPGE+NL9BLzi4VhGY5ron27ODNXeeVFODtCw2WShtwFnTOG
z3gZ2pgXORq+708onAr3HgA7DTI6cF/Dnvy8O8ofU00zPwc257eJFBB/vjhBCPChG1f+2BWcOcdQ
XeFySrltMAbxl5ohaeN18Ml3Ga1ZYJqrif8UbGEcI8++okr4M6pip/Agw4eIR65TvA9xFuJf6Yco
uqb8dvOrIzIFuckIHVHQkRmH9xiTFL/cLFwd2aJ5IlKDIMxdeZPM+hKqJSKJA+PUmsQDS1D+6Uq5
Rl2RXD7vHUqMaWLy+Lc6T5rOk7uLn8t/SVk0T39RXk7qoIcH4m6ziBjl/QJc/wRiGfBvYp0RbHoC
kZc7jMWBB5KleAUFxoF3JdJN0Bnm17/564drTyQPPf1TO0jlp4ny2c8Ah109KqiZBqzZAvuwUOoM
5i39x5zKzvOiGsfUrnagTLf4jAYrRsuB7fv+1ttxrZRioVg6vTEahyKRDPnHq9OXJNolGCvIUKHU
8n3nw47FjF7Qn1ewLgzDGihRnu4tk2GWTZEMjjM5vJ+IWyBj9TOM3cP2RukAiUqHwtI80lgFx3SD
OeK0cHJrYHFNbuG4P8SVpviHAd69S33Nmvh+8nf21hDuflUPdwfQ9EetmZdkOtYqjbnwUrzu0l1U
tdRPw2SOW27JGO28y+jeh4R8Mf49QaguEwU5pPll8e3+GRlN5T4QFLtSaWSQqjl85CzmgeGgS2gv
qtAC9YMkP0Ufrb6jQkIhrGvz2EHuwYKueYwreHTdPXxmevWv+SYZMTeM4yUMZQ5G9kdZdnx6mqBo
NYdwxp3aQBPbpmprqrhbHydr4uSy0nRxOrCag8d7DmCj1EjlD8PvyV33PNtTP56vpSTWhviMS0xK
j2oHmEfy29LtVMbcwndsgytcISdQeLu12J9SW6MF0sW6MMKaoOgD5NF2jICAg1Fgmmg4Ygcha00a
EcvynEHKLKsBTLMQkK2bpTmQU5gYUlzCXq4PIfUYujlAsPXHf/CMq/R5cU3yM03byWOky/SCvRWt
CReH5K2omX7OTL0Y+s4cr54Mx4WfmZOi5+Qu+S8YBoJFgUdE1QHKAbeqAd/CFc8oTsReOZ3z0+fA
Wz/zH9gduAneHVKSMWvXswexR8JHQQOqVaqaqJY/+fwdRUFC2FJmd/HoEYlxiXnR88iFM/Qc+OCX
+pVyZ5Vz7r/JZBl42IQP5XL9LfExwM9a6uWKrBOC00mtm6Nc3Qap34KeKz1iPehhDDH8xVxEgyim
+VAdaxmlKIyQIZgPJPvyBiYFZAQeokhlycMpzOtGE6VYeFcdVQ37n2gr8INEpOz0axM74IfsH7B+
6XBsYql9+sYbptJqGIdn5Nh0gB8BX+Khgmm6VZm+YdEaFiT5LdXYc5WgOMrZ7Rv2bQ17f1dCFEm+
rc8hNBWZtlWGJaUY7uveb3Q8oeUMqK7MyXoXuz7ZCMgersA66fPnGhG9fUuIBx5XgPz7dzXcKbbw
FBL3aKiPOdt4VRu7zfCL1RrI8zcpjdJ/NNxgQa0COkKW7Quc3neA6EgpCAKxn9tiF5jtpgQ2Ns+G
KkHlVr6n8uJCaAMP0IFHQtldbrC4AvMgVTv+mKBhvNOP8epE/VY4to4WMdAFoKZPLWXyH2wRN7ps
XNU3AgkG9ngokPzMoIjaCGPEwF0ezPFUDhdHSaxcXUG3MFmQknIdJo/Vi9AWXWXUJgmgTlLg24c+
/1veaRe2vTqLrDcJ/pHv1jk9pZGwLGegRQ9O8Be9VU4hMbSZnAsNDb/aiM/GTauRHFkK0oLvjE2A
En9xenyQoHddaI/VANCQ1KjrL9guLkEMJzJZfuPfn225ouIRYTXWCDpqprj5rZZF9EaxIJ6PSCn6
HUWuu61iJXLtVyLW53z0ePk15A8yuxn4Ix38A8oBUlAlA70WUhnSDdd3lscg+0AQSwjLsk4rWYhp
RKH0jOmv7bJ1u1e4OpVrWMw0Ua4DUQlCQRUo7VgbOQfdYm4qFe3ebSxXMLnxt6Ic7vZhnlXCPQFR
h5B+dqzJxSXd5g1z4xq3GmHoZq3Ypsvxz9ZTDibOTxQrYXDl9xx9A8j3JmAePeyoWuzpJxU4qz2Y
6s6Ujd52Ef+2yvxHLAutYCCiqAFALyUyz2/RwfTg0E67iB//pKlf8VL5Uw96nQOTH6yVBJ0GcNz1
lIyPDaojjgX+AWUwHSEtl/Ab8guJg+xTcnjm5P6QkCLR1A5P2YWgD8mfcmfx+gIlAnHMZTI2euRY
JErpdNuKL1wVt3NCgVjc61/aqhCdrEnJKq0yTLC7oQHW8BGI98GGl9/U2ZsTUg/DbbJD5y9NeMQl
/a7YjXXOrd3EDUzlLL+mZPRbfd1gZiEH9fkqjJ20Ytd3E+IASzMdLJZgeE2M+bMbMYZhJSzgrNHM
tGSTnufG7f+e9mtwJIwUnWGBqrwhLcVk+UIbiDs4jXSVuN0eOUeKhHQgS4wuxb4B8Eb4OmhVFYF7
3nJAY4wt/kWPuw8iQsCsAmOlDKE0KlqU3Lx0XgMlwOdzIGgIiRKimKxSegXyJvahp2vx+WWkW8hS
MiAktf4KByKY9UMH/vTHo1IfoaIUsntXNEIcT3wGzv5wLZThfFbV6G0VEtKEB+IvA3WElZxVzROD
PBaMUMHDvSC08ecs9gkYH9gHf1Ki5LRfwKAgX8glppW4q8QDIvmeqkEAAdcDFCvc+cZcssLrdzG3
5y58QwTuWKzKxfmuwmY2deI9Sq/jdYm93veKbWdyWkCSBgmavCK6O5TkHOmsUUVx+ROnBzoTbaiw
4FuuB3f6n1+pdIUN0VrPmVvwL2qGgGEuroQFhkBP72RBwOtHeWWad4TpeDtHOCfhDmwhDsUIUbDL
6B5h9tIc5faYHcNATlkt2uC93onoccFhM4U07J0npY/ZXgSLguuSTiDg43ej6TdB2W41zfHxwlJH
xbk6E3aW/vd8olYGSSyoFpqmPa3xvZWkv38nGVJXTq58G7mIVzos7K+usfpANOA8Gi2rOu/4ONv1
fERbBXN7toSkarDwNlauCKGbwu45Q3BKclZRRUdIz/7JAxVqik51ht1VXjHB0a3FybxjzZI0ucfV
sW+KLvHd/vovwPrQYfTcowRo3ko63TgOJcrBdH0aWWJ9tsv2/WRrUFGMjxIHE+plEajTMF89mn68
ETmBWiZZLSryduCYFsjBw/SWD5IxGfhtNabPlfMBsJkatV1RgGbuBmA+4WRATQ+3DD+RxfCRkdL+
E1RhfxxDLVVnfYN0HL8DGc774knJWgKY7kjce2qcNVv4K4MusjdM5lpAXN67U3yP/mCMkkHXdhUB
Vw/qjO+TBk8oXVmNVmGKbozV6TACniuQMbXk8u2gSccjcaMgqOj7W1DYJEZ/grI8MdfE2nUd7BkP
tBCF6NMf12Zv561hqaHCeizQCc90GH2rBzZwdb9yUKKblzcUnNY5fZK9xF/HpYEFZCPlGOLPltX4
LqQhTNqlNKxzX5l+O5+AbtpvdUCALE5W3aqY1gOgeeHgwHFB3kDtxRlWxee/PpFKac/P9By/B6od
RTyoEIrxT1ZBWKBuzcLt/A39n4hrJ+jjueAyxDrBpDNFyT20G4a+8klzA4ta1AKAA5ydqw0fczFr
zOL1ee+0e+p02k59lPoVV8nqlbNPCBPHb3vZAMia2mXdooyzV9YMHpMET8ytc6vi8Cew+SjdqW9j
M5tIgabhlibz9e9bmEhswjKEzd452OyLJdAoiZbb8/hdpFYB5GsTc+F0ug7oXrzNv/MSVRTaqTtv
d9CSxfcWcNBl/XaNMZGtvyL7jHAQyCVoFodhQlJaj5kddeLDxg/OVwrpVmB23ahK/l0ccIHykujM
sDs8k1tnKw9bkPAY5jC9CmqfD/pRre+4wMu+nhd0wHoHOmuGLEkR+N9YE/ot+bIYCYS8U4ZZCL9Y
FYd2fbDejCQtZ2VR7DycdY4bsQ3UUYn/CSd1VGCHo81SPKOgjJCPPi3O8M522aJri8Kw/azm/TnQ
3XSlHIWfJsO1JxAkLoZKSHQKqJ3OaQxXbhcG2C0CDTiQ1paVj0/vbaNzNraYuKSTGKgHzlNS55ic
hRHBSjS3JKF/C3+yZaW2XdULhBU1oiyCglQqtEev2Vpn3B4RIkuOWmqgr8LoTZIVPtcnsYL3kBpv
pZ/0OOJg1nZ1dsXIWLad+1RoZ5PtPDw978AwPAR1b535dO9RS/VVls48Dnk6gxhGbcA2pNhUJaM6
k7K5I3EmiqIbzv767/uvAk8fHZobVckbYR6t1gUOY8MRt3IGkFPfoDIaYvFvkjDLI8dRZXaZsCSN
uQ3gOeXzZzR1T2sM5Sa4bhfJCTvakpsVODvJ6gbEuCWmaVUgbNw1ao+Z1Vd2Psa19NW05oanuglT
9PlKfzFk3RRYNTiZnEH9XO3kFdxcVJngDWAzfu23ONbpKcxjyh7x35xnnT4fpqc5S1H+0qy4jC7Q
z7cRqijiPXwxibtxWcacKz2FTm6ghlLIQ7pRreOE7IZx0AoRwK9Ie5CUgzNLdFUqqfQF5P8Y9QkY
jCqd1SE9U5v1GZExEId0ToEcuhX51PuO40HBAEmAnwusYoULbPcJ5tjIY4I6KsxqL7ZSa0hKp8v5
blxvIAFJ05hECtu9f6qz2FkPCOP0eyPb6KskbDqXhofih8etRQvoVWKSwHd1NHVsEuEdwpItyc/Z
5cyLzeKwte3FXsuHriz9GWz+3OhCR/uCMzDnqhV5drgJNYO/t19+7OAII5NQbq4/L1fCOw6LVhSS
lasG2qi/S8jROOz0Fmq5gyLVVrd/LApLPDvNBiPCawG0efFJqilADo2ZMD7Ad3sx1xwCH4nnECCW
wSrq0VLKnNtLsH3RVgIfH8HPOgzubg1S81XFsVpccs310DvKZjwNd4g0OQ+fJlC3sB4fWo982El/
kS1S6twutNzt2lbNKv+eszQb8oD6U3Werigu8soKPftQPWxbqxw/hptjpPOko4bVmtBpvDjAw7GD
qKDHQ5TGJSvJevmnhLAtEs18nfiUboJZgnvyrfUP+I4gm96pAZNYlLDhVZ/Mh8E7swznESrEcZ3y
EM4BtldG/EfTz3CNASQiCgn8a/1/zDqJFzh2rgDTI6IiYPYHDAZRd5lLQYwds/gprEj4Ax8uxTI+
WJDTVsfBupHzHIUJMurkgksxIrsVOEHcm6eoPJRZoHyK9LJbiN4v6x/sk5mc0Q0CIEjiz6TOPeZz
OWp/EzYNlaLwaSAGqRMQlG/P5UeSOYVNZKDXxeXVfGFE41O04fYec1cvlawsJ6lV1f7oLbKWyeGX
zCH0OXew7SwNzkFoOZ2x88XpkC48E8GxBJ9P1iTQB1Gqa5WUd8uXzsSqdiQYvsrUBYx+1/FhhIa+
lqrV/b6cN0hhlyxM2jDY8+qeHdPD0PRs6rpWUeUmkhohhfMsc1Cjf9WFtIh2igcDNJScqTKo1pl+
VFixsRG4tBWYuiYaSTtQVcGNFJTHYMrPKGaT7mPxp95DpgxqMDU57767mQ6VNY3tOKTVVWvRQc7w
+SeU8M+XiSpC5YCUjYyfFUf8Rhpvk2cW6J8zjLJXBcA0H23B/HmdolUwF1b4nuIgZPu0BZH+EQUG
AJbNJxcCvfcFxeGrACni9ZFdSXz0WxVGKiWUqEy2CHXFQ12XyaNKObRoJGqBEeLWoTQt0kMIBDYo
7C6Gu6jho61/uBhsGvexaezRkLp9UcK88L4nZuaEeeK5+pVK+FKvjVD9goi2907glYcd1d4ytEQK
iKLAkDeydApjPRUD1NpUt2+VwNmxFGxZFqjbQVYdi05JFYnYQse8uOGQbo+vvE35HPSNSTCh1IFP
eHI1nh817hzaMdS9akurQXqkFpvTWrYQVYX00ELlFXr5RuB7xBOCnkJD33+1LKA1eATuwPpQfG2G
Pr74sp2sJgj4rbGmTxpANyNB9ZT+kuhzYBOzPsvwsMngwFgvth108e7GLs/+2xLWkw3WAcGb2eCZ
7H6WO5YW17D8R1RukR/nqxG/5Et1ECRN00O78l79yfe6e3TFl6gSDmz69C+YDUz7DMQu8cA74mS2
4vaACTHYFik3eFlk6cjZkPJOtlNFt6MxEESpjo7c7NGX94kKbexyul0VtoAqWPazrPWaIeZITeC+
a0mNs6oUPSOg6ELnz6ewPqlSMC2bMNInAeW7d5bG0yUYp3u7PlqFDsA95L75Oe8yk4CoZ+sEVtXr
8AyqA3Jb1pd70+fyWMRz7J42iARYHAUWcFHmbApcS0tE+7AWRYNKZrIiu45k5TBszIsrCieU1qD1
ZVXh0mM2lbmV4nEwTotuNK/PfBr+D+HHA5z4gIUf6p7+lcVN5YvUrV0S2dtoNbWw6Etf895yEzuS
r53MFJylfmqvvM7glr25+qKeUibJCi0FXL7PV55ulQEIun2v0To4LC8/sj1b1nLM6UWRYpp7I8jT
T5KinehdkyBsjWpdb8YIs7MIjxuKb4KydqmHSSPDtAjXf/AGWdib42MeeeIrpD7zv8YNXrTMAWa/
KxoijHNnYMW7UqhjCg5jQiW6xjH8iIWjPKY9R0NEspRf0Ltff73wwtx8O4r8uN6oftYQZQ7GBDNM
2zoH6rYS8qMdhUzsODj/rZ9pMCySvqgcfPRuyYn6/m4oLW7ZJ+iTfeHmUUCdx4ajmMkTOEdqX/yU
MHr7Ttqg9/oQ9MoNBbNTzv/sKtpc8KVg8PgBJvDr2pHSCy5/ARFe+SWMwuuRaLZTV2hpFxZGLPO6
+ngdSN912LWavIHDuWc+gpbr7jrNVWinFzMCyTAgOsmsgN5bfl9vBHGIXWDO0Xyh9S1DY3ivTWdI
fC6gRd5m1GBwrQ+hmvTNuFQ/eM/KpWi2acp694Br1QGdvz4nMYtvFuo6XDxkiQi0f3LtuQe9YY8j
/N+T9bs/F2F+XE39ggJSlOJA6Jb4TuMJxXjTCcmFJgdE5HugiWNVwdDqduFo+4mDC02w4I7ZeILH
v/Y4Wm5iieRMBJVw3iXkCtV1TlOBwlpuN6KKUnGtQ26B3UG+eha424y+cbGFgE9WrnSlOdYwJRnk
ofwjVjiCWQQWMOV/Ac+L+blCVCe3TbdJj48RX6Lu4qQn5xkXU0ydyM+5cRUoP0+D1pNCNs1P2Qi4
6H1uPzqlwzPpqezYVXByAZ0zmJ0geZofeyx8JW3h4//4VilLVO8C4QnbCCZ55+0xszv5vBBEep25
NCRRIvujAnFf7FkPaRJf8SYJIpqChjOLaEJGcla+2iW21hKT95bYCoqkPzTRL0p5jXgJtUFPibdJ
We2dfw2KNsYgdVQccDuHVHdj4ghLV1qYNpOY6rsQZvlxU1/ea8+xAyQskPOhyeccdIA/6ug0i4Ie
sO1rmTsYMGNOMyxLLqeBSOrkOSFBS69FUiVn9bhG6zWBcSiOF33sJOLwdjLVNBD9aDBTx36K1UVJ
rl44SMYcgtOFD36x1G12DqJp1xbQan+j+XG8EXYELYBVGicQZsrU+2/A0MvCAfS1kKM5F5WOKsAz
HmShnV5px2m/uj1ul9wA918BwCQJU6fKyC/M0KpSU+wzSTvYYAjpEpFoa0+blRnSyxgMC8gkLZd+
rU/aVay/P/wERYurFW4d/MZnwJfpjLh5g9CPQpkVSKl16vQmU9DKPXgVstpyBxYMjVukRlbxwDWU
ZHmH6mw1aJmaOtxIIHrSxxQE1wOJawdCeKiBmyHhG8EvjROkNMkHFJUce5B25Ra/4n231Yg46wad
jbKEi+OuSi7GfvR6Ny8L+eIFl4msfIjonEjBH/UuLD+taaMoxjiFermuWhjvUdZExWASAbbG/+9P
f82AK4ATelCjhkRf5VyLhCiM/0ViqNgnFbij64WyS9shRU/eyWn/y/6c7Ca56X+jYoFspOYXm/Ol
dt5Yj5BYmbxk1z0IIJUboixKYJEroOzvLWuHL6Y/3MbsiPy9/3NxN/OV/Au41DQoUOKvwtYnkaSZ
TCh3vvrr1CYd990KcL2L/T2nwMU1SSEnTmiX5ysA2xRDcjZIcOZdam+rL2JhlKdfG3EDidXfpQHT
7RGmr9v25a3hhpYrTObgJTFCLl6hTVej5vr+fAnALkJz+mWdl8nUjRRxNxox5q1gKijhPW5eRS1a
vMaTEkX9YpBW6FLBk8xzdC87ISEUICD9aUWUDUGM/h/1/O73I5xEKZGxmqD2Wh4cOBEFKp+dC8M2
LZr4maCDnBuJNGwI+bGjWUb8VWi+MjOEoSWVtJkGlksDy8qzjjeJhgjN0aG1vt8ZNnd4PlL+mUg0
Y6+YQB8vidF8Ly5VDtJNOGAdVMMIca85z8RWomc9/gExrbr8UfaMb0cPt79gYH4hb9zfl6yfYNJ5
NcmEDpCl1fTwdc/OPb2006GR9GHt3FDAGNLF0vRFe5AYWR5NGHZE4LS540luYlsr5eXt0UzhA1pB
OVS9c3GK/ZS0B/Y1zuUbLf2+xX2Z5F315AuwXTEDnVtqyE60fAdFyQxCj7oo7yss1hl2D3hZVRII
RPKLYhkqDCdN31PSRQgi09RheavOOJBgnCLOcrVc0vU7OGt/itPA51jTcgFvfncQ+8gQQKS7ZhNz
BVu9oTwp6qHP7rLW20ZTpLy4Pmh5IMmJmGXm2IUarqCnq1JXW42yig46t6eWh9wr63/mFrsRH6NW
n+qWMVU0LIj+bOu6Ea99z5mm/MLMoWU3gwBVqXkOjqvE/Y80MJlaZLMR0dv/zw+52WySiMxhOX36
ge+ynmIdb5jFStssaLq1YrQdJHNyXqZO3tHE2STbWRK4JpEsn08XaljiwtaLpXiOuKUOCbNdy3JT
Fu/AfK+1kOhNZ7g4cPvbnsJiSn/yEjIS4Vof5+t7iJ1tLtGEEZ7GZGdd5WTWICxCuX91TY85yNOH
kyd4/837v0Kx5pO6TrMaf1kn852ZQzZ5W3EU9fGl3LcPp44m5hWS69D6YJUK8n99m5a8eL9fCoR6
N+JAUDAksJ/DkriDPKfjvKclhlYHZTLNS7xjMF69Dtigd34yr/gq9wWGHBDXqXDpjEWPNosq2Xz4
ppDfLFz6ReLrv9baAT7sGdtR+jKFDilxI7Kdrsfx+JlCazOfS8nsSWMyZuhlpe5R0qgOlXGLIAJC
aGJEIbWcJdfDJQatdhAnyMj4h2XN0eyddGrMIFVjrjNcDsYG4MILKemO1//4NzimJJVH7ryCRhpz
nRL40+twW1Rl1vaKroRrsmkHoBa4DVbumnPamjxcJej+NOTUOaqWhoYJ09BUK23AsCVlGbPcAC0s
b9TerzJS0Wik+5NVZemdqKeKyEfKyD7R/aSOJU3hCtT5ozX7W19xySJRAF9JJ81VC9+HWr4LN/om
8nPOIXrMtNowKNZ4DibUwJnA6C8AkAxOQ6nX5FTcLYBWnIpZp4rb1/OWrHwoLdqXMIXbBk5BikYb
DJ6/bZIODm1NoqqGO9iiQ9V6XEMwvm1SDMOA3zpr/95LPTOENdLibxAlryCL7bRJbw99+/sCUVd2
47CSi1jZOVVakrdjhY1sdzFlwg+kc9UkYTjD0pFwxbyRkxI7jEhVl6e5cEAtQaqB081OtWHX55Ge
HSIAsOcMgo+hBQDexL5HEaaRcZO2BFWzh9l8CBLza7rnJSDh3j7cthBfPKuzwDc4WSuRX3XdrWLW
toTlutZPIWWqKWr73PszE3MdodIZqbquyjOElEElamRzFl2/cKyMH+2/FPHUU66pEEog/3K2y+Jd
qM4g2s/804ePbNaaUwZDVmUmbU/gFX+RPMfj0CwjSIJEQ6kGemAbZ8sJH43osm01I59ZGhLBvw2T
gqbPToKLZlYNWprBNjW3gUlxvY01Tv4wT6FcGcc+9IijWIr1qMfzdo+fUrIUVA813xht/kLDN5H8
obBHiePNWk0TqRrSAIhTddu+NJl1YZunhCZefrQp1/BBpMlLL3gowv+GStWo19Her3kHWVt1S7t9
ynBZ9v53hPrAE//AL7s3Ywcsb8JTNp7Rttf+HT5ANzfZnzVLAWdfG+9iWN+hvGVfrgDkAshxrtvJ
uGuQRzEXlLOR5TMd0foupYOWdwJpQuXltXFchRzJL8YMNXxE3TEzmnYhnouBZratDmUCOXurOEpp
5CiwNT3gjps6xI8RNh9cw1w3pvK47ELe5+CWfZFBRs39xl9Zjn67sMCSNkwU2whdjiflm9v52Tbt
Mvh/m9UhYI74HPDkukXDMs+C/OOQvNpMT/VdOinlplLWrxxzbe3UTBwRBU/QoDd9ieQ9bGUakWEJ
bdvfHClB14XEe+8z4/fLZh1rMjktuZ5rOf9TIK3fTUsau0Wuz7KBNuNVZWe/fmdZn1nvn2lmNqDG
1JHsjrhO1XHMkUvKuAARUinh2PmDsn6uPANB4fSCAB2fKZsq1puVAg+XpMp/Obgh3dct3SmmQRqI
vifcrgSvel+MpUrm64cTni2AgR9P2miogczLRZAgcqowoCo0DDUtCAt8YMvgjyCVbfQ4e7vS5DUU
pNPSPK1GUjpsAP9XbRfOVf6JzbF6cmHrj8CaNUg2bq6ikijsfqTDaxDibqO7hEbHosMfEq1hRgqi
M6xP0VR0jl63xQgDJseuBcalurKJYm88uUW+8yuVickSvbDdjWxI2VKT7nCXi2nS7Rdc7Q4HjaiF
rOicROu1TgFqQSGpegpFccfy+QpV5MN4f9eHfZQ/o5ngSm8mnJLI6sR9IN5aTLy9I/A/uBULP91+
4t+slNn7WCzXS3DbCIXHa8v3arbffKnf2XARrodq9+fc7dEnmVS59gMyJURCKndLJxD9c2kNncCS
ah8mG8U5pfjhCNQJ7IA/ATJohK7RFLthAXEo4K209/hieYHxGOgwy9ROqvKVM17Lvb/pKdbLGUfu
lYKJJllhdbizbIlHJDwJsyo+Q/Opi6Vng/luGcy8UU50N7LrpMSTneRNPYm0Lb7sUg2GRSCpnC1f
nezZNrITgXxvxfIOhZcwSvK9p7tZJxDnaWQ4RT8oaOOEIikHhormBClrFcBNFIjWIPYxkFbfJv7c
Zt46rV5a1H0gAkK0sg6PhxNnTqXSPIQahbZAy0kbwAJaTCkRXMh+09sDUWHzK04txZHJFuw6JUk4
Ac010hyVbpnRe533gCzt1UKVNlA6UfhRSOxlWRM4yo1m7dj5M9uxORHIV9a4Xz1VvHAzHUz4UxGE
vfx/2o61JeRYlRZCCBrlv2c4vmkYJYcjcKRoPNJz+kZFvAlzgo2dvQmmBZIy7r8tZ7MNbvZYOaRR
X4pDfcly7M33Yt6bqg9EXoDmIawu9GSyqBSYh1fOZ4WUVKdSaVdVFh7J4fTBrS/wup/7CgkD8gGu
n8o0l15/kiieT39c41SapCdY8/74POpvjpZsPkjBtrJyg1QC03j6ctrJr1kAXgws71H+fdvTRqR3
uJ8ZgQpZOE0wl2Hmbxo8dRtbpIsu5PrUlmSMDBoyvjXAgOULMoBxNBMdCTMifSNaX399oheVlB1t
2T8aAGSpHgl4AmbBdYGUzmYS/Y+IDrtjON4Yot0jDPZqRhT4UwrzKWhEKOagDYrNAfJuEq24yI2+
LYqMUBr0vMV2XjWusvcu41Q8ydD+A/+oGHUvGKLteIggr1KTUnogUmBZwhlXreg0Wfb/s2WBRwtP
MR6ArgLhXQx/rF4KVGwPPMSFJ6QcSlT86XwhTnLOy7X7OO2vCx7gcEv7cF4y/cC9btBYyJzmu1jW
HHNMoDz0SYlcSCrmSgwr0rOQVs3XVAIR8ff4MROfA9QR87wSxi63Y38xtlvIQAIQcO/2btMxnoFv
vC6hrsXSATq+4Fuzj6Hb/N7knmTjInrrZVxobUI9txthl9Jy6I8jFC/Qt2JrNi2sF3qjH4H3TLI3
rIVH7xSKw4i4wpShIM1kFpxRXCKz2Xi1uu0Mi4aLuIdIT7ZiNwQXWfwEqPq6J+IEg4bnAwrEUxE3
/bUhpYfXblWViztPVG5iVcT4FIDIek8M046izA+9Wr9SvNWTyroHpX+NXF/Eg3oQgyn5wA7ZoUeu
g9eDve6lwxtpI8O8Q6DrUAlLD4bAOZHnX2EZWMuwc+o5sDMnkyboWiy2ioZlj+5xh4wFPjgQayxG
yrUnJSnYBF8UKstxKvppnHChvnrkkKvid4BzpUKINmD/hjsAVXn6HSnR+RcljjD7qzLUKTLpCTUz
ujgmomnz+4rH7xFrWNZGJ+nBSkxD4EIYwqpjssNl8QKcXpE3FAUp0XGdyoeLuWWqtSO562qiioHA
/rYddS3exXsuBHjl4eLqX/MJo7mSEXq6KGX5hxnw498wh/L7v5t5nNGED7q3ozXoRxbb6PA2bPLw
vxswWMMUULBSzXQGUTCjoLfzzppAbdTRsbXN7F+6CZCOz4DLQ7ibY3C6L+uFWPEpAcOM/j2t6z0D
63xLiWpDi6jqt9+wGKfQfFcj77mz3QrVQZ6ToD2Pxi+09y8+ANy622KvO7tP/5ovGY34AHOXdz9L
HdLy9EhS7GmlExpETqIyF5wBB4hiX1UQ7mB/TqVLcfgmrhh/fodqNEoD/GEvQxjPJkz2N8RKMQU9
KjHNvXkLwmgWQ8nmclvkBqjOs+exL+OZTjnyq9sR5G6Vy424EwsJLm1274Wyn/16aK6zGdkfF2Fx
p1Nk0LJdd2woHAOcrMYo9EcvwdTqfHvFLMzea+z/22vJ5972JU1STBTAMvK+LuJrIPyUUEjItmgU
uPhKK7GSWdtNLys0CuNWjq+sJ1JQioDdy/CkZeXoG+8wu0JOsb64m9JT4NG9blLPk3OmopMm9S6L
mPByNqVOl+s1JQbO8KQutPoLu8yJ5B+sWndWa8qhGH/3OTa6TUNmsV4AV13bC10UyzmepnoSSzrO
2HSh9lDrA4fWebUbms/BXuB8N7k8kzs04RQdek/OM7h3t4uqwku1DCUaKVzCDsHYodJ4BVZJyBwK
a0XQd1zDsUf4FbTIukJBhZCP7dbkA0Bd8ynAOYuDu0CKhj1i5d4qwjedkK6j9gNtcAuzxWOA0xvs
msXSeK1/2q2hLNNA/BaApyD7E6qD5kkTwAI/ueaNEYUUnNMfDVvYSpdmcfAsdJ6Zuf2Bjmx2qMLb
m24RKiqV8aJudMtlU8scPVmvQCgs8ms6B8wxdPA3p25R9nZrSo4T/z8Gg0IrW1gum5WApGs8lxhg
nmilmhuSe538Fkw4DM9E8IfSA5tSSEV3U+FQsYYuHx8tqcb36BeF8rnHlJOgy6bZ033wx6glpHU6
DmILjwmkJrH21d5D2yZsV8FYsTpZwN8w9FtlWAszOENjcqDjFHwLtGrFm8XG8fd1M76IYIOxlpeH
2GqmwnFEKxmcI3KPdmxPR7PgkvYEwKGZhZ3bgzADbvRwgvhl67zz/NoRTROqujfBGYF1CayIXTyW
MFZS4D//+NpITejCINLl+S0gaKu7qzWDOSBtcpPDZxSQ14l56NPq2PAqmeBAs8ALRLmEhkORCtlv
1dQtyIskT+Swmb3NRJQuZrtLHv9X3inRJ12GxtFdFcJe9RsfyR3AwK8E+Ci5e32yoVU6R/gmh3Xq
7NQH2mnxQjjxo/05+sQ/8mzpCMZ4PQrotf1zF8bOH8g12i+byz2MGqHLwxTLbR7698ghdhz3KrlM
GIMr3OdEoWPHqx36h1PdzVs175Bw6EYJ2L+ySoRCPRwYM9u0qTFrbdG1QLBX98AUi7AZRa5BOaue
nxafz2ur2YRLjb/25k7VH1hhXNDrV8KLv1rDZWPEsuFUz1318N6Cci10PBNP8vpwogleKKPDhdE+
oDn/CXGlCQtKslSsFcka0OfoqUq0n2mCutwili2dOoXItAfaTtZM6jvlsK47n9mx5bVgcGAdPBLk
Xs9CHyAtG0/XuwUVE9FbX0jVSYbRPmgmcJsluXgChaaudz9rdiBEj4bAWyuzNFitIvA0wYuLh0nr
0DSn/gE1t+qbrIpz14jFFitwHLKR+csAlFHPDdjp3/YMdnXkFeQ0yARMEzuLLedDgOpR4ASdYtvx
4tdR4j5qs8Trw6n4qV4Pcr0mBc7tKDoxrTSulWGwUHCf1YejC/bfOCE6TMKqyQdWsiSomgJHyBwu
dq6/nEB8E0tZ4+mbtMgnTMVExOy/K2fLHyVzb4fzDf4d+Busa2yhDo2MnyGMlX4j8DrBMV9ZjHjF
JgPQOmAwE0ZqTM5nfMzR0MNponFrYXAXIMTC+eNpgldpNOpFZS10q5tydkANgbpJMylN/CqW2cLX
q0y5FNtMCuiatI6NhdT7eddV0oSGUr+k89adnAXbO2NlbznHJtn5Pw/VxXRZufPvRmMkECeI4I+B
o7SPG+nf4+niVgMkZJO7CEOIf8C0L63+b4g1bLSoyjU1mvGFYL9BUhMEUGfj82erJFPgyek4Cfmb
M1B8uTB/Pli15RuC/EXFrJQDbFwOSSHy0E8yIEkwYU3TBre3h1TeDEb4yhaD0jHGi6/54v7pUfzW
UmNpckgj1BjVoAQot5DWvscivRxsyEbQjm0WF6nc9wqJt/sQ4bsg6tNP5/QVnqeI+QnMRz0l0Ewt
yNQx12YY72YbsNNtrfu4h6/GwyX/sKSfTbjMe3SiR+57v44+xYr7a7C3yyHOPIANWOeaGom1Fpen
TIiG6BDT5p5oVH1kR0SwLT2x6/xKc/TvBIo+79Jx+8vYpCgOmsRzXwczW9zIyl+eWqfRJ4ORzRay
RvAH9Q/AWknAmXp1APIWyEPYaODow3zMn4O7kjauyK3Hc7b46b3NTvhJYVGPebEmfbjL4ECxpgvF
g6CATiwYfkQJxFQk8j1jVQePnyL40cl3pZtiXRrLCZYrisHkZ0ua03y/16Uje2b2tJ9QVsaa/gBt
4Dtfk4XnUPUd28sdUpXpf08Hu1tEm0KyLOb9ctaq8QwyVdKhpmqMkv+DMl0tmwpltsnlySQHlpWu
+qAmhvkRQLN1lkMAHLgjOLYjQtlW2Kae+j1y07sRYfgY23hLpjWUF/Nz7erZCsmBFcepYESb8vWk
IYwpffB/ZmFeoLe0dyBZat0Mn18P2THDGo0JmiwAi5SazuHNi+U3Yj3iC8wknFrw/Pjt8dNqKpsy
iY0BbvSXgeQFiNjV/0je/SB7dWjfTLZmkjX1vdjXlHlqxznAVTv9RrDt2QlTuslVyzdgte85k54l
OxX3VB/U4hcqilA7mofoPtZ/YV/phthQksEjlrbpV1kQmm959B+568O6AC+pEdro26JhKM8MBsbX
fYPuKJ+KWNtNHtSjrb2reAAnl5yKWHyQhUbcirMUJ4RDpu6XJAZZ3aTivjuJFymnqb+tMnp+TO0N
ZY9EabFa0sXtDE7kd1UueJC3ETvgOeXPzo5snPwkhyiODI1bPE3zDH07n4m6O0snQN+fjZqAhOfa
gI3YG3yosWjIEZjIGoz9WvC8BRZ+1NGwXRaFbJ6933tWAn8I4wg8AcvxIJFscEBaUtfgTDLixxdF
obZH5LLog1uJn3NVesRID/h8uQLyEHtK0DWYT0oAFlT3S4KC9clAU9cPsYmmH9eBYjG1vI0iFD38
DJ7FKBSLz7y2yAO/9L6mxHYvS4zMPFSf//thSiT2iTQST/3MDRMeYDEMVWNpWRqUunHfoR12sV8x
bAYpsZBetO3+p+spVMPICZRcxw+KIDGr+fFddjMv/drs4xy9xxLbGT9GRm8YCBXgEPX7IcfiaNLp
nHJUwiPKjE1GNIDTZg6JDysyGeIZKrAKqXJMqoHtQnb8IPAO1StFtoDR61dROUBsUTx9+tOIvaws
/txuKaKyKDm7fdFMDfOs9IK8ij1lCUf1iMpquo6zEj/ZmgkpMCOMFn4Lz4WacPTl2cx+5ik8ZZGf
CaeaBzD5Jo0fbpv8/aMi6zNnm1+3AZo7oCvtv+FJeMgT4cI645WhK3X+17u6QmyEwPKwJtNMy1r7
bhhz/ZZIulEai0Y4xHXjBMn8pczrdmP+mCWnjhRQ/7qVLYXK+Xy/3NymbQh895RM1LQ3z9iRNh7P
weW4smTVpT0HRRX9Wx74c5+3KTEHIN2osKbrUTUB1GXW7Oo218nkPn80OH5KAkBg1o5CvjwkOEWv
SCU8XiC/1KphQDdKhWTLxN6M7JYoZZt95SeqJLfi2xHmIQbUOvptooaST78KVkOAwuAsx85OuZPi
d7dwxyRlPWIekSNLvEiRxmomMUyi/bnRuAfhxAzS+19G6Xwv07/72iZMaBdccCu6q7KCdu7OieVe
2Xtw2Y0k6zGX9LVEv6DJcdmIUzHEOXqV4wM7ng6gY7dV24FeacCRAPENHzT+ihkSqHl2oATTjeq2
KipyyqTLs24QMeKu5YbIcgRiA6zTp1QFN+nec727jqvAVYovZL035Fs0mcrdEumMNjHbC4Ig++XN
vOwlBKfQxQWj76SMBS7FQM1HFh2p97xlrrk+7TSdrDU3iKoDUtsNuy9WaOAjmC2TH14us72nRbjp
0S2gYGGBlpA+n0kh9G71c+vLy6aDkoH2dlwIcDF6jDIQmhL51fT63uVWCKhuxQQnGJNpk6kbhgdj
ycfOCfADH/mgln2sABFSdhl8jfCOUnlMeXkcEKjH+woEDgZMu+0Zxp9xMaTy1sCFal8Ui14dMpA+
gXREIrzyNy9jpIxiKOCpFtOwZymcnmc5YFXcGXuVIS97KWEUbZtRnZzORahxtC6Lx3CA+Tg1UbIB
Q5GnSDVEmssbz3GiXEBhWWuTlOhWAVElJ5swT/LVp8uomspXdoDOCSt/SgWGT2vkLF+0BEvIaoyp
avICKRhNekCwH6NYe3qLLMP/4L8HyzsMnxKn+vP6edrQFM623mvaqjE/KIzHteQ8qgmJ0VftGA3a
YHioLoinvdkZKg/Vz7U1vzgGtWRxKOSYcOPUNMr233I6PnvZ0dyW9CEpMFvkbWvImB6SsYPx3cpK
4VCcHIPUxP43OGqxinkTczykN26q7+y+gx2WNWPBliUZLAYdIRTpj5Cf1YzITtCc94gT3/zGtO2y
ZZ12Wg2vYRjPobWxY+YxmuTMUznsTIzKLx+Ehufzlr4C7hTdikvxmfqk9HRFCujr+7ZlaOywSH3+
ZLgbbk+Dq6l12zXaFHB8JzskaPNvhZXuvoLMcrxPgeYg4gywZ/oIj9/ZBiFjg97HpqjAh/JdMdyo
UO6xblfdu0rCi3kPRaK2oNwQArNpXqakJ8VkbhOEaZFaBgww15toGLoZTHNIc+L6oYIwuHT6/F+f
+2DIRRjIRO99ML3kI5rTz6jYeAq/NS8hcR944oHZ0+/3lyLkpaGRm9dN7QLTRgnPVzopRa4dmgjk
CJm3zrfX9L7UNViwH7m2XhL0gIXP3F7l3SWQZcZ7FZz1/tm9BNveGH1jz6pkMBXgtiYLTPuvFspu
3udEEawfaz+XL+/W2pCFn8cLxKzedLKNxJe3dGgyNyqAL+mvB0pl//FYEtltoItOe2WRLIZkeXQA
cK3ODyNZR85yVIf/V6Siy8z1XX6uh3XIcUGav8KxIpxYQLVnpHVi9kRMrKzyBO8d2e/P4KVjXheY
rRWOcN9gY/w7zFdCcSOh+IjS9X0OixN0lb3g+9HVtMqD1XPOJsMrfDkD+BZOlHoMLHy8DLOKh0JR
vBaV8MkRMehtC5qtTdiSzNaBV0AMYqK9TgSnZ46JmSXzPTscS4NsfKQYWzsfb1+nfrL6TvUOuSy4
llSDIJyhqoUuDSjltyCYpBq7KQ4sxHGzQ8UlUJbkDshnoAPRuzwkwIwsljHCixRLHTMjYqbl22Lo
IXe91mM7GWmOyY3PZzE37L7vghgKypD5UZipMhhZpqTopXeOSbLaQ2YS9XIisgL/h7hbZH2iDv0A
LVGKzIfNgdaYp9GCZ2CgkHLqugp3syvuDxODkD3lHS1Gg8pK8cSqV7tec0EhQRzYWxeq//2u91cx
ToRFu5AdKWxf4Wks1nDfSwaz8N91abet3SLPFQuC6pfYrOEYt4p5BIGxpirAELMrGOPlvJmZ9I0j
I8Tzzc5/KebhjZ/x/b/wRoxqGwv6EnDI+dJl9hiu2XQMVTfocpmtW/UyGM0rL05WTzUA6ajnMtTG
UwpZDqTFJFxWoYuMODoqviihLrDROf6O1F98Srby/lhW8EfKGTNBEvoPMs2XxoNjkM5IT2b6UG/F
eOMzR9V2nftICTZm6SnTYU5+RSrDXl189RMU4JLfuQJ+eQ+2m/bD1UVHhzDjBJITpsPymF2Vrw5r
fQfHeQR2OAZ3n6hbmdezs7rQUItu3BzxczG/LBr+ch0K2/VE+xV18AQ8s3NOJYS7mfbdWSgDMjRZ
oZk+1Gxich8I6R8JywDkOclPC8/5IFn5dl2wdzRSt5htypjU0i0RVQR65SUSIQeM18nb2RDGkKEo
qDue+qPT7RbVdzbjjygu2Y4O6mo9u0bUP0s6czHNpLF8WAGgG2rM4dxIPGkRWfu2lcHuiAQ6qm4r
+rkM/37Jl+N9U9PQ4QrCuP5QJUA+s9D2oN6xXOfS5NteXIv2chUE5fbvCHmnVkMJMVhj6ELrtVsk
EZUcj7C1QTbdIvbwOfDdDIEi7JfnKN/kWKO7etfC9iV8+1Phq9uDu7uCcnIgzep2BosaeyglB30z
7gRz+6E1Xakdw1xiveFk9xfLJggMM20VQoDSA/MxoIYWs1KoUozWsDwJXLP4DtzJHaweEE5ZpaaE
uzIkdoJU+QcXtQSsV2NniWILcGrprv4+QKRDipR6oIjdPffyWPckhySP/oSEse58quOG8T35X6hC
n299zEPAVqm7135y6ExytiIREj+ywvG6WFRDqzm1NgeExklru3pP5V/gm80NcdSdzvedaG87+/Bq
jvV16Hqh7q+YkiljD0pDzwm40ZdN5k9gnUV3OiOwAV6cPQPD/Q43eHDBWtSp6swlFkAtiB9Y99RB
lCEhjj34A2IK2eyUynxUWxLhijs2IQR2hmcc/Hux1KNBk5EOjIod2L8KK0jDH5lU1Bx3IckQ7Bjs
3BaQ5xkANVxVM3YQ+gH8EE8NJIcgbjHtEnwTH+s52TB5Xl9087WUWkYh96Tfnm2m4N0IB1MjEz7x
slS5Hpg0gSymgqgqY+j68Ohdh2cf9iSbusUpXuxrpib+wOoEUaldr4wbQ+sGOTgR+DmCXFA04jrg
XYgXbonpynFQsx6vh+EWataPBuSD4+hgENqLdSkcP4zWusHD1MU7ID+cEcALQmNcoGMw9oXgCcL5
foP5kRrI3wD/Di0bqbCcjXg1ops7uq2/evPH9R6N+QIlSfkkS6g9vlZl3nMsYiy6PA0mMrvzTPsD
5/bL2MrlkNwnd+PwGf+shEeeeIJr2eEz+K/7ng0S5DzSx3XqFdn+JYkCx2yRfwdHLebkLOBNJYf+
Ca2ifVM1a8hilItIBnzhfU5ztN5CRqck+1BD1kCooz4mrYKUcE/hvrkjHzy5HAWP5lqT2I8vCF6u
dcvf18lbS8xObG9yv+pZtLJuWYSqteDNEqK3uDDE7gmOudV5fTE2ccHhDVGLEclahRUnys/RpO0i
FpmLt8C3VRY7YQBV6r32uYTe17c4JcnGYgyGT8ncuykCGbQlaeRCqiMKpncEppQ4qR3Gjq2Bsysy
ezQvpA6g+eqX9f0UefqBFRsqk5EIHDe1Vdb3gAPbuMDlq7auHnYHucYvIV4zgoWP3njkHYeSBuqw
iitgsP700bTFtTm1Q6gfBy3/PFVWe5Jxgi/DvpsYIDkU0Dk05fYm/ay39kwN8WLG2Ul+plqJj0MR
YcA9k0patngyrLdG/Tqg+3Xbgo2lAFF+KJu8jZRYEtHRww3LgK8n709/1xkBgvsBeEkLxylBg/UL
pnL0JlFH65V9y5Sk33vMLxxgsXchpeuRBEaX8gY9n7eSDI414q4kwOp6FrlP8cpSoIRZqCCTeguC
JAAFcnlLz4ccEpcJink/AwmZTSzuK+k+Z0ujqoCRqMzh+iDk9DzdGudBjyeh2AgAW13Y0yGDW4n2
E6jDPdKgR6081MerBTC2dneg6Qa2schcezmNhb5rLQB+HcvzApuaIUUBfza4oDKV3Y8mfiin3x5z
JNJlhNj4ff4R0pkAhlNW3gErHSMBszJzDHlpfqb8W9h5CIy4cQUZULydBejnjJPQKxJE9bg3D3vD
K/pA1HUwJCI5dEb/ubc54PlKnbCF+0uN+qKHzOUM62DPQwqBk/V903uTgOvfCA5Rrhxf1wuOXRvs
ORSqhjTsGAeZ9b3YSXN6gniJQmpMsF4JIiQA8CoaeHD34DvhDAjBanGKArQTLzG0pfwnk7HssgQD
mzxVEaR3v+I/RMsp1f7oQNtUPAS87SEY0pFhgqFn4m6HSGPoxfIyzQRPy6OeZnWwqR0lxVJ1PXIY
Mx1IpJd/2KC2Uji4tx/zu0FPi3vGyHCzozNtFxmo8QPmEQEaRILQvs1D9TySwL7CxTHat3TFEuOw
m3fAUhw6UBwiSfCpLDvplH8pDYXYdTbitqdU2Fq5Pt8pEofpqsCjknHsMcuNz4dbuGjcvOXlaAQ8
Gr5TVZUBLs8um0MDg7bAlxZO7/aFLAFLB/DO5xauyWbKL7zkRVi3lnGDfuiklC30Or8S02UV/XE5
e9ik1EPcMHejhYsIvfNXFMBS+Gje66eboTAZ6nYfcD7OMR723DGpNwiRuZpDs7qlbAdDs9pFnHYc
reSHZ0Rv2pJujV7OSpysUtaeiEmeo0Pa9cMiNqvV29nhxB2wLBh/po2l2IXkNy0p/po/X1W8jweX
ux2ygPh7fd0PMZJaxo7ziOowURDODV0/tAXX9WGvpTrKZSk04P/K5bAsa1MG0/M97W5h8F8J+GOo
8buPz8oCrhiofCBEs9g5Bc2i3Ocm2OXhhNhbKlY2AvF9ajOfIoFEKQjz05a5gt+DYDXS7GwhKXuy
+iJlX+Bmj2c7IDoultkyDCahIUV9FOJpRuGFOn4lEoggDZZW8AAATpBAt67dR76jR7QrV+1NL6NS
Lf4+fL/20uLXOPUwgacr5fxObeRrgzD+o2ln4cFzr9GM+3U9G3Rh0I8sTOM+ec/gXIGLOYPXFbJT
re7wDLM4wIg9uBmrUPaHjFcdbMLd1H2RypVOYic4F5mowLzJrHLghV98OqzzmGT5Slw5u7jxKqT8
dz5c0C2b2CAdgrTZBT/5/oK8sZ+0Q4U6VsiYLQ2ti2i/x9PYLZNJLe1mZf+SMoEQU7i2HJR20C9u
pmCkWqWRcN8lTBT05bCY6KHpaAXkhINimASrjREd+nmgcVGtv7qK2wrcd69EVwHRI+qUhYpZHBHx
1LjxeeEFjwSTQb4Ds7flogtSvRdlmQw57g1qems52tCJ3tg6cgeJXIP2dq39RI5rFOQatcT00mlA
C/fFkcGLQB/cBtkn2e5fXqyxQiSvG12hnksfGamLP+fwmsc9jyxZ05Yk/0bMyIGTncKSA5rr3gIJ
vAfsPka13OZ7OmkbtKQSy4dkEMhffTESmNyZ4chilBHtYBnrJtGr0vu6SUndFLJVDR3Lb7Y/yMJU
nxXb3nOXtMqWyh8aSaG11Axyh2TWcAvNiY4GvkTgNUNjM9SJBfo8lfV9FDzqpHYft9x+yuDvxGFA
CFozC+4p8pKIMa0cnpNqBzruwkNMWjXurubgT3C03MbtHdhZSa8wvffXepwocsH0Q9gaBn1cOI8R
5GWFKqkDZbfxAFd01KtJNCoHnToIj8nK1wk6TDcUfLGnD2yh4Vwv0Ty6ZBzNUn0yeRAw6e07hqvj
xQWx+VE8Ti8Mhx0w1o4hqeAuoRQNaiPG+M1jR3OUFxAF+obxtxL7fjwxgIw9WUydyk5/HMsfvn6W
IOeTmtAefG614XrLuYKnfyxwHIREn+yhLuD8LzlLcFNRQr5ghWNOQmVzrJwxo0o/9BRSBK8EOTz/
HQpId0+i49SFcrK32T5hS6AK5+pAX51T42xtSkgy2Dnmr7VdgvzNXp5memjS2PgtEeAm69X/3oX7
9IEAKkpC1kj35XUdu8/T+wfqE9kkapo1y3od4XMCeU7u32HqHFStUuZA50wGIg05ByVOnlLGXgIA
TgUUUyMIQh1RmVI0fMXE7/exntbGwzHqDzIy8tbc6i0crNYOGVMrZtWEwevuKF0UyJiAc3gr+jBy
jXgYTnf//s95N93w7gFUEA6C1pmdFb90Con7EwAWrlC/RYdMAQPHvKA1aUKfksIenypOpr3OWDQ5
dSuIzEMm7xvYFFowthG6fw+rHKF7lmj3xnHAa/wFYsHF3K/aUTOgS+0x3ib5BIg5FP9cIASRq1k6
m3Kezw1lvpZLvi+bKzztOtcjTE8KSzHckqK61oQLml+D0/SJ5w8eZKNcsGZlKuRcOovZr9UGP8eu
C5SNfzBgz1TlfpymnNgaLWnGn3t4elgA9hORQjZRmEwBm+XiG/dplcxZbdkIxMjURhMwP8GRP1SW
quadKa3Z4oYd2Y+Ct/rCPq8TvascxP0DQG3M8mDy0pidi0koAxn/e7biRLMNZbBJWw/m4Lxv4Yyl
dGxkE8Aq6tI8O+MTJ1AMPMMIxD/S8di94kBHqvFjDKZcfSfyN3/ZRrnlixNWxOw5c87NQC/WnjfM
PHdfYpmhjuDW3LE1324qUhOGDOhMcynRZD2y5lYQt9QT7SUz7CMOlqZ/O6Y/t5oAw1l2OX4PjMjt
3wZH4yLxj7757ClfB7B2hlppP7yOafc62TM+V6RgiEXnBesF5uP5s165ODrfi+IAdigQqAQRNb5t
tya2GnX7qR4PW0rFCgPijIj6xkh19rPf60NUkg3q27yXkotWRn+4quSfLUPgK56an6RZbP/7LbGh
N3KyGCoQppuaLKl+/ihoaX2ZgpSmbdUUdz7yDaGqS7+y4KyD/qU5SUFy1WaR10uwtSeV3DLtgpvO
kuQiOiUlNhzTM90t1/UegCPlgi3dvDYh7zQ+hGZt6SWBT0/qARXaTBQjnsFdYG1+p7uCLFZSMYsE
fYJAS4DCVvSeWk28FJuLhyNsqvzHUHm6rsV9Bayw5TAN+sWXtoG3nyaCjojuF+2I72z7MxqXWHU0
DcqdBoxKE0jwvnp2T5umti+TN9KwmUqar2nV3gfXGentMuQoysw8dbobJXOwY5IDhdfTMKV7e9mn
kqFqQdamrOOElI131QTnnOV/vE9S2U4yG4lvnzfzdYytgVkCzWYc/5al00MXzV3xuwPChChKdlbu
zty3Dv07hsWClIjUNYfDlaszMw1SNQT6tfbBsnfxASrzVPaMI9Z/P4vJ/Wk1d1spusKnansXxLI1
wyyX8W+fJ4v2BRXXrIjPvAqZnx4fWY6sMjwvbGs5DDcHae/9R3HlCi8pzLqT1JkrH1m00c6OMHZR
3UefZOmd4+t9pQQ2HU4Je8bhjrVRmYhVJqQ1qfpgSVo3y9ZOAO3pmPfBlSSwEBRD7UAOhrWr+dZp
IZsdclQFeWT+UtQc/zlnZXoevqBCC+M6Oa3Yrmqp21TYeUQ/Qxap/9TLdHt7S5adnCNufiRpMff2
Qus5y3NJ6mKpr3Ug27OrMCcGz034jB7sNujl1kbK9L0YmDfEjmwAazLXB7g1gbHk8qnJ2Tj8CB3n
+RcbLPHmYKEha98aQkr+yr1Ffz4DFeDENAc1hvd2eGlwTja8texrQaG7d9llBii3OoJFACJ5Ghfk
Yf+l3cChQkIDUUTH+PxAuUyJAlrHxdOE9BE3m4EBVM38P7PqtzkTZgaNm24SMC/v0XbbWUn3/t7L
C5XKvB9OpSIRCcIsugvexyzLQhM2kzbyqeraL0haTk8BGc+zPmxe1ONoTSsDz/T9t+5dHtH3gvdA
H1rsSAyijHadSqigEXPln/UGiufvhdeUIjrxweF1vDSe+ZkvCxnDvmiqZics3UxNdLrazMFhOHDd
/xRorG4nt80xreYjD2jAKOd/cmoFZ2BADHDCanbDFFwUwDWqgT4dAPzuplLonMp9DuSApbDHd1Cf
EXpUlNPT+tJASrFEibRGOZDUtFNTV2oYN5Eu03A08YFhA+p1/6PY6CnY2zzsE9BaqCoWpR4B4CYR
9LmJ7A4otP6y6xaf+0yy59ARPR2CVo+Mjt15DhMOS944yJUnq+1V8XqIt+PmHNEtb7f0aPc1V83A
t2c3zdqA1wZ4P5r13Hhts+wDv9IoXx4EMlIUYcbE1IzuIjYIJjBQBkasDKn6bFDDBWpu+J1yD3JC
vE+EeKOJ6H/qcNfHlqxzU8oPspVYUVdPqTP7CkIktWl6Io5ZFfdAeJj2STNZ48Ohq3YLCKLyoGJ3
g55b3Y1ghh6LcPvOavY8Ojeb77msbOhZc0hSArE2qT9IK6fEsYez5UlLd1FMvPfQxe1A60ipFT32
1A5HQBkjLOzYxPZFGyMz5658WmOQInRbxgpCKyi7cj+q8d6DbavsYCJuBBuXbWg7XKFBBkFGfsci
D0ac17uvzwJE5gS3AIaDs/BUyS/AIdCuOJcrsgBvtxwoNs0Mwp4Q5tfaqPK989rEuvmGq6v1bYmP
e5mHPieR55E7KCUPeixsDGxzkStXua09SXDBr1zxHKE8TWTzLDcRjFNPPqyQKlUChfwvc4T6HEmn
PtMGoE+ztkUgjMD/4xOhO70EPUKTY/ii4HzKxHSkD8dzMIAp1iE0SpicsSg398/MJDoCePIR4vlz
vGDCga7B501jfXpxIOuyWvknIVzYhefDM2bnS/+EOnWDAxfLPujCRNOMhlWLLpJnsgUM45hexEwR
fe6C0wdaJaQThs+92ec07Plto/goPsHtHJcW8gx9pra0z7OuP4lz2s1+DxRTc6b2N7MfoM6GWJTD
IHLMPxO34MgYBsULwF52ZPF1p8KuNXdK9D16dgQrsJ09O6/4gf3t0uyqQNxPH9EYhd4K9gRq3qDb
KmdNvX6RQODqv1qcIh+Y6oRoEHIxmchDmCJNLhr+R5ZxBFbOtKQfYbW+STJ6Sn/RcEW9Ix2LShDR
HlyQAdebOhZe6WJqGsZqgc/RqovKPVL190no7cwS0uKWmzBIeiVZm/r4YAu56VuOvUIsqVw/eXeQ
BixH2Q8hb6hcSNhmJ7hirw1IloAEXEhUGnMIcGkGC1kbBr6TsuqOCM21RhIR7z6XdWwlrhQDW9qM
Z2S5axZgG1xABUuexmZ+20pIMEv1OCRuGCMlqgD7HBb3NmgzgD6Y+rf9xPfvui1NuEHSrxg0VGTo
BkJPvIDBPg8OxrqXQagBY3tVzF1O1VLNDKxt8yUEkJfj4hE4IYVYyd2vKhc8Be0ao5Ueio73qlSl
rJiwXWZEHeR0CpiG6wX5Xr574ff7Smye7LWhZQpvSLMWn5oAv70KK4tYd8MrO8AFtvbAVWqTklHt
bTw8xLLuB0IW3pPO0Wmlp/D+RtPAAEIqtBxW74s46/jb5ZS4X1+BydeSbRDsq81S/ZYDIOJLs7UJ
cUqIZz8icI1Jr9mFQSqEYWXSI1QBtWHhwKYJl+a/vsQjAf4GCqTVy36V93/Y4/ASLC4WdcV6kp5T
gUHO6bbmo56+zOBFt/nJ1idRgoXFM+SsOFB1Rkl9q28uEzVeI9SUZ2VwZsI9M+Q+9HCG3dT4CW5i
PtQYUBUH+OfDUG7w2Vx2ed5AArpzW70oUu50p5kMYLqhYEcOto1SWUuQ/dEizawkxghZLamjMZov
f+CVwCzPAGlsYvf0MyEN54NuLRbdx7bBaRtWZiQFWQe5GZ7b03bsRegEW2++H2Dk07qvLND4M46K
cve/BCREDhDLrn3ldDkAs+BY6K0PAGL7MLcgsBbiEimkaF+pvXaECTTBCjO/P6xb7Wex4F1IAYU1
0XYtTJOfm36XQ3uqVOdafvEaVICOLvi3h6PJPEknC/6DLGDFgn8isFuM827+q7yBSFNIuqg93kKb
4iPl2vtQjmFpJKvjxYRSp0vrijY6vWZjgp0YccbPL0Ox27Z0eXv/C0zyOW1lmpI5/QJDOUwCykcK
j5uuNpqdT5dAoVYOpLS/rvvToUvs3kDYOzRQDqvQH5XhA1xMdIhCRlHW9XOiKYuQ7c/FGBL+zyFx
ax4TW9tmok3z/L4j83557LzbgRFId2B0sGlqg9sLLKr5PTZSrmaerJPC20EJ0YGkAX4cOsCWpphg
yhWZkIDLoRzQbvLiTHuGENjAbMuStm8JF9zBBvVKqGzlW+6KQcl1IAiJV7lG6LQufwhjpAubJ8WF
Zos+tA9Q1ZavroGT5QLgvQHsIZA8uy35uWuCeIAIUablV6WuzR+H4cSMKVn/AM+WqzPEaZp7XHlH
Rd4oOAt8pDNpfN5LlP4dz7+QuAslLhe/WtLPpBeongi1RDIgKxkrMJ3KrbUvUWRLWCsB5vYuHn43
EuwebkkVNPC3R7seW/BchmEwBs+gl9C6joyu3mTNL5t5elqnnKomlFIBJuKWAQNP55azgqzvqu3t
PgAawanlRh/uzWFLC6QpobYBpp1bndMG/oRC1kmbsf90KunrXtYIsjPU/4k5AFQXI0iK+wGwL40p
cHvPMi4frwcoK0a/Cso65hu0KknGihwUcH2gurlfgJ0TWMQVpkP4aT2WGU3GNYB3kX1hVIW5oOG8
iRof0LNsq8EfUYLArDcokFdoqHmmbm7aKnVczU1hIdEWADOtLNITFO2kjeq1FME2GKxQW/0NbzCP
LuiN7zDOinvZ4pFmFwtFWNGpksBeiit7G9hLqWMVsnPfY3XHaANRxDWg3de7guOF00XO488hREg2
1vcr7XtJHes+ZL72eerGSl0Ee1VWA3g0tVBGR5rf0VlUxOuypeUzvzF4lZ70jRgIOasds4eH5x7a
tpEIZHKpNe67AYApNcJeTEfliMS8VdAT6ywclAY9dU2nzCD2Qwm1THq7fUsUap0RK+stdj789VpF
B8izFlIUi4y3t0vIpFNae2LDlPZH+h7bl2Opnyp8b7Rg6L1y2lKlQq8bbpX7ByIa4+3v7PBfF4Sf
dd1wjZ0ex9qzTY7vD2YnMh9cm9Am7C+UyZQx1sEE+cLBaZbcLXiGi7oVg9yH2uiOUV1YsQR0D+gB
LGkVRdGlgBhgaYPUnvqgKAs7M3B7B624NMCIdeuTBWI34yLy0b32eAZ4KJv8AvYbdM4NeeS8hYR/
BWc1uGtLxsKeFhry8sJPQSsYPglzBihHEu/jJ3rvMsMWXzZQSVU4U0xI64gv+EJqSQdKXoZFP5gE
sMyN/krBeekDL7PsNUqAqJ4anmszO6dib9Gh/tkr30G5Yhx/ndqOp6JFGTvRL/CwZQ+VUVAf0LEx
cRjjx57O7Shq8qtYhiXzB5Iyh12D2oocUAucw9MTRZNsyK837WNrpcXlnpdoK75jIMQagVODicNi
TvvpbaCQ5U0gxSmEjgEoI0F93AYYn49IXxPG00XT27bwRghShcycFv9X5Z2KbVcz8u97XTgxPDpv
K6UykNWlXsloBYY7t8kJG6oD1iljqECvtJXd7qf7K97Zoh2BHTWPoINPXeH53j/nYDRj4muKT2jn
2XM5KuX9AByepLiTrMD0HRo1bRaP1zWQJfcQWfOKaHG89iswZCO3hTk1C6ByslJnOU1Y4Ma5IDue
XJw4TRu17GEx8PUK0jVS+S0UYBhhwUdAyc6TdcLpVt9S1sbXYzsi+HGQhFXK1aEQl+HOIRM5cTHd
nifmBgTP+Y1GS2fSFXmgHW3wmPlavWQXQ95LaVjMHreD2nO/+e7bMTBZXw/0/TIULwUe2PO4IkRy
10X9EuTjH2/MBel0Vhv6ozNZKby4zir1Zik30LHxfivkRONAd7/rxtL8IvdtvJA1yK01ArPvzoG+
XvMzXgHdV6j6wMf/XtRSXyqr8fqgsNo6yMKV4qxzFkkjAq/AH+CSZtJhKSOfewZjY3Tj0bbgF2/l
GrTxIqhqwBliHnGPdztXRWp8PNa1xLAXW4xBKC8gnbYJY6R+zvYD4+yND+iKdumDXSEIfnuUjuX3
RdSKmIBWSEf3c6K0zm4tcZxuaDUaqhFGylVFXwbdpJJwq/QfUuQ1pXu4gGt2vc7nbG1m1Oq1dJHn
C3iAoNh6ilb/sTWf2sHHhPtVdZPsZQfv7nKDG9dpxXjLz9MS8G/NX1ZpA6GUY2OIcSoWAdLnJdM5
f2YW7X/mNIiEO67kry9fA5+lOD82UgXTptPPcHcUVerNT6CL0LfXh3ij1916TxV9qLtXQcsqr9fw
Ax/8cQWNMpLJS6CMn4A2FGq+AKDWvp1/VxqJ7xK8VCtqgay0d6mtkMfurpvthxLlW7FeZlv0U/uD
u88CMazuahTn+MP7YrtCaWkzHnef5bcVzM1BOfJnIwFhUeQQBk4cg92vdsIQpCOCk67hWMjSiFkT
VF2T49LYw3uU1/qei6q6Hy9A1N2kgIRdecgw/EstsqRvS73Sr3zZY+h3jDuw0BLlfedqAqnm8pmj
Vk/IZfhoY1vdTXKjaVQ09tVCqqhXibkUYsoNeD1LKHodop+1O0U6GGv4BR2nqVdnNh/+0PxM39+W
1Bl8D/NK1gRrpZBIZnvVrVQn7eEBaJrP5AUELOS6iScoeqKBLDHKLEzcBaqHhSKURhg9GPHVtHv4
n/Dr8Inp0LJz7huVMR9/7PuFlBLoZH5HimNUndchAP71x8Dqi/Nv4lFC1QPvNCuf8BGFp6n96xlj
28FohxRCpcTNPQZ9+RCKb0M2/1P6Vstt2Bt6Bzg+wqofb7vSwaw98E11fEIkyrPhtA3EE0jw50et
m4lH/jqXgb07lvbDOIqm3Jo6yCGl98AsqF16fMMKePqTxOyD0pA9jMZ1XTBqvC+BGvghq/0yIg9p
/5+42f7jKdVhAPRzZ/AsguR/gH8aAm0n56wq2QU2gYCtNRsIKNgxoFIz9BLtDjLKg7KC9BlmFpF1
W/ovwv6wAPXV+pOcFlREX3mbvHwqqU+vaDO1A7ixRIqu5TyyIs0YIcRfhvOqxZwTzzr9Kmi6Lz5n
5YdL/8L3qYjKxPxMUviwFOOqpA9wUim5ZpjvkPs64NRYbIEgCFWE4+m4s2RId8TgYm6+X3ILWBI7
lia17uNeivjIgeWymrBqrRWdoIiNEhGUH/TnnACY0uaEJH+ghGCGc8EmXONg6i68QMxLW5WhliZA
N6BhvpvRfGyWnVGeMpx5abZ4/zPiuv5hTkxJToqGKw40mqmsh5FiOxgbj1H/VrCDWdTqD95ac+cg
GqhGRwujiVvYt/5a/1qAia9+LzHYlj+nhDV946+Ahu0gVIMiY1wcSWXK+zqly3QJ/cK6Xy3gQXXV
UFLHZwsfsX5VHBfYxr42LhAtlSRLK0XSxU4AK40w3iQZEZO/S8hf2jI296h1E/KjapQi+nEH+Nio
nbimx0Lgr7lt0sYv0/74uxn4h0grM0W0O1V9qLzlQ+INDHDifAhenyKOJ2eKdNO/cnVTSLNkUXWU
/LJQt+aFe4o+i2rIW79xGCEJI4NKd5My4YQ1h4m3Wm92osGnFe4P9uHGd34ot7N/9Ropw4q8mGUf
8Y5XrGqUkLxBOmug7kBXKNsz4QwQKKsZ67y5wvWNVOzMcgnKNeKiXwCpf6h0EgE+t6Iq7Q3WYx8O
Me5U9aNJWY4wE7BjrL2+1Ib6L8nUjokwpC3LPnGajxFomwsbvjmw1vQH+EvLRpXzrtFdn4JxYazY
lVRfCxvrZ6kB1oWb1yy5yBFbMTRi//AkWws1fDncfhlHkTwsGNYOXXxvx6BCxKr+75kkFVTt50aH
iimgXJ9SCvmYrW2P86FmKRGS/bqUN4JiJfsrJcbdFX4mAanO7uMMbLtkQc0wzb4XsJ5i7QNxcnms
SYFdg/zcIl7oEaaqGokEaMA2xap4mdkgK1GbH/CkSxmo7iQSssYfC1YYGG57nfNJX0O5AG0DT8a9
2SAjMSG9oEvW8pWK5Ka2CTe2dOBnUuShpY33Nlz6jKMOcK/tyRdmshp5fKVCCN/yuWUS9mm27OSN
jLCICaMluFnUgluoSd73XAtEnoJw8HuwrsnbYszb9tdfjIyW7xfLf2ZxmW3QjFg9VKJArg3ReYm5
x8HCpHum/h6NuNdXijrT/jl4hTYrFN7WEtl3JuoU8RO6xzbXtms3fSrxjhi0uRyZ4pIr4H7GBUyQ
LKr0JUz3HfcjfpHsiVwiklmyTdZJiDjOvUT+2iv1A7ek7XOgkvsH4WmS9YbUeddzIJJIS2zImjXp
/+fIiy7LsnXwcaKC36GxNJ2c87YtHXJ5ZLFn8O4+f1pPC1n/4gtNZLsMtHomJFB9cdO8UmA/QFcI
TZBJ2Jql2Zy1Vq2jpcG6P7FOZw+RMfkd2Kzp+ZrNtnIPMhSLtRSnMF0dfycjoXk3EFb2zLFEQyaF
A+7XbOH2GBzlLKI2sSjt81pbBGFF/PF6xt9q+Tg9Z2W+aDDlTDlRtN3N10UYEtLFfD5zDGuZX6Es
Y3NOek/DpNlU1x/E8cwQGwZiEupqfB0uUR98x8gn569vAuJAJq1kA4e5EQJakff1UusBBbrqOIL2
xN2dLqZ/bO5FWeKgcxPLQT19wK20RixYYaPFUAunfZlZ4volm2W399eHolwFy5mSKJ6josTeREU+
2z0wEF+rw5BYBxlbZjzcsXm2DFHiIWBFhqcLMzpYRaEsk5Pr7vJCBXcKPZPbPmDk3PitLnUk2dqr
uhAUFrXdBNrN2aaEsmQNLrKpGlZSn6mqOLjNo9q202syBzGEUrirScLVTQXz8DbhgPuxOahWxSSa
k5H9gPOSNUg12M5dzqLYQQ7dbiuvaQrjSNfWDJ5W9mhuvCayZ4jrD9rlO1/3SI4sL2TeMlme6XC/
iWl6sECTxD+v8Jy0C9EE9HTh2zJEXaEFXcusy9MPDy7SMFDcsLdTs0qedw2pPCcvXlo9Kho4XLQB
8mJNqzKutz9/sc0XYYq1aVXUFBWN5BxkkbelyvsjCfucrYAgoSi0ze1mSWD90je2ZvxYwfKvCAJp
ib4i2oKbHkBzd0iF++kczbfN7IWCOMqbZuJBAAwazCxxVHAMfvX/uz9fU34KUHG1lToXIHU1HLzZ
I96Y6xeF7iM3/TkSHURBtNbP40Os/Fa5+N+7TiMIZKNOxbv8grgCvrjH4Hwe8dYvgrd0HXHRKi4I
Lz8AXH3XW4UIDP8/rztTO/5hGN1Zqec+OKoR3PijCcHSF2yXVOkwx7kIi5035bORRWRrbG7+W9ME
YotLn7ORjbTG1DR0MpYzAbHMA8UoPgGyxuI8TQC0V5VRuSKuMNAYpOWJuVc0JVJdGCZdYvyQx52v
o8WmgBzgpkvhupjy6ZNE0NSUTL7pWSZy44HeOGCD0p0ehAp1diqJHCsu3XBNfSo2QH18MFr/6zSj
6eWCknOZRzgi650G6jX8dZuFsGO0l8zXVyAADYIUwrCgiTQ/jz1e2WwYURt45vvt3uWkikCBarvG
7lCU9fC+jeVLwxoCPWnlO1vJPISYZ9gxxoNs9NEngbLop9RxGzp/7duWO1W2VukoLrrfZgM2vxp4
KijvxgadMYE09cUIMDjHR0I2oZXUBvQvYUwsXPG5fQx/Dd/8mBbpo9Rg0z85adL33MKihKSfDIaV
0pkLhWac2h1r7YS/CWlr8GutY80ybX+X2tMpoeCoPfbUOwYiHeUB23sY8RU9K9dywAIBfwaWwl4o
Vwl4A97IVP5t9EtT4z6G/PNJfrJTZOZazIH77YKkYX68pjnb+U6L8nLH/+c+g2a+B2JROgidHvKC
YT6H5jCpztW+jdYL1naD+ESxFB6jy+v6QSRzMLk5yX4/kfbMep3bIE/RFzoaGS2Ch7PK/mKwGrHu
Lwdg+xqCLtMvtjx87dfcryY85+wDJbH3agRVjU7DRiBAYFxyEmApO72I09wsC88E3qPc3n0D7oBQ
Uyn3EyFVBdS37JIq865vz4tVOtXte91zQHuVbAlBdl5Sg1gK+WhgudeP0b/K9iNP1xZEI9h+/JeI
kwvSzUOOa2JJ/TdsU9D3xuqf1lHxM8RN10nygyOtb5Ita+PsIz4h5BJChSoNqHffWsRxXeXEBhGu
5ExhqHRCWmktbNKKEqcxcAMBqiya386f5UN/vhnDsR49NQ6u3gnroAHJc+WEoCQrxeTRYvuGURTy
H891+qpTJxBWobwDjTKPOsGNmQUIJlDuSQmoQHYSTnveS6z2cGD/+8FXxZZehsXq3ECtp0+1stnP
94A1UvE9W0QpxjY46ZfPKLg1JhVFSTa+zsxwN9Mt2zsdmXTCxmd5u7vbXdHtr8QiXXF9VlMcLf0Y
Mpm3AszZz8jvEsx2NTaDkF4mUqpmhW5tfl5LEOrW7lSgf770M/fx8cFUnB02kG9LXrudOoyItTjz
7TPVHxB1imzKe5wja9qGN92X8D0UEfo/fAOXGHHrKN9wNyi15/JMfBldUOfwa/Dsw2A+8quBsueL
WBfOWEmULzooGgoxpQp6/i4Z2KbIuVx/DOG7fCrJo+RGAXraenHzxxHFiWv8u13pj0FAWINOqT0+
ePu8JPok0vm+3ah1jEaeUxDgnohM+8+yW418Yrt0++biH1fDVyLW6oi/o3aQzQ7Vff2OpTJ1mCvA
AMVFgLzYxwWeyAhEwWclxZ6CCQqLFUi7vLoBsB/+2vykofivBA2a4ex6+Br+JIMffX971+UVyV9L
Ck2KPfkOQ5uK1w309LldkTs+bSdFFRex5KT3YUXn8bDKxuYHmtUt4oa3WSo1xp/1YccvNMfu1ur1
Bu4HaOW25PKh/BOix9tU5oUY1Q4Coszv46LF9fuZwSW45CL8Cf5rBEJWoAKLd7n/IFdqoGWHeqdf
vOIFlWtjE+IgkfwEdhVhs9qCPfEov9J8T5hdeEMTAjs5XrcGmczh76fT2+RxxqsUHdGCl9BP/Dba
D54YTY/b+Ib/uzewLmekZpKSMIYWlJsA8BBY4RJo2yjQDKST+NMu7BGc8twMd1dwpXTUu2fXbvf8
XLtZio58NcmOrVypDPELJS35lgRQ5RegmnYDYdUX2GIRv5CE1DWnSrRXfFSuHIKElcpMrStjEjtX
ewA/UN4JFN7KP1Z40GokqDOxNcbLCHRXCP6ZnW+JH2ZWLTtsuyU7roE/D3YPfgG0ZMT1dF1pIJnr
WmMvkdWgUxSVHKY0gU5yPZaoKI9Gssvz0Ds8mnuiaQfjQTwBC6GCNEcaWJVEHaRmTEWnKMpPQNcl
oywldIQW3N+l7jYSybVcrFGXVQdYJ5m6xsLM+4aYwsz9MEj3wauWTzAcJ8ODb82eioupL7Nb97Rz
ls+2NGZA4iCJAIMDUWEjl2FR5emgLPI9Du9SAk4d8p+Frm472YxlCfFLjszlsjQZGhdeW6YZgcDc
S/8e4242i9W0MdhrZj5cwMELUUD+bj4DOOlo8/1R6eaMJAt4VTcECbrr0t4DCBph/yMbHHPFVLC+
LBlrgMzXJUxPvBt49PLFmywbYw3VMnHqBf3s/2o+ZxSMBdSZAlMFsFvXv8999XUdntEHUGag8Tnj
rlcHCSzsFYv34/AY/GyuT/xaaspLG4l1OQgEF67/0903fajPYswIm9Ojxt3ZBHS/Ec2hmmfBqU5p
ZXWt5BlTNSfmwfi7WN/xrUm/lLiFiAoGqqjXjN1eVZbgU/UspgtEPJZkjfcCgUxeBpheVNMDJ/0V
roWi1d4Ouw2xy40bsU+bRjuFhBFpbHdAOKWhto6000bb1q+c5oIy4gfqRtz4PXRanXwPHpBm8Qc1
u4AloWiVHHqSc6/E1buaOd7Q2VRyzkeqGPJIl0ifaE6ClSPp9/i4/O6I39GChmHi1pzhgJu5BXHJ
zie/cnZIBkApSaWcvUMnMEXefTGUH13KxiRaYosHBQVuZiOLQKf8BZxxmI/4AeyPGho3zXDXMcX0
aYR8b3gZGV+Q+iEgJHPmexKCwmKm26Dq12Va/CWOwQhOJM1kJjwHSdYbj9tRYuO7j2IZULD4SWBw
DhJmNOnrwgxmEoYaxEZCJRSDrJHCWsueHqxK0gy/bVrxCSELlzAmck7Ay85OwOtSv7prPhDedk5a
E4MQV00xFZ3yarNtvXWTjkY5Zq50OIbd0WkN3PEJ1UHE++BZZeGFJ/4K7iX1v/tcsQgxR5+qs19B
EPkTDBYrcSCGpU4LX7dK5iJuN/EAjWcMAQ70w5hZn0J+f9j6bnuC5DS5TJr8IFtIJJfp4ZEh4j2p
9bSVnwpEqWRU9lmeNVnCeoDWXg7rdmVrm/m2p5XE84K7D4oSEOX1ilO/mvBlNH66Xm+BDY7m+o7b
fRZaeuCJIHzXmSTJ6yQy6cMHCvV2PJu/QCcI7MpZepFAt1xTJqbyr4eTsDq7GK5rcTOBz/CZTVaH
wXMV+m00TeFEaDrjg7Kh/B+fZOztVE6hL8sjAo9zLSojAiE+aMeK9t+SgghnPvveiOZaAoTcm9z5
8B6/h9sIbUiDSrp8FsnauuI0mm0HZFKjsWKnE/TXxv6pXisfa2bV6lJWcsuk9hTL1UoKsERCCsl/
eiaaYe43K0hlEel0Cp1JfRx0gWTR0Tq/4dFr3HjHjrQLUKELV3W4Qhh2IaIcLQMaclYEAB2LwDe7
mkz+q3DcNASbwphyqgsnnBmvGtQA/1k0ofYMhcbpPSPQPOxh+wcunXv50lFDPanngOYZFjSWd2Hj
g/x3lK+ekjEMlDjqG083K3HasTspEn2hvJYJliCb/TUVgBFaSS1w9ruSrn7VApHrNvBnobqVi2DI
OF6UbT6Cb+kq1tbE/VPICpLSdcvuSMpoU4MNif1nEaF1k1oLZYlhmpTBCrM7p6Ru45UtpRtKGN15
UadWoPZs7LXSP9SBSN5tQeaZ6BQohGUslHJFhELqqNuaHL7uSYKsga+GDJjx66uBqt+xhBr/nQB5
RoilDeBWBX9HxXUh5uYXAdl9ou/pFMpTwnGbC1RM8nG/pUydz+KHJ8uI/Sx8ipqeYq6dxhv5MAjw
TGQs2ARW5UAY+KIZxLTF1r1hd6rxOSeXzaQQV0PE+GwAjmjsIRzEVYNUXfJuXxJ2cPSax9AolBEW
0/EgZK6oq24fZ5P4a58jsJG4e5GoXfNh0iSn6LfYmMWqL8Ou2D0GtKcQHZQPCaaWD0e40j5HkvdN
e0XXHKoCjhKlAwYAiZgb4iHHOR6mFWp9pxd0OGiwjNpqpL++MsMiS37Pi1xtcVtpA6bB4VZUWdKv
DYOTcoJJzzWqv5SgEcCRVjT1/qahD946ImnSTqIVebP311U4f5+knB1VzgI7Edn+CJ7hBC+lRXF1
NajHXCwHYYOLmfmSjbUtDCVnpAoVZl0mRFXtAA94elznsIoP+wwpnoQ6qzQBSoDKF5VOj6MWBaR8
ax+clxK29f1DOgaxttiT/pvuPFMB4X0CecpM7kG99R8pEG5W+LIrblx9Ssx/eo1uFgWcqCcFE7oA
POwDIRd3dizv0XUrSlbTRgM6Wtdd8Sr04S8km0vCp1JMkhy3jc/g95W5AiWRxIsxaJolSLtn/+iW
GtS+68I4e/QJhMnW7+0ZJEJPDjWynbN3FyuhKlW8FYrMkvmX6UKzHMPt3yrhA012xhZv2KtW3TCc
7YzdRKlKicUAhmumjmbvkaoOnFXtcsgURWaFBXddEnsiMdKHD7YsS4N2JEfyUP9NVfsQ5dAbfmdA
AwZ20DE9stgrg3CN80EY8gzwY5XucoZknzZvH7Ld1J2Obu/r6NLm74JQJAdl8YfeQo+MmKbvLK0H
66JM88QJpBLj2beRPCD0rOBlA08sgctchLpUGUo0kJLl5hHAGVjgqeC6q+ejQwa7ZJ8pYBdUJK+T
slbaUgQIbpgddDsDC7uckzak9NHK8K2hwcF9vQSUtxCLgp8JgbZqqMGv6PjDBgCnuPCbtza7o4zD
hTjFl9d/y62/0w9fcGYYzvrB4WZeoiQIN7BVr7/Xm0H/+I0Ahq3V3P0k2DwTGO6w0CjYy2c/crvq
sdYAYdMKQ8x2FZXfQDa4mgOYg/8N6pilPxS1UZvCfpE4Qybkp7G3sR0uMqScDOzVf4EVTMZbFHL1
bEsPVwRhGu1u1LXiq63DZNMCKCyQcUAUKjFfUwK7lchDajw4LnqWLyr3dNKy7nG4LYIhzhith3vE
UggFPSsDgUjkeWrIHEvqtZGqQRigtX11ZbSDhNZMb4R9ZxDGdcP4RgOLLooyGxcrR9mWQXCIP0WN
wspdP6DH1d27+uANv2ar5PmRcNbTGlKXTAoRa8v6yopeu4yvcpr3d860MXkbVr83MhQKk77UVyiV
F6Sflgw1L6qlCGXvj+J49GeBFHyCVXyj/kbpL/+1TlyRH9XW9PoKfCYC/Vs6vee+dluTsawbTNtM
8uHUDLPUkyBO5D3taRlFIh75YBz9vYiSKlAF31fhRb9Ojv8UVW1s4Q0z2IzBdudaNZtjR+bq6+43
11NoB105li6vCfpU/GnAV27c32ZOQzqxYVdijz194SOMojV1e6JaAnbGlViSYWiRXLVHmJ1XEeQP
VQaSzN9IbNztC+c1bgbfwGcvoGFZz4jVyuJRejm0oyMNKf3/pRNiFiohf2KYUPQh55agJmoa6PTo
dea5zWpbKVK06oI7axeyrwU44F8OauX/oQgfG1JIO3vZy02Zm5Gq7aHTd7J3jXZ5JMkk90F/v1WV
GnIdksW6PckqcdhEWSY3HWFx7qQC3FuvO4551qXQ7tbUaibMjvWdx04RmLsN551ifNGn8TQrVnhe
gaTaXOnt28c7zEMiymtxiM3jvd7dkplvo4PYtOfp93GSpZ9/1AvPJVxFaLWopYmIrT6ZN6KXqCHs
2vLEp0BdBvKDQthEzzyO2fYgrJzsxrOW3LOhMvgNIHkLMe4EKc70Xn+8OvUtKBExo/nAgmZ04Dvc
Uc01fCd0fEfvICC9Oci0Tb8z3fdi8pY86k3WNgiagW5eLXDdxQIaFXUWDYaKkU43NG0zNuTQRZ8j
FP2BuLH5M3RaYglCJCnwfXM/g8xFVQtf3LboUNPNbLF4d6SonTtgNmun/gwQJp7aAyk9VJuFNQE4
RVtgd2uYRecoF4Ep3VuK05nrtadBL/xUc1U4bXPzEog1m14kiao1fmyV2picUJnhfWcy+nPMhz9H
aUKRKnmZWz4Ll87+V41CkhlQkK2zEvNN0R/l0OWE6wGm4ZNRULjPvLLV7AyQw29cHVwApVEp57rC
bJ1sTh/SkOAObF7eyOO6jDx78Rus37X94sN5gtiybC3MDokIX8we4TvkgwkV6muAN9hHcC2br11I
svmlFie0M1WCM6f9FeCrFeS4nS/VhfR77qb0mZK5gNlVy2vN6tj14dv1yo/td6J1/c09mtTsS43m
V6uog+M8tJWwv+PjjfJUjI4Y2ONKfeUsbBsRhm6W+hVc1ofZXIdD9ioVjteiIj6I2TMBKxObRYnK
JvX/R7p2fbvzGUWDxQSHyXH+XJWArf2/4i120k/Dk3cBR3JjUB5KuQCd+4eS969Y/ulMQy5jJ3RL
qn4hdKiy35w2FYKQM/Q7QT6dxbsF9NBwbbgPf1lGelV8Y1sreX6yCK+1Ko8as4GcE3WG5JXScIak
Iylgqo8IuTazK1N72rstlH1dxaNoKEsA73Ooaoy9c4HFjJZ3BcRY9aYu5BzwAOSznIF7syGLLeYc
YUWfRTnDf1OJYMBXFJRbFt8DdsvMUFyt4uaR42niYeefNYA99kOjQntGBLPL5s+WGfgNJCUOxApA
R52xZsvIN1ciIXhH+ZbVFJC7hVB4+jfTeAx9o0ZM28Wmlq5sK0Z3ApHqOIgKgi3AFRp8mliAEHkR
+yWLeg564vYeNASjbV2A64rd3zCLTrEmrpUFqjlvMgnSXn3TYYJF+DfXa1HOzDwdfHaSK6ACvaRx
OumvMGCBRft30Ili5VTGq8o/F2De23aGzX7cv2Z1R66ExbgF1XW1atOm8A2y5nYvAWBi90oPS88X
O0xAGmbUEDnT4XxRQ0CeFcBW2LaMd05Ggdjz500+ktoxiq51oDTMlMGnyVqtx70MHG8Lnu7+s6DB
+OuJ8kiFKfRHKyy8lgR9xTWA6DW08+/g7wdv1lyVT673E2vOT+whSsAyrIhvBvgStj/ITd8eu7ai
F/94YUhvTpeBiz7Q/OTnrCXwrkQyf388OQqtOCkVxvYUNruNDoQH1I+2/FtHwG2X8wZ/w4MqWw/f
zTFuYAki8pouyIgytBl6ZSnCPJSETfxq848tSOicuUPNV0jF/PQoylzaAov6YnerwTlwdbUoGiy0
O01xZ56MR0LiSbIoYAj8G9S2B02OYJhb1d/jV4GDRpu+8irhXLvEVsmUcjWRXGzVuUZg7Bg1EJ8E
kRbEYoxwQLy50Nj7BQVEh8m6jcNs9S+a2FuapLxSCQx57cYj1JSeI18O7eRVv7VrWCSQyU64zEx/
VmYltd+pwy+UCdXA43jnDBnM3sBGstvLTsg8uRuUUltBrx7T2S2uwDtJW7xTHO4RicriCDPP7CgW
XUNfxLQFXHCH5ZHEYAZcqZ4AraZ4J37hU2q93QriLxqMh2Fjcf1Gm0unrd5H0jPye0zBArz9CNP/
u+ObyA7Eu5kY6a9E+TbR/l9EUb+D29tTJHWmd4bwOkNGWYLMoEztUSfHHk6AvK1Douci7sDeQuZx
swQlMNmXXHlz6eJrCIqzd0RIo946IW02IbygrD67yN39CuKoqeZ3n/3WPdXiMlMD+LF/PuKLuzrX
BILO7GDVPl1NKg3BzGgVQcWByJNG1PW8mcR8YQNEOc0GO6J3sphnYVtH3DohCUQa0ZpIF5Lj5YAa
+sfwFNXAjGpIwOOCKfzbCsZpQuudCF10CimAURZCKERQe7S/b0Y04RB1mw5jafMQs+SxAQRjDw3h
VDFlacSVAQ/sE2r3a8SLFlaQu54MoY+1SdKI2gFAo84vXyEusEOuRZPBZjpQIFJ5bicHbQr2Po9r
E99tcKIgmdrjyn+0lEg+DYKjBzvTxUS4j82+SK8EUoC80ZtucKO8wqwiZydj58bPSi1rBbCGGXJv
qNmuqoZK4WC3q2abEy+rONfXW8jmwwWqWOh9wXa+Aobj/jyKZ5ZnCttCkEkhBdA3H3tRaEMnGiLN
CdR8/OQxrEB65IiK+kSGXiFEDD4BQ0jsM6ndRR7De7Ek5oudHDgJRHi+kqjLs8DZycJESIpB2uaO
BhC7OpAAu+ZsOtDAQGlMry0mlMqCYEubsWT1OdG/OnciymEYFaT23A7opyicQ9I152a/H5j4tYqY
tcc23SzLesuqrWHDJNpG5zcJvxMvi8PJdDl4VBu5/pDAeNUMc+pYy7aVur201UpMzCA/l2fdXjIu
8C/YdyJ0GbfuD9qtyDSQozhmnzDaB+tjSReAs9JZ1w1NhF8GtpSN14yc+NeSobuJ7YKOd3pYFHvu
N5PgPeuP0ULdO5zRh5zxJ1OPCSlOWP9TETxl40h0fo7kC4gcPuqhvgJirCIzPtBk9cHkfgYzvC40
/j8lL1EjmRh9rRFCL4sRbFsU2/qZW4viL4NOx5N/PvTkkKJSp+3vAhDbjB9BFAtxYmdsWYlr2gQe
fqXPE0cbR9EvQ1o/qJsP9gSl5CHEjKz98LEPWJbu60xs7PLoa22axGRk0fbYyM1Iq8GQ4tBXqqFL
G4tjvY4ZZKvG4BU7NPEZpDTu+BBaqgRMygJsAfRhto2h+SmYL6Tvrm1Osj9pGQKTnPr/ITSuHs1w
Iq1DwtUn1GY0+vKAmAt4jeRHq0UmAAKZYt47aZUXJHsNUQXGoKapQ+dwzbMUbrKUP2kPyXFwOQ81
CTawnSxlu2bLiVkPPkEX7X5qMMNSUs9QBpzbCsVgAsP5zia5olqVMPxYyl7ruFhR56wb8QMKQ8rr
Pmxt8n3vGDj8CrSQYVS5YZQUKve2FW7KIH4HUKGeOw7T5cUTXaxHaEHIqpWjGNDZUxpr/eUxXxPB
gI8XnX8zqT0axJ5ezoBDI3Ts8y3HGWd1jT4/bn2zD57ae6CZQ3l8lDfuc9Bqhvkle34nU1QsS13/
aoXYpKVRXRetgYtpLDn3qI5MBydVqWZVPBpnPnmJplNBCzBo3XKsLx9wIRiY6FTqa27oJ4I89QAx
i4eY6d60BOeUcDjSKAFxcf9Zd/1dZ8l5QyD7+Wmd63K9fPpvVPMTGSMAj1z8EKf2UI5oEQR1yEEU
t2J3vzA2liP8KWHUciZt+jNx2ObDmHllb2WFu8bVkeUCYTKbkIaTkPgFwmdoFC8a/B8kVuZEqu63
/VzZUcCZNg9D0qajqgndgcL0guH1u+3+eM3Eui9BfP1fcGCDmkWfInRMZUXz30oVnbGAziQx4tum
HiLz+OPAFDqzGIw5uxLmwBQNmvB/4PhO2ysl5M09dTnckVUto4QUFWlkqOzClS3fxVu2kh9nr8rJ
LTxfet+Bp7GtcoualmHVt8BJq39ND12VeHnVL+TnI9kHluWCVsrzWxkgslizZuUMlzqM2fTG5tEl
hMVKioeJcCZ1g2XzQa/gcqOXn9mJIUS2bUgUltmHMcQrj9M0mTiah+6CjUuH5YKUWuiUfBKIntyU
2z2UbjNat0yskq3ePdN+U3j9pTbC1nWi/bssaMjFuHpjUxGC7V1xIP9XfStwqY1V76h89xWo6pQB
hVNsRFVFx35QHp7MU+IHSsMPRaUQSi8/bNARS/g2EWhTdQ7iqbuKiwo0h68MTpnQPhgy+NwjkEU8
XTILQA3NBP4c1mgr+e4Zqeh/8+K+0E84uhpHa4O77nV/eOw/CKYRhnLayG8YtnlFWVmjaDRJFeEQ
1ynNrNCWnfFeEI/Q0byuirUKmrHDppbGDWReXzxVXanJ72FdKZ+gUBB+CqBlmZPKyUTpuCGa9kJY
fSqYfSZZjQQnrlmdGWYpqqbaZ9MbAUPJqOC/I/m7Xkea8iz5mw2QI2+DyfmOG4MEE5MOGw1LsJS+
bMmvoZC35qD7i3p5T4QMj89s+UkCXOxm9zmRSk3jCsaDv+O1Q7porvODL4diblGM96fTXtIDS4xD
aXUJ4OimU81gboJacD7y00lTdqtZ0JVx2SRroivMjOnSCbHsnL1DPaUi1XQx2VMA9F6H5KLP13R8
yCNuZasFNgAVpBPo2TzLradbopb8EL0BLZMO7Q/E7EtM/5xWv0pT+Juw7qgKe+lKZbyovKDeIkMn
dVn74odLwXsvddqV+mUDcVfaYon/Rp71iDG2FRujak5Mvk6N5+s/5V/6Wx20Y6CDJWt37Nb+BHw0
1x8K6HBE0KfPcdilKtOCLYhx6+50uNR+32zxyJHfaesxOBcbO+OILmvjiMWu4WcXKLHhdar+pEZX
TOS/GzGxPKi3sPTp25t3MBfo+wlWdUp+LkGlB58khRDk3Lyh+IWloj5s5ajv/E0e6hDcunKt7Qy7
pz1/Lq50nrqg2SHh1gGg0OkXjiAmUCasedQhTKnrKAXnDGRbjBcCyx6tH4jHaWz+hbEFGLt98iSs
8Sodmk21j8jloYbdmQJIEwJQFuUQ3u2uMp8zQ9OMRi4FWnXXPRwQTmQ35F7fIaNEYD5zJTHeWuiP
U1T7DWwUeW7Oxz7JEwo7draeS/MDCdKjYnA14I60oFIQgehCfo795+NXVnIq4Ro6MLf96PJORwC2
D68ztGF+C/UwW0Wi5kI5rsjN0cCpRvk6KBSqHadtEBVuJrFmtPvaLTwWTJv91JutboUvEZUJngY0
lOmnpWAZmpBojrtbitdmvRiLbtI5r5HXkMj7ho6D9X9X9n1taa7tC58128Z8xfgQsdYouF+ozfZw
3Bie42k1UzraI4OsPkhj4Iu90M95QC/mqXcfsa5KGdFuRAO1q2Q+KW4ELs+DNiMLHGRcDbXCY9h7
b6TmspC5WOSveEv3XXfXDg8KPk+PPHgMpTwc8FFhnlSMmxQa4bfXxL9Jjmo0HHG/R0MR6uRt5ogI
LUzXa8hWRtAnu+4Wc9HSk3ctbtCYyF+6NooyHC1LtJlVAIhrt0z0jx5HLq36rM5dhb6yQh3tqQMT
wUgptHUewYTzQcJs0CcecYlbs6IXQyuvZlJKi2qFz0+2QZqh9OMRBJcxpGnjutNSTLxDDFUsjLW2
h1gTNveil2ciqBVPMaRDApkfMmaOmk9KED4mh+4PfmilluOEApRgpeGlmWlJ4EyJAhOH1TeLY+xm
7j/OJowG/sZLIVTZk4pIfFgASvnQM3BHQd/vgqGU1oHSA0sCQ2N04l7qWANLKgGHbGQS7O6bpe9o
iIxwMZS5hNt6Opjnk6AFV5drZrgUl8V+AbXzkG5E1ZzfNaudOhtSodEIv7LtzFejRvMMQKF51tZX
uSJAP2cfed0vstY/S56cZx+FXHgubjd243q08lb1A7FtRHyUeJ9EwlQ1eDELbxIdZ1h5F8KV5+KZ
51QDhp6HZalBXcW5rcOKWu9ULfI+qH1XVC7sYGYNDdOYM+rdjOhFrkxwzb1Li1TaMdJ1gHg4rObc
ji7Em47gzmeFN/n/lA6YGmqXG4YI79OCk0jsVkTis5HegKH65QCZmrGG1urM3iXKaNqehnRLqUHE
0A88Lx3iIBy0Q7pnRmE1OMcCbGMufi7hL9OPyC/nX7UzlCgcU/xL/QItB6+Z1wCHYGYaIqifJs23
iPPS0xHalbyOCxLWbttZyryNVfdL7ssXqbC7Luyw/r0RwtxKFJOgf4YhUzarf8pAt10emlmelASb
+iymH9QLgZYc7Q7ZdkfqV2EpDGoxgmFlF6vniTiRpgqlvbU/tQk/5C3hSIDwTbsISIWG7C8rmUPl
0sRHxbDf9hy8VLsSf7J+tNLuUNRiXf/C7SnW4OdaAZNLRdjuJFJDsunfkQ8orsAagJArURQHRUrC
CuZlM41JZQbJBvhncB2ztm/E/lRv8b+o3GVy2Ipev+lJ8qoGuwnvXhoMC60gxGHE/JqMgHtUDBWa
5HM/kLNC4ja+NJXTK0/ab8poec6sWHdda60aGQbNsT8XVV7luOF43eN0HMoBiP+JvB/05wvFVHZD
XiScl+msowU34bNmocSSEYbFvdEOXCof3f+b5IS6mMEO/5gc2LawlZoQk8zSjhG0/ChLGErgvqRB
Bd9cJXjyoZ6BVbFrLeUWtJLYcRbE3od1n8xjIZDA6BkuiWCMiOlbKjG7oUQTtQdr+ikLUbsbGJtT
vipyXfXMcvHtdby1OeRad9QqnSSGZfjRZGvIfmVNLJAzKpqAhtScH/8zaGDONG8yiIfCbgvPzok6
jSViaUEMvdAhj/ZI0YqYCAo+zNEyjUNVsBqsSBEHGAiF3Tgz6pCxfOC2OAZVkoTlZFet2q4bO5d4
LGBJT93r65w+hRpXfoYgz5HIPivsBMRCyOv4zqid8dU180BwlsDT72O6qGGJQuufXFUHfbIfyjaP
Evn8OrDfGa9mx05JWvOA8+loa2Qv5AGhovAMtgtdF8V8g3hg8sosAqet1ZX/vjwHj18qoyVJ+ksZ
YK4xwqlN1IT1Onzo56R6GwrCTAyuCSXb7DFKtZSEn9UHYxt3XB5DCBrLy2mFSt6KAEC/PI5Mdvgm
2UuTjhNKlEvG9RwNQ9OsXosAbgLOtVndM4oK17aIvAjV87aPS+b4Gn864Y1mIwtDpIYAcADXZpj2
VlVbMWTbvWOqoy2j8ouf+3xPVcV41Huoh7ycBsZiPLOQMmUdgfDCkzgDok39p9nc+DqqYScGhOQO
BFrw1KJJDyZ9aOxasCCuAgxoseaOoQbWA9OpC6TD13suRj1MnyBqz14QUca219cnZWM7J0eTfpSW
+p/Tu/CrBvOEH0AEMj98rxhEjzN9n16VVR0ckppkvd82/gbawxgwECevw2VNdPczhOh62XgW+0Fc
RRjQdZVyr51V2OXckr98GIo2ZVvT3xqTxvnXKsX7s8ouau+ApnfJDR9IcRhxY5yxYUuBMESSRuff
CEcrdQmEIHgekWjFKWzjPWxuXcHsou4Jhtp21U+rk8P4iA+/0FReikgYjkKQUv9V1RMoflxzjayk
/sHfVVIcWvowM8tvhB7wrqidiGO43/0SlbpcMp9rlxDfhktidWANCCNn4IIW9yHKl8S3zVD7gke0
aYSXCF4/k01FcomJBwyaWXNOTKIsosbG2+YNbC5PlQ25BhOyJ/c1FjmR54qkgnfMY/di38r4JOyk
AiL9jdwFmiOuUJ+z9snkKUV0u6CsxZSUIKqp3olzPLxahBmGIjbtjPPnRFV/IV+savUvXqbGSEgb
rHxc/2aEfAJfTDwFNs4aWSz6Bor7LcLusRb4ppwOLbH0jWNJ7SY46Lfizc9TvZ3iyYZd5Kca3m/b
J7JYgQ22ikjNe4JEtg9ISGXavhq9liHa44NztpX4tQ3dydD08lTyArZkbMsXrwzGw35FZJ7goDNU
rC2O9cLcMNrZCADQQM1z4kCVa8o4OvYEtQr3yItyNN80B/lYs1YJ9G+Uk7dbxMgr1XBo/x0nSp8x
SrPAIuqxRUpq9WLFMKmYZXCOznARU5g+m77j+v8QuZP59jeZaTJ4m6xN82XiGUD4qZB0ckzapRkK
Vpduznxguj/D+yxl3f50dEt5hb6HDklvXo2U68wq0janXb6qjAIulBD/VoYicejcQtMxr94kky1e
fIr15QFoHU2S7qWqVVpuB4ocQhKjmnTO093HQuETs/ZB9jTuKyGwahIjHQW6QLnkqPjjeq4D8sKW
qYoIiStUsyrpS8cQfL29dPvOyL2xpEv++fsEaOQqxD4MR+9Ze9S9yrFUFsztx5ZBp3L7JBk6zH3M
VYoj7FtV5cLmNPmEFruMKkucYRLio7ksw9gFxpWRvKwZPVPf8aANDGK7LNSD9618z3cO1nXWW6wI
8UjipjWKAfvGEwPUkgFDzd2AZ6tIJ6L1q/loXkB6XTcjIVygOLrIyYCITK9fBghYrjJL2pwzJ0NJ
Tco+xRjZ3QVmNBG2XvbsIiFrNaT26tnYOxhF8JxXw2IzizMpqloSAqvxACwvqABWoqQ+ixGCSoz3
SCNsnO+BKAnKIQKWfUQoJAfuAiAU4/owWokZGHa50dJVKjdHx2xp/9XqYY4LeHj+YIcTaeEsKP9b
J5d1M1NPrlT4HLNDuWlvs01Onlp4h7srOd6RFZoO2Z1wmQeqWIeGNPKUE+OUeL6ZPhcG/qRiW3B1
6d7XiZyjzKiiY2L9AlUHhG/YmQ89f24dRBZVLHtb41f19z+9a4g3msvlPPf1BqDVNksMQbkzXC0C
GcNvpFFQhlHAavTFjkLYqHGVMXF4+Ml8SwV9Yr960fsg5U5XUfR/QGC3Zw5T0ByDu6KRAA11orzh
c8sg06L2yNH/8x3uJzDkZwamN7+H5nHapDJlbMQ3WPLOivbmKLabtuQmKe7zUVXd5XiNdtayqKPs
P0vlC8nbxOYFYcd2GwDKImk1BlmxgimjEdKP2KDHLAHvGmXdn0D2GUBiyqsE1hN+zTHGYMGQh361
H6sptgr0yFlfI1nyniVY8L31mfjLGgItgHolXYsb8pDKFOjQBnAFvJ96Kb5CKUNALTHHyNuQJwwY
Yt1CETE6CKn/HTXAI3Lfr+M5NSg0E4coqt8MVHN+E7JGIJbaT9l+2Z47f76QANZU4CMWqXOoPXph
kOySuCgufWSz3bEruOCcMljV2lIWEkjp10ZVE7wOjpqq5KWPVAFR+y8uFpLeOIEgOtVfdtqOfhje
y/dDZ0kGuvRB264j7K38mnKNMyBWBZh1imjabeG7j7rAFtlWcknTnBkuaxeLxPb12/tbSQ6S5N8e
S7QChCEhfahV/7kX6Lrht+VDTT1Paq8Xlg5CbU733u/ZhpsGrXvkTo2NW07rcz6/4ZUqBIPvsdrX
3D+hTXSNMNQcH5+QKRuA9GQeg4TWpvJkol6i8yPugQwNBqB03hVjDzsnAPqCi3GuL7Sgs4iHgmfu
n8c5a1Ukv7qtSVZj7v1Zqe76eLfhA8A5XwXniAkMzXCfG18Xxl50Nx3bv0Jje8X/mgl87lz3j6oZ
bXGGTkRFC2M1410QPdEiR6FFO4GcBYero4nyKc/dKzZLwqrmOpy/wwKYB81Ujq+S428CkBER7XT8
ktnPt24ZMhZguIJEWyLWnwAHqTUh4d2YkKc05e4XQAlk5lab3+3ToRVLeRSEhRvsalK//1WKxg+w
kddTbEQY4VJV1rA6TVOcx4xBHiuddCELVF2tMpVQZztjbrP1OBWRIqmIEOha4lKr4K1FBxjNSszC
fjPvYdFEexmp+ZzMqtuuGSLH37vhSL7deH0s9gJMNpO7WJnnNljdfEwK/xoZG49NdSCmmhknC51r
eTAPb0KirjPVkcATiD1wqRcrCEotL+1im+oWtoTEtHHsjUsl0sneSzJV0a1jQg31mRfHDI1ercyN
cQ76r3G4Q1k6svy0kPt9X5Q/U5/jEtSHUQcw93q9UIthFAqfDK0xe+vjwNoD0PoPrLKXIX0JxThj
ZXZsYzus6wrL0qyz2NoBaUXeAISQy6u/q44uxiq1UFHsW/CmB52pHTjUyRguzGaCRxbOjP95Pd1O
VMW7nmJXrbMhSP6yCTSRUcts42DbZaliS5VxgqlKweYQkM3FyurbGb4MCOWN/CRveSDV2W0Xd9TB
DaK4xWblQR3k9a/XHypOA1Y+EKR8qeBetZn64oC0NH8om57kXpKo21X1LP5U9uv7ptiwc97zphVg
5VjyImi9BaDE9wD8xg3df7fvZpgE944lVWkcpMtr/+XIKRs/DYS87iQsCchd2xitSR7awcipZksV
2cpa8iHwGxcrDOlbJK+uIk1aUV8vjH181qP+JkIJfu3bg9ZehACvSI/SwFSUhc+WWDGAyblYRy8b
4t2aQIf9aqTsgygZx4TBzs72Q8utpeOyKkZ0/cIOJ9sQsdkzM/EoZDGpQ48UFSClUFej5rncnmHo
oB3TIUPOPWFoJBdKPvq7MWWTZoujaI5WkcCHpXxfmlycYYDx4ZzTSU9bOtxJySmZfRYsVzqJbUwh
OQctzscXTqk8K7VyeNrhqKEVdXQa40oYSWD8zmO6KtghvGQ0YeSQl2iqSyHDsNoRPvm/rs14KXJH
syaiYa81XIqwOq/G5PZTbOjF+VzVbFBwYETm6cy7DAOxHNNzKnvPrYNhN2AJ981z8A5xZhKBKkt4
UBtqdHxUgXOj6GE+4F8qzXyozYNVNeD2B2XZNrX8Cr+3czZJGe2WNaKd0cF+n/ox5KNnqDQG55dg
bJaIlCaW5aacjDNvANWr4eFyWmFT6IyIFMdjUsUmtECQb4vD3WV6uC94UWMZ6fNISRCF7BVZVcom
oXF7X0jpMHIiXFjKqImEG01AUcVuBexSH/UCt8Ay6TdEtq+sfOYC6qrLzCQN7e04/5wzkEQ/3gFT
hpBjj4FSO4QVl+WT2tydBaLRVZcwv2n13/4j/yrArTFu9TPY6ALp8vCBeu92DQjbFKcK6PcY7BO3
BJVV81wNGxEWBSRMfKrnJ1aHdWhkXACu70fSzLcoxD8UWEwmVNMPlRAmlVzY7R/RAfGscKbnz+sF
eneeGsftU9gfodkGmQ7Ep+BQIQv+95a25gh3DGe13K3qDm9k71AGy90jyZ+BxZmB+qtNerOH39IQ
uDsEQ+VqKHJUvj5gdPbpJYL6nMncNAXYUmztEB0KiVWOSF8jD2iEmIgGOA5rWjHvmHmNBI8tcgOm
zEAFzuQF8LZHLOCjA9u78POqZSdp0t+xSskQZSri1oMa0kxe9IiQ+g2HTdFC3qezA02yLjOtY/yl
fYzSVTBaebyfYfkfqOlJI5v7CL+D9l+gk6DqeQc3vzaS8PMhgmHsb8ITXKrfJYodkof2FrzupRSp
KVQZ87BNIYv104sSF1LfuxXaAUHqxpiNokcHjxlvjxnEXDKMEtm8TvfSiqDBYfgcOl8zsi9jWk4o
Ja0bROdkEC7xT/tDEWLy7q4bi2lbMxrCgZng5CVjOmFuBicbSgetX0E5ASNsaxA+UbpxtBc++u7k
vYv297cFjOWY0Ei3B749x2KG9Zs3ZRjD/YWe2wB1gWGGZ55NvMTmEuxy01y/ULdXrOHNfjKXbYYR
KIYYHD0j6WbnU5NNmpCQio4eIJlqQQjxhHOHnn/UFSrR1o6II1YG9S2wYnZwaUfggtTU3XOExcj/
zayMWMFMb6VWXd75XeL4jdL/78yIcnuMRz3IdsY+OpnUdjlS1v5lXgv7p7lwpYN8hF2KWMdyccWR
72X0s4wTkd+C7D80D8YeBg5RJUuJKtb433RVokH0i+ca5lh0WzEmyziqTgzdokxVuCIdSyqj5uTS
/r65X4aViwYNkFgPOse62EXAzxRwyeWLVFVNmIgxM1hvdtsiu5KFzKdJoP+HNRFdop/0rPkUW5Fo
bncMDZGIVBiTxbHc5IFigo1dGnMNoeAENXcg5N4bPJRc8vITjzb089zRuoFUw/FlFe9iCF/tqQa0
0GtlhCvmmFd7KADEW0s/ncaMFUt7dXS59LNB0obeqxspcAJwAIZKxoAsYBcFUt0EbJdp2BDxzyIS
omXrQPLNyGfHet3+WWGag19Gw4kX+YM7Fz6/OY6m1ZxWsC7t44KSk7DocTjuWCoaHOnbr1NqTf4/
qLwnCW6C7FW/zrknGIenHLrPfjQ4kjkiO0fekXCek2FJYFn78TzIG3HIi4LCCt+QkCeLCRxGd4M7
wyfs9lu3nkgIymKmdzYcemqWpLbME5+mAUEyZsHuSP9Gplv1sjBUJIVq3Hf6HgWolTUOfRT5nVel
6miJqot/4A4p/8Y6SvnsyMaXII1Q3Jm7Q7QAYATgbiakchkGcfwgj5NuJY9uyNGEp8O5hCslD3V+
2p+l+tvwLuaoLEeaxrllRmwvVPsQ/OwuYZ+oSuKXbA9yVqz0T6H5NMdMU/vGoFTBWDSFALkfpstD
K7CAeIOXSC5Onzg4nnov2BhDI305iZyX9nMZAVRykuBCJUieAjuD2OzCIOjRM34VVX8VmH7CUDZi
9x+qW5plbsbiuj1jpcXCLabcrGAXxzvzjT2kpDg2HRNdrCoUFQ4crf+AQgB3nexHBNLdEiOzl5Jf
Y1y1LN8WB6hPo9JALxPJ0omYMSBH8O6sJCwgw4wRlFz4k7Y7nB4nkhCxSzzPYeFMWPfu1aVXihw4
KeAwn3v50GYKvnh03hmE4FkQ1CVchtQGkPRGJN33FTfSynyw4Jh435GUSPfdPmLjiNsK2ltpMHLd
E2fCVHxnzCfUg6CAwDF8KXVwuwQZMMxPLyVxpZqYqgqzmWhJV07kbFM6+PdeCCXoWly3jUUjdw+b
s6q90hPOd+5oTphnEwsomNXR5QuS4fQEVjcAgudr4tyamvqRtqKm1VPGLDzyTu1nak1AwEHeEyVT
BP6rRLbaZzrpZ5at0VCs3liUwzjV4zGcTQHERbg2yX7cLFN/Wi2+qt/l2eDWGjYQhaoEErw/pPEd
Jy0uVoy5Au8G4HIlJ/Vaof89acMlK5+5BSGGWBRaxXvLroEvMwg6ULAHD75pbY7RJ7FiuuBY2aVZ
YLVH61jQ0iEyx1doRRtREUimMA2quQtXvQUmc6GwPSakAtU3M0/ffMteoHWsJgVMdItIvaifQVfj
y4Ll2MWm2sE0QiM4FLyMBllZSjtqhwZjPaGTt+o8uzQIHK+66LNQlTC9gZUa1YK2wjy4Ie8ZMUeZ
vxKi2ANjeM8vKT3hwPhgi6ip0BaEH3QiERIk18dBSRS0epVqm+KF6jnd3+VXGdaBozk3cIgNVbHa
DpWIxv/dkopoAj8s5u02DwRvz6Vr9g9mvRSKBIV85kxOHJo78MAKbLoiF8lJDhb18E/Iu4zbW3lJ
IoxM92prafuO/7Ew6W6AR2rvjZqdAGOtLz0v1B7uccS005SuTRa2i4s6L/j/1uJkOqQCzSc7TDUV
v7uxOu907LHornBCrId6Ye7/5946ZC4/yldDkEdw6wXWWRAmVsuyLYnj/K+Nr1o4NOibSaqFgU4G
45iF+yVAUrd6QFS/lwM0avv4xoJeawFEN7Qm45PEUzjvxBP+xH0bZGM9TBDnjZtOVrrsjFz71QOG
GbZJ9MAFT2/ilU7hDqrB1bm0rZ3rH65WlNVDl8QHd+iFhESajw+zEAVH9LwIJxJcEuBkzTr8aKxq
1+gWXRnRZTfpLD5rGiHT/mVDNO9N0eJGu5bJrKaN2tc/ye3WqKD+mMHWdyIdHopcgLe89C1aQArp
BvYWk23KIeuGXDCU7oaImusDcAXF5yUpLMqxkMUzsyWnLQqvUm5E6XZNSR6ZDM708dOy/755vHzN
VXu1kWVb7RP/JW7HBDO47nG3U/5LrE8fERY8yv8dPp32ivviuhUnmE3NQ60em0cGvMF7qNMh8wG8
MmfGhNuAfdJA8AvXCzDkhklB7B7Uekec/y6G9jQKF7d3QqMiiiAXyh3zCmofELUG48nSAyAabthe
Opa2tyWsUCboMjrqzBzTZRS6q0yOuAVIq+nwwcm7dDJq7VruhewGqFyn85+AoN7Ncx9BuH0coEdE
Z65QwCnEno32yqVBkV+3943A6TsH/9K5QYOZwfYAjmCgGwiF+YPrE5AHCeAiQ66o3A5B3+yCdD5H
RFHdf2KoT7htew1zOOvAVaVyQPsYSF13ynNI4rxp8UQo1J2EJdqh1JQjk8jh3Zu1O7JJUpWy4P+E
3f1ipwiBjxSSY8LbQt8JuRCaXtFuv25nayO7LwFm9owCuVkKrOFqHCSUtcMb1GVe+5RD2zFSWAfC
BNpHHHevKCYAaI+5tJkLER1vYJUeRAE/X9srCB5NJv7CvK+tN3gD7iPR7REKnfWxKdAUTLPd3qzv
sITfJ4KUjOfyAw5q5B0nr/q9ZYKhMyGd/Dk3g0hsKDtmi5d2wvr4C4SC1ZFhdU98XXGtAf/TrWbo
tt68+OOBhv5YmHSJATkxgE/AJNhXA3UwMSjzc+8mbP2S4oRjQ6uuGQunJQTQ08fM1XtxJqEnUTI8
gLysyZBVdKauxerVChpOZw+Vp8qIi9n4Ji3zU+eP879xzT6h769ukrWetsiWLSSEiMYR2GVrywGg
8eWgNAkjwXKhzek1DxW8f4M5oNqAma53hgOFHdZ7xtHpBx0NOWtUrKGEJ7L+jzsf7qotOKEH6e6p
c4HaEl6nFYVAMRbGF9kV5b0NzT95AC7j5ZolQUUACIMS+0Hl4+qolVHPChO3QXgIdWJwjapdQZFd
qxWp6c3Qze0993+P65ujaNo8VvctN/Cc+/INQ8HiNLHW9cmfIXaVQNSsyyfXq9AViU3tbR4BBhdK
QXmlgVTDBHXMpLZK+QSXU9ZuQobXikn4O2Yav+rSBceTCwQ09w+/Gkqe90cyEHUzW8D4MHzQZHEL
sEoEqLU5Kj8wOw+SKArsnzIkorgxWB90/mB8axb5/OiPXkdU/SduhRRLUcTyrxa2VOc8GhnJiD3e
AdwOHitPta3K++09GuQNxsqRPz6oHxTl2GgdNvLLD7j6JbyqECLXrbq2wQtlgQe5dHM52GtuKs/w
VfAJGZ4brEHubE+IbcLt/yTTd2ra1gIatrQNADZWhXECGfxBcFoD5u71a5xA8wwNt4iMFD7nvCei
wTcJwgXiCsUP1iitpqvVfFRQ/Wy4vrm/vtj04Mf2LenklllUYj1N51b3C+rcKFbTj6s+3csZj4BE
fKCPvyA22u+hjCQcuG8irP5twHdlHTbHpBjghl4fXOtiUkHTLaB9FDazjWlEfAGWBh0eB1psb2E3
0NFUskTP/muwxuuvZKFULCQ7R9+9Z+DtybKvoRG3YxhKq4xWEuemJfzg+92nS49RqQFAjcksrH8A
FmbFx1tdEg/7Vh2hRHPelSy5uyJw8d5urA2cuKKswY6+aDZWYFowr299txjWXURtJtueQ9kimiLs
Bz0WuF3k2Id3b2ag7fesr0i1J07CnY1q0iTJnfpvHpX5TYuwY5QDJDcYxcoJny66xVPThu9Z9idx
mhXwOm/Iwp9/pg3iaTmiQpfOSSy8oJBBLq7r7OcLlxlFtYuVevcErBGzvW6mGOgvQMTjYte94QHk
NNf6gWA/1Y8RPtRWNdLS0Wmt1BG9Z9I6n0UfgWeQpbKDB3W5zBtY6aepdluEjABcfItB3IucbmHK
pInACQufPHjPCHy7oiUyvCqHluwXnBUZp+Q2jfdlVSsBqAyZegL62huxpVBl0LGNh3F3JAmV7d6e
X4WCjNBLOBvHv3NupM7/PzmqvfyxxLy10O0JxkWwvREkSQKJj232SlAPeVMwFKp4/G4vvnWAPgVL
QFBW62OTDWRNDxRQqSL40Z7ndbwVDuXDSsrIddBQDLQGj2vhSnV+CFVIF2jy+SKWSl2ljM4wOa5M
AnIc6gjqRFvB4cUeI2lj6izBxvGQJAn9x4J+GtobZNNDFB6mXzy6fYqi5LjlE217mc6Ot1ILNL+5
0LcUplsUC8ulDLBAO6iSb8firB6IaTXliBtIxIDavlKDcEZwnaOqBwFh7gmhBXLVnz82zTpUPaMM
VpqEWYyPxNWEnYqT/CY3nPe/O5Cjqnuc1ixXE5RrikjaAhcCa22+pV7flo6MRqIuDMG2qKXog/qs
J0s0NFB9U+GvPBNQHGJXI6/xgxiHCxqZxuJMkHg5hP4rccLxTlE3UGJgUYuMvizRBFGPqHAICcxh
HMhLazuRou2phEWNN5B3aTZbu9HkC1PLi6UyGT+AbOZxBOzv+HPsytiP3W8BLzuReqicSLNGXYRv
jR1gzGus2WZZd59krcVIsQynJ75TdCh6eVpGZyh4RQyEzASOWnuw5PJBmkAL22ZSC7mHqHzEN7OS
nqWjNJnPobTmBR4xOZSHN2T73xg56msLpVHg9YuFy6mCNj53Z4pw+dZIN8id89gejjQ6f6Fog4zE
UBP9n6MrW9UB2Cfwo+ZjBUpfssw+Vuk0kjUY3BiVLrox0EAZLWjePIAoRopMvTdYQc0Xa3JcGR0a
EZsWr7NTjpedQ0dUuIkIygBRsqt21lqWMsEzOgXdVI9oRwYlZn4RDQOhHAG3ju+XdwoJ3NwLOaN+
QYyyqFJjE3OUZkwzXqcfVPOgBCsNeqnYTE3+XL4O0rsNkU4of0O2JqcZcjnTJI58Tl2ESJ1ajitF
8jV4oh9GCmUY9G1Is5yrR25ImUgmnX1GyisXu1hvUbsgyroHOhbcyDWnLVTFiYj96nAgCaZ30YBV
ysOUpWW7ZuoXNEwZ032yUiZ8Q3LaLXgShgLIAYPISMwq7DpvHU4L6pQweDNlt51atMt6L+QeVS4Q
67FmSISsiqfW0qKWmBBv8gp5wEi9XioMstAzWmZaq2LX3WHc41odGqhOC0z9780ePxWgnJJLADFv
bDMPU0JdqiKdjpHfAylECCEBT4TorWrWL2XyC3XsVuSvr1rU5KzUf9Dwc4cWEzNYEQRmyK5HqG8C
ZpxsXtEyKQ7wHzfNe0V8x///is9fpjuzqLDFBdlBTAHISU/rD6d1PeeRjhtJ2y3hp/0KgFXbaXQ0
0lRLuxkmtvoS8IwA1yDTOv04zZDJE6nJRLr9FPWxwBpheoqauYPBfbxQdva9GJFGxU0bh2fhorkf
I8f246WqQ7aLnQhV26nRDzg4u/MxQO2i3w5R2dJaeK32mlHLb3omlAInfncLU/ssQUAKHs4YzmEF
fPynHkNUUW0FJK5TCq15clDvdh8vhJA320deIiPEHeKISUhIcBMD6gXfxA2baGFTRbbf0IzodTKd
K2hABS1L7wGe88b1L8kRi3xp5dY40h48+e3xnfp5kl9FwQ9aeaiW6XDz68cGgL9isdOblHLatlwy
uMkTLqdFIgCfgStHanBQ8nWjA1e0dYD7PwJB0YarZAMQYn5FWqURjRPf8hND4sFDoWnMC8Oa4voD
fcxwiSj+ZErSiRshAQs5mBghLo1cNh0/eS9OfpLa9xdFq17hU/iAkb2azsYJ6v0kMX3HpxjNERHI
g1NrR114T9z/no1pn6X33fpfXmKsgK1GWYElmiUB0v4eQUZ8fmcGnzUKc/6Sn2LzwClQScvkXWhT
jW08T83RcnfiM0PqtZoB8w5LEcDnGIpZX47Y6Bi+FOq8IbU+0ZtXqv32n3ZzinU9pFxN8euX7830
ipbmbmZKi0w73e5ueX0g7CZANcWP4DfWh1JTfzQIpv3BdZQ6xMCE3tmSMSMGffL27HLV2RRlgT/5
cZmBV4KoKLpU1i4Iaxvd0aR3KjPu0tOlCbFJHmUL3VsEcOPxc7VKhCo3p+mS7ccUqo8I8kjWW1We
RHIrGpcCNgoT0JXu6fLmjem42vl6pejF8tFBKRTWw3laduU81NgIdZFjmCxVHr2V8wxGtPp5fCar
JffU3KzJ62M/RNLA6Z24+bBGFYdxbbufKc3cIUo6P1NWVKggsjJDWTxEnFAd6zwvoymdGxqaZ0Qc
+c0e3v4Fykeg5uXGUI4MU1qxuk9sjlapY0jvAWp+PcoMLS1ahsYQ0grxC2igT3dLAM1Rn3KPNx31
75AmidgwcuPiLrS3qaIWMlh7HN+ImlcyF3kHKmcVgyHqPbyz1FhJ72GCywXHjzTkf4jvr6sFYJhL
e04+lfsmpKq28NZsXdb3x6aDoYyC/dZyxgNQqYOx7sQ/if4Iz5dinmDcPkNO+XTJe7arvWGq2BsM
sLmWxjouONi28h2QYxCGA+xF4gt/Rv+PVPVbcuGrHUQUz4I7wSFoCjVtFC0C4bt+zVFIWjp3wtpC
N9Xnc+6zNEiGfIWhD0OR78FvnyJ09/yivWAAfW0xJrhG2prieSodMtMQniNKyigL8rHTrUcE1Glr
n3Md3Ip7EbJPUple09TuwCjy+hNGXH9NrmuREK/I1JIth333q1KPi4Y68R78acAL/XtHj/lQ0z1o
HWuAu1Thfnx6RfWfu8i75pHlMtql/8bf6+643zZmlCSR3eZtHb3sKKavCu03+gE7DsfUKohXsmpy
03FGDtxzBqUqBEkKcw13FJ54KBAO9GR6AG3jzyeuP5nzVU4mrHFT5g7TdDF4UtjyCs2awl0v7IWX
Gop+GCPz6B3SxXRn+m2mlReLYhjNuXzS2SLcPXHZfQLhum8rJ5NT1Y3QpTVLvz5zH32TCyCWPKI/
F9sBC5UAaev3U2q9/n2g8bf+Y1ajcP0zVmeUCd0o/7gaV6SVmaQQTT6UEy6KF/uRNCEMWdMhO8Xi
5ShmKOm0svT1RiyOtJePRmv8CcJ1h+/l4kTHsPfeM7pwYcq7+x53sVMJFET5eoucE0ebWASjvK6j
pQAIyXSEly0iq7SYFr6yFGca6ApnMMm8SXC5ImYFGebrqHS+sG/x2odQPCQDr2l7pR/buDyjA1/o
x63vr5W5VShfI/JS8cwo26FUAg2HjKwNBxNaq8Gs9vwMKRSSy1BWd/43/EFKVY3uUDLjJrYgTDJn
9tM6VbYYD3+JMmzwyTAl9b9c6zFD0SccmVfS4pwkzzOWumyy7E0PQMXWM3GHa6bkpin7C77wMA13
SgyRKS/voflC9Dmti3WzpuN9+HwI3frK8xZImlUg4pb9QyH7UwK49twmBfF/aWzlprrzX5x6srRy
ZL+aV6CkMcnBrav7IDjNNyIdUZNmSL8ILm3+W5asOgqog5DsGP0a/4LaUytz4X73i662i4iATGZo
AVeAwCvNElaWdcf1icRH+Wn6ssexSpf3cOKaoMDOr+ra0/Ga3RZHAooNTTVdZ5vmvl0ovtNP6DjV
3dH32BeO7c3ooZVxivqhmb1EmFQkyVA/GPeK/VjNeicTCtEpYYbR6S4Gql8cNdVAXW8keVHpqYPa
Ktm6dLB7EzAJkBmjI9O+vuxQJZDZNW4BbhI0WBEBBmp68kElTtTt4EVLPweMOF7riHbenIvksHfc
ip7ZWgJM3DSNY+21QSLa0WXWKNyic3iQTI/OvYyNT7XpPJ8JZT3TYEXzb6bhonVhV0HZ/+PixHl1
hH/Ckr6ZKntOQkTsG5VNiS+kUcPuXZOsfNFV60EKk3ve5TBP5iXhXqW0p4ICMRpX7VVdKATbjMGR
fseApYOLDlbx/FzQxg9qsrCpnNg/6ZPOcSmaqnhr5aw+21zntszW7i2tLYzi6e5SySprOC7xPMuX
B9AWXHqh3sCmpPYlk+wz2onDJzVK9d4O1Wnys29sSqF/VplDQcorsUTxLJ7/TQNX1QQ/scPYPRVT
gs8CCbfmLtUJ/4iGKoN6pfrqrg2dPqAG8I1sAN51Rnfe61EMbKHM6DCm53d9WLXd8Qj897P9XouT
JEH7+wyEtBFv+fFxhdbfe5FyL82zZ3Dw/eWryH2F4HWQqMy9qbqZv5NfTuVw/At+B1ImTHsoE6J+
agNOcmePQBF//KJuShz+F+MFo1hmoPFioHulDQ007X82fIvxCUwk23K1h+lJwjlM1dQsA8ViR2OF
fVjndTSOwtjMNJhBZOz/Mej88MPQOAP3/o2fhKPVop2KUE7dA8SV1n+w1LqjRoDVs3XEaRh0pcha
yB6UQXsBreSz15BEjKl7sUhgryg9yC5zLJyxfWgovrDSymI5fCg7tJbrQlUqjC29fgR30PJGJIPn
G3md/5M8i7DEsTcAr8dQTpjn3LB5rvaTLoJe0of8JysoECpWQQwsswrvAJ9RiZqW9+3682f0/5Pa
PCbT1JX+MAKhqt6VfKioMSZVrW7iF+6r05nwuM70utHxJUnxpcs4s0NAyJ5+5eeBK37RuvFciBSJ
xtJ3KV87a7sYqKzWwRWUY2lNF7cplehdM4Qxh2Awic2dqwcLS5zNYop7VKqWeqkwT2YohBWYCip4
CEmmvY+LciYmmIQo5bqyR27NyQnMCRdah6KVeYMd0VxPM4eIbkR9uknJGtQ/XsOPIeSV9SPr/gTp
vj3mGTKHk+N40O0+uLW+3yfh4+No0bZuxQYQ2AYcqdLrbh5oIDjl8idBDUJW3uy5XJ5xcoul12m6
3rQD6YzC/FDgcC1FkF6gFVG+m9ZnlJ9ACxEor4YNSJF7CSgTI/or00lpk31j3Aj3eULrX8rivqAM
Z2qXn/CrVSNd/jSmSUh2Pp+LdLE3FOZTK76i5HOzijStu4XuGESMkblwrFHxjxu0GVmJWpvrzpca
h+h0/cfK7DKuTndC1zY3M8y99Y5awlScMggZRHEnQQDRLMML29jkga4ycK0QVs3i0TjaqenYOdf/
ejwMH6pgdpFq2Ml9VAbXEqg+UEaWhXrJSU0ApjpGwH3lkc1rQIt2UphofC31qjTuMg+xSo/UIjFc
/5X2YJAMO5xtWJSM3hPoDAhc8+S/IUnXbgbNhoMgvuvUXPlfdpMT3pitRGpjPDpMVXhyTVJfsYIu
CMMBOt1ULCchzPiL3HYaEMFuv2lfQ8jxnN3c1rWn8/4TdZIU3gwYaquPfBRIOzuezyoGoDZizp9Z
5ZpVvb+11Ebg5KdOE84g0Fko7gZOwcF4H2LCZrVY6YZzonMCfbPhzc/OPZBxH0BKe+VLhgtR2691
5Vn0Qu+t6MLm9eyIaDBoQrEew/3FNrqidWaNbHxdqu6XRTePHq/ra9N0KeA2s1h68rLbB9wVV15x
lUf007S6+PI8Cr/KqGO6g5KiGQOq0aVLmk0668zAdxpUTbUp0kmteYoUe6l74l9UP1jhICUDZIzz
4WHRUzIoCB5n05SJw2QjqESaYPLT9rK4XTzsE4srVB0AqllmEPsRmTvuo9mPlV3+ynEUeSZovqpu
b2EVQShX4pBZkSDtqeVReAbJMrJF0yfWVhFl+YcZ0kGe1lUHXGTJkK+I5jICLZTb9d3p3cHkjUBJ
K+p6fRTOY6fy2vWN6aPT4tupcJbnFkXG6nwwQBygIPnqcCHo+slQuxS62bk4nQ9UwgRPrBA9z30n
ardevh8uZBdTNVnR4SR6qEsEtzlDcIA9yuuWpzc0naKYOj1/SpcSixSsaCCD4ibSlSssbyoUuoyJ
MMLVWqrNaBPTQsRYrm6WKSwWenDSya2oQYLBvHEKm0jtCAT0sKNruGcuiMHw/Esez2w0ZjnWOR0o
yoomcmqY2eA81gGvWg4MTd6lIYK/RFv4gKPaLXu98FmowrrmQmuAZGmGz9bQqh4IB0y1GsD1zNyD
SNpFUGg9mMDZ1J7jEq/nsiIBzvkxOIGyj/RA8b/BQNsiTMCBFyjNFw5853x2cN8HOcx/ueG/pZPF
kjEZ0m74tr/Ta70J2zO1GQVyRX60q6V27dBrpXGnPSv67HW60sjcLyxlweEqEIxG5QCxeYZedgSK
rAeZJclwoIOjZs64qtUos98nnBPIjZ3daSBQ+x/NZzLg72tCbDryGVeIPh3FUdVKhbyj3hFm3HdM
t+MLOUh+C0uKmc9cEta0fvoqCPHwasnxfJcDqwXJW0PqN0iQezYQfJJ1KW1+Aw8Ay06ZQ4WOTi5/
REwDOqbG4TAYm33gzTQs2XjnYLLtyGQ5cySsHvFhHwySnWAeBeU/rOfT7fZZb+dK6RA2RrMLWjiO
/UNtt8wpWFwU6w3+M4aPSXkNpivd+8sBULHUyJxDRz54TkWnZMetJ85Fjo1wmV8nJrAV09JPxqBj
uGHnG5YGW/FyYiZUGDXt5Cq4vKGPBitHHcC8Tw/NhUAu0CQpzyBTlofm4kmgzVul2YoF7Z/7FPb+
/04vgT5dsGlIL/hTgF+BtdNoySUR26v1HpR3FEMCeVPNdmhdhC3UvuAdJfcf3ljI9t8sdPhRaztQ
qJdRyKkucwNPXE/Uq5KajctyxhOD7TkhStH8guZ3dlauOSa+E9TdB1MhAF6etSDOCekQ/pj4v3qx
3LHu6++oidTIwx8Vy9aXvF1Y9tEii5panZ1Q9iL186LRRjf/iEunWJmBf+oZPcVI1csOnf4zbbuv
vNnj7W8J0dLHCMcczTi//jjKqiPHWmBzvHiORUbtmhs65QiK817efzEsAzxhHc5pYgWgrPNdv/5/
j0cP5zpJB7Q+uLXKIHPy2j8yDOld6iI1d1tAumRC11BWh814KpGj7ntIqLtucx6OGdqG5HaaAvIF
hd1d3TbhDrtsGutcIpjs+tDkozFrqjnfw540CiUDsAZfGblzmztkM/LOkfor6bkR9lp+maI2tmv6
NSKQ8hGhRU/p/N8NE9JKOa/oHjKsghD72UJjQbftqObqDkCIfjNSLSNTMEfZ+QZF3bWfgx/Avhul
du7uXgVqhZO/g/5mdr9qMJF7prAz8mc/v3fS7KaeG4EaiYcUNpZvokdumQjO1NApG8MTKXW//pIj
WKtYN5qTj7pikuNhOCsEXahJOsq7P5H6KJXUDpr3z6ThjIpFjbR8TSspmiQpirV2UVpezKbxR20P
tjW0dajW81rjogr/CDHRZwjN4q4qOCVhh/dVsNi98i/KnvgU6gD002u3gaZUgjau7NxkFMsKsRQ2
jYAXFxznrpZaoVnl+swryR+xAV/CUVU99cCYm90WFvxX/dlm7T/Go4W6njGx4CCNRZHaDrhwMi29
kzhuFr50yi58RiOlnTC6dpHB72EXbcjhjSxtHBS4NuNVyIwc0xab6sFgeAWPM2Y4opPuLOLns34U
h/n4hOWjPPxwDPyp1QyjHFOt/n8mI0+0zQftf1MY1+QJVipjIv/bJmzshAU+ZWxfT1rW4C7K/ljN
giGTd0xN4Bxo3VXTTQg1Lf3kdHcXp9318plvSkMweMt9SKZsK5fLxC6WjINJvIwnlVTdzgEl6aFy
vsOsNjmk3q/hN3KlrWKkeviqi6U+wBTf7Ci/QlxDeWZpDeonAbA2W08+I3IWmGpZRJD2yGaCTrp7
BjK6DVZbN6FiCdKZQxXWc1QcnXCETJzmbLJlPINSlTrmRXvPPsxkOoK3FItLTb9wq8pAPXvB8Yi6
KbAvN//w4QANvikRItvAEFFw5UTbIyrTzlur7mfMnxW2FvPmXDaZXCdp+mHzZrzoNBBH3SANgzM0
4CvkJUM5e5HEgUpsjaVFn/DCWpeBMRMsafVOK1c3f3a6L2SD9FmGLGp8RcJwZ9QxzVTM2nL8TMIW
mIGdBmVRRdepLshUrQb+nZefwKQ7Tn4G/IBnpVBUFn1wTU7KpmMbZnPFUHz8MkIlBMdwLUQycNUR
ul1GGmjG/dOABRa80ijmrn0JqSv3WCUwKr0WYxLmA+DEIix2B7cwx3yDYulDikCk6bt0PtJ70sn8
obrWhllXiU8p5PtUdMpF9msXnp4HEZ5K315wlSZvZLPzMd3GZtyWffG/wZVn89iGAgh9bJH4KTPy
vUzD3z+T/lYpXkOMgT/SiQlk3I5SY6pjOigvz2rlhGVdscZr1Hg0ugNBRdFhEFxChtwgF9hX+Zc7
QOC8dcWMGS84RgHXTL614rtMic6cj0MF2ijrvMrugY67wKuZMIvlbrGCSSneFK5tBQV9xaa5Bl7c
Ap8aKyI/DgEFKwvFk13dN3f5Hc/MymWe50dCgiYQheVAzWzYjt40gSwuqWvPk8KUV/1YhnbLEWMm
SuBC1kGiVAOSLk1CRGX35wPgemOdM+Xo8BHI7JOL9R9yNSMmgH1+Ix8C+hVGxfIbMDWw0SN0aPts
5zLKhk1rNtvzDP9y1WyHuU3gUz8tXMU+R12UnzJuEeICBsFNGkTg3/43BL9L1XzbCaqePP7VVjfR
aKHnOerlJvD8HY7gmGKoR3gOdUsQkDfCmS+TtbaiKOEr10QufcNJzrYE18EyoTvUuEzQs2aUqOBh
29xWJb8a4mJcQkJf2DAWgVIA+bVUldpq7k3050SuDwrViWvJChSGlJTCfMv32K9lHG2yoVdlrx1O
GkEVw3PMQNfFUyI+KsbQ69bbl+OKcI7EvELsbYOHWIBo9M/NZ/YmlEPP5BhccId9QuIItN4BdhKg
W3PYAMwtkNpUulDSc7zlA1hTYN5/aJoKoPMZfFnPHPlKUhJUrBGIUEZwyWll/rZnPZULsn2TtnFP
l4RSpE434RWFUmOGitkGg5QOPQ7hF2sXciwHxB2s4qSgCIyTkVhy0WlV+7XNHqRKI1Oh8dSkYPyY
EfrCjVfM9DgGzByoZXNRAJhBAcoxOYWTJO2midAVEx1cc+C0AC9eiq00VJDBL/UDuoh6oTiBAaex
vyKpIe61ZDyxhmQNyV5rLV1NR94Ec6/vziZeWRmSJghaFsvMfVS5Ff/YpKz3K1u8+vSz5i08H6Uf
NAis5yLKeqXM4xwFZidbi2NwfJ5u8HrH/4jIM189XsBfZk5TixQGZ86+jGdbUpPjNLzPzS29U2Ix
gLLX/e94A9y9ddMhOCU67AE5L+gRIsM84eiLPY1uk5C1YvlP+bLZfvXoV/A738tpcbeiRMc7liY2
2mFqfPDAn4v8Lde/hcFU1Uxoy8Wa5CIK+LQF4vC8PMNRojehA/VgZJygoLxeBmSUo2BhynT06ciH
l8Upno+BvXScyNLMax3CkYUb3kmtC/TxWk3GwI1nurpREQ3BsXclukb693mSne4Tj51YqFb4bVvp
ca35Ud0fhZ3Ys3wEh9jNuSgp4WzrLN/lKx8oArQ7DQs3uPFSzGSL32IBjd3jLep1XDBwY0bQeSuf
qDeU9AfZ3DEkcBXnPa10P5uMbCeeKP+a0C7V735qgByRA5pX2o6lrTnqbMx/RyJ0vNjoSvpHQIMO
MCOQjtmhGZBwuMm5tIDpcgjNM53cnJegzHgwHTFV/xk4uWvoGujfN19cD1alf7FTFpbWCO7gduus
6E6vSu2WD9kCyRyOa8BiLSc9sXV0YHXYkMBGF4kiRZofJiRrbJCMgMnVGM6Ee1Zk2iDELlq/PFy8
ZRc8HSD+gltZEmTPp5TkiwDRvKXSsWB78b9qjNp9c6Tq48oavXLtYcV8czBTI9kwT8+7UcUOQmQy
kYzRGtoKxAI9Ur+yxoBavJUoge7jH4wmyRFZBdUbgnkZ0gnHdMqp2m1sTxRHTZVimBHvp6rGWyoI
4730xfRoOYvWZA5rTw2wNmByqTtRR+jxgpmF23ucRtvt/MM+qZW1wHPXKBaMJxtAF6iC8nmwikRy
0+p55lhW6ia6Ffvzp7tCDasbM5BxIW+4oyJBYRzWq8U6Gc54JOMi+mdm9orrhqip6UwiVE00l5yk
9cX+qknkC+klIKQdS9K6CgBEaMg2weAtinRNIGH9puCSGCLZsYh2wvMqlONqJG+jUeYP4LexGA9S
+RmMWC2JgfvAfcptPOf6XVEhu0IDqduPnWWyYjdXQo4UD7a4bfMGbmApEwGwG6g7C5mBzO+xCyAf
fJ5V1/bzj4CY6KDKZ7PD867Zekn9vyOw+sRhcIBp8ySAqQedSbyCndsVDfeYPCRIVJJTpR+MUtT+
UwifXF3U4lhnJVKNcy9xOW3rwSnfIaLMMAFyxbU+/oOpwiwCmrPFiehR+itEuLQWiVG0C0BhvhId
v9RDT2ViAHdoOSMe3Ts8HetB/ioubWN+UURc3XRhNoLfRcGCyxsf3VraOQM8RxqRJAY7edeuuJ8h
eQJzhePUGo8dHXUo90kbxDG0L3BkbpqVwsOYl2jfJJYMXsfYJkrBGy4IkDX+4Rx5M8KaMQjv3vaA
hO2hWR7IXdoqLmbaLXXkAbB0MUHZxDiak7hnJbLEQXyjpMUrUBTA+CvxCdSKmQmYXIZVEkO/kwau
QfIHmxb3ueVqUtLUKbCr1ZjI9IMk9Dfwf2Q6gyx27fZXnFK7mW5SyH3TMf7nOYYxr6NDFrAhKbY4
9GU0rEEjEsB0HNXrO5UqzCvpE71ojCOIlFosl1b9B3gEk7GjqM385MCSogR5wgS9C9yYf99O66Mb
mjYPJhRCHjqNpmyQuk6WKXJLTjjcaonaRfD7bMPViF9vB0pl9ey5M8FfphOemmIPjmj5jSRgfb4N
hNwLgcLUEoB5k6+Pkn+JB7IKqdMA+yi1D4f48I1LOaweMdiD5t+QA4QZ+0imhDKx2mcl4lnUiybh
B7s17F/8hXo4aECsjAFY8u5m5kIVu4HIwzC9Ub/Fs8FYob6APiOHP6WRpKhe/jzK520gPuKxT+KD
CfqXquQsmE2QdfMuS3sDEhkDvAOuc+UfMPmwgY+t75wkz6N3y/Bpx2cX0nn1zPZdXR0h7U9/+6v0
eM5UcsmopqWdID7mmuEcxTZ4tFkv18kuOguEt1BsR2ZqXFatxD5j7uwoKeunbFOHSRZ/zzquOtv2
3a1f4NJVY3R5X+MAnFalTOzGLVbfD3UeO/7ITorohBPy1Y3HcERUGHBbvyNubW+S9qidtF4p8HDz
I3+nWj8jZrQ/dtYQi5eJQfKGDb99uArn88dVG/EIOE9HbBP41p2vfY7gstWvkJpq0o0r0krSQ263
D5H95Q3c+vG96XjxSiFfEZ6cLoud25Uon56kYLenhTnhnvgdc8JucvmKjTRNYKub9zNJiS5/gBEu
yJYiSrssbXp3qPGMA6gfzkqHyxgJyErLdMZTwDZ2phmpb8YTAQ+3mXSlwGejgJu+IQQlsjVhtWRy
SSpvLS7LhdyCW0lMXBx35OTYPPoyJF5hnPeIXthoLbMsOU9zpnCQ+OaMml2ZPUEU9XVHqx4JqSPa
pPazKSdxMk8lwkm7TVzOBjJp52gfZlLU+dSa6wDwu/jZXwSRLDpPgCYjl7RS3p80PRLGSQN3zkBV
U4sH82/eAz6P7N4GF7ebhOjNHxd52H/XHF1swkjTve/yOaQR9npjy0dd77qKEZ+/hFOQE9s7BH1I
ojOQLfUidTtZ/c7o8+6/oyb4mxz3QE3kzYx3ewabGajl7us1Ot9fNeq2CObdBtdROWq8hTH9andG
TZO+SOMrYn5hvysH7WH37+9J5m4WnMJPQzmenGoRgCJEQl0VLyYVaK7I1WAeMu/hoSCZKu5ln3XW
4YfT00vWot7Wz1Y6S75ON2Wi1q1Avh78fd7jhloK61f2lxNxQluwKlE5nX4TDlmRgCpqIHXS2ojW
DTpQHHLXD0XA4p+ndqJEyPqWk5uGsrJa6mDdyS0hnviZznEwHTbDA4/QIPEwZQYHs06TYWe09own
EBXEenG27/XRnf05DwtCyvjaPxv+b8jytMYfir2Uv4znewMoWugAjPIAs9hy1DtNhzVzaulZgLP/
3bg5/q8BJZOKWsIak1WXTTwwBVdHfPAngQO6NPoeJGw+ZELmXC1yQnujJjywok5WgW+kiQA6mZoC
pUHulh3lKhFFjmDZOIxmE4/8lxbvF9JzdrYJfejvpXIJfqM+l7MJ7lEtE7/cuZuEvkB5UZGwsPXQ
QOhUm6pLfJbtz2Uifh7ZSqcTbdHHDbq3WJSRpBNZRNgsOixFzbeWMIRUZDsGmLbrNVaIoNcXMcmk
/03JF0/RxYICJuJQDZ/4uwW3D4kKz5GoJ+tVMrHUSu/RJ5fF6jCpi0yLP+NQva8kvdo4EFKBEup/
t3y6oxYJ8kFLZxonNKkZ4eATRbg1nZhQy8OFCBmJgrTMXXMCCELuM6C6n3HCdQpD0KAiN5TTSIcX
FctknRSwST+jDO6WB1O29QTBs/JjR8m5Rdnw7PWc2ynqqYor6fEcTAQc+ViYZScNDh6mvsu/Ja3+
IUD3Tanlw6evI76JByrlXrea9F+HndyrRg2FdvAllXh577LecQZPBGRkniHt1qLUgUFSqE7w8Gi5
+3wL8OzPmpRE+fKB/RS9oRtEBmqZrsICtii/E18wl8UORenN5ZW6xASXqxNy2/ir9pp2rFvLw9Vv
sLSsz3edJirVXR1hgeogd8W9c14XCLK40L88B2CAYalaLLlCkn9sj4SRbYc5dijHfwqVRUPwiQJI
JEx1wXJLOnmQ1YRUVwJd7AU+0mTzSBbIpENmVgjNtZ2PmAOZ1X4QBz06YtxgfFdEYPCKRnZiJ3yk
xO1i0yR9qxpUprFfQyZyBuUcc/TKAg54fUePFCjEp0ADx/9jB283G6bXLheUIt/OmNa+Bo7t0Gnv
8JW6JnZjtV3FKIUtSVDT3e+ae9BbHjFnVLNtqIUun964Wdc0b5iVfp8URaRrT4IT9bNuh3X3osM7
lHXkc+gwSgc+ESHGd5VLFPxFFSqKcn5psYKaKeFXliZgUVk5RMXeztVaR7Hmoy4HjutomkUJjr93
lRqR2ww7/kCoGcEInqjPWieG8rQ8uCPHfJLbsJyb2eSdMyd4XK80dFc0ZTwmTMZZHI9WAoJhLH9T
VNbim2Jruz3p1fNyBzuyUGUiDj26lUU6XgjkUjBivd/9nBjbtJGeFB/JDrr6ZoVgp8O+YONGwuX2
VyppBdaPIQDvRfeY6IhGlmfmicT41mVcmmwJ8tYk3cDzLU2fKS4Vh4H9Tx71tJmHYc5wcyjwy/1N
zfeuXkpLIGoKc65KNtUzRqpZ1wbN8xqKUl996dERuktv5B9V3yeTuSAqBO0HvHDFSGFsjiGiwAlh
6LldgE/bI+b+5ZZ3JJG270WKGItcHR8vIdQjbc5K9LiUDwB8mLikydrCzBoXjM7shF+GZarcqlJe
dK/Hz1l2O6GX9uvJS4L/irZED2P+N7V4g2uiD3bnH0ImQGIvpN9Ix79QOKlxt3WUH1sXRIWEChto
d3MD4p8E5cDia5HM1glBgypdmtK2+UfbdG19arXztsfYV/V2fMWXOV7M9nbJHOACG7GZ4EV1OV7r
D0I0/pJ2N1t0HCn7wRE3j8enHXIAv5iiNWmOUEoNm0SKjDFCaLRQHuCCKf/UO0okCNqC2sHusreK
SLBkUdjzARuUQ6x94w4IiGWInRI/8nLqmoZNVHIS73GgMcpSVgJhj7BKZluGo4LjM7dUDPUx0ah/
1NN2c7a2UQPrv+qgojiPF863HJ7+iqh9hoD41mJXHIV94c6X3bnpLY8It6hlKT0NNOvgxFh3IRrT
jiQArQkGgICHU/39/TdOaAKfWRhVeLut0rXzf3NQsBtjhQXJhQr6/YZQdWkctvOukxu+1yJBo27s
8WbEVebG8UzR431oL9JT5RMCttiZhFkA05vCeErnLXrMOrx/7NKfMRm2Gjp0JY/EMv+mH1YaAC56
Z/LIeX1fcdGnBQoPik2tNe/jiuB8+OR391w/GdLs8Fj6IghvFkJLl05NU8rYkTxtk2kRt2v4bKjj
LxRDkiyqoVTGyx8gZo6r3vYpUbOS+xKHOXwvAaOXq9NDver/FER4ItdmXY0XXiBvCORRUdS2yjvB
kwGd7UWtCqUtpe6KJctQyNgdiyn40KRJx8mbREylJOGbXw3eFFwDUKEB6jC5tWvqv0yNw2ggbT69
YJGY4NdmwxUVls8LZ1ENIkcntHZuVFKOKlUO25qARLGiakfoYOluIyDTskC5gC2KcwtzClHlV6I9
JEr0HN2XBK7RY4YiP935LP37+3YNm5pEKpQV3/MP+fCVCTi32VDvmxXCMlbqZDc7y+pCtw4Ba2R+
8HZmxJhLNEl9wfRWOeys+mkuHeIi+GVS1ls5dPIr0yR4Ul0UaZ4TtTygKet6LoBOueGGB68UcyZ9
VMr88g2SOzL9Rsm6cEyIFJz1vyfHa8CP95dyuKssHCH8w6RVtNdYnm6L84Z/V6yQYopNNkXH8vg3
hG/7I3V4Uct58e1cz+agSYApJw950zV0pwzBQWVjnXr3NjMuD40Os48jT3HjQidNMu8mOTWsJjIH
40pC7FXeRVUUjJBVP4JuiVxb8o+NdXOHJEYr8L+LPxQi2iJQvqu5MKsUj1HDrbxCMEZ9dvfid6RK
DG8J3+fXVGv+QHsjSu/qX9DJKUcybxEOiUMCXv0wKoEcBu/QNTW78zBKK8lriE8AsFXcx6rk1p/w
nXEQxE3kKxWtNpKgcEKCpXoOCh7ZZFuewpZ2JKDfN5dnUcJRO3BKZte7tHG8QxfKULIEq5f+vHTr
GPJHuLzu0eFKzjUq3lh0i6b6DppzGcohSoPs8ZfgVMfh1bXRn7sMSOnm89NjkyYd1w4jh/OXOMBF
VE0plDoQUVDGQbUdoQg206usHx2mepqr2//mrRvry0AAIsiosw71H26kAcA2zV6I+uv8lI+cH8o9
esllM88GMnwWWm4+QGSh9SgO8G+XU8e13NEuRO27j5eA+Pul/C8ZqwCbu0UxubHopQD9ChJLkYQq
LSvfSuKCtqFZ7KD7d8RdNtGf4pF3NZdaoUeHs6RpIpwQ7k2GJuwXGcXzQvYaxGrYByZFdQGr8Xzf
E0IMqoO9zndO/rJDq1id/E/pCKlGir8WORmMZgOqs20+oF5Gy2NenH7slpo9XnC10c2BzsjWDEGy
I/iSaY4SVKCByI2bPa3fHhRt+mvDIqn11iHVZvVhBnR2g8Z6U75shMEHasaXy8Kp1laHWJ74Gh84
u/WYO0TnwRsPf0dmBd92IaYc50/YUAbMlWmPVyBkEFG8apzCZLjtGCssY9i5QxXhAMwe0H7T0jLr
Pr14Yi114bg4tg2vCMkSOQDadi4i7AABmwjMDg4I9269/e8ox7DVI/kc5uTREYBdE2neQrxV49Cj
DRC9O2z/jxTK2GuKflNL8dMEpGPb5dUMrmV+pTXohCoub/Ixd78/JbiKHKHxMWq27ebpR/qGh92I
ezMQH6l/tgQBtLp7FnXVpkWog0y8eqweNqIEC1QAsgmaC2j28gkjQBT7L0IeYmlvOHYMUouOmgUF
6HYa2YJy731cJDNIYHf7HUGZC3T+DPuOmlBNLFre//Uw4iKJ81XC7ligSCElF0+dUQLua6y9KeUY
+fMzmN2qF/Aab+3aZvAaaJxtqfXCtJLjrA+FmSQy7GSdRKl3u17RnKCnF782xf9iS7VDdZGjUCYp
uES/mrbJ9UHPav2NSyWrrHShbXKYMvMJuRKLkI8bZWrKOTEXWj4DmSSM0OVVpT/rlEwYq15Uno8G
OMvlhXp8snLEhafJO99QWeNxFlJylWmccUAZoNuVBftxEm1fCUTYxw0ybEHazVfyet1CzOvX1KVc
T+D3em2mY3uVPbkf4iVx5O3rtS6ymLzPi+WUNPAJZq05Qhfrz+wyjPbHrUppL2hwc6+1lueEbQa8
QEmwqEOZ1kmNYnWU43xLMhNFwMhx3TBKRszKIUYLzb4FeLlXM6+kLfx8/NiJLuaTaT5riAlnxw2D
8x84UNyMCrjiwy79j0s7B5HMI2SfLBjDDKMhZ+2KkU+41+GGb0M5aq7sfjTY1WqGqXJhNQ2cnXXn
Sem25fGqfP5GSLSIP55M9fkSehCMTRtrcxC/woiUPWg268lLOGAtIvugKHQqoDLwuKnIbAca376x
XfdzDcC5sRV+4A41Hmp5pmHH4CZQ1udM+zaJrubAuJvri7qYOOF5gfH/oJKe16qi92oanp4ZeAaJ
atIed0FucvunwAzI6fsgOuRliKgOSfUQI4dKCoox3mbOAxtUW4zsEtvfgGDv0rIqOY5DwPd59rZj
f29R4BoHX1Oo4MdVzUhloZYpUws57v4maPWX6Zo2aa/gJSs9AunbZyRahp2nSQTJPxG+JketyIwS
h5vqJvyALUYfuTZlxGb325w81eVKEbzikmYZWbWZEqLOuZa5cYrqOOMD5dSyQC5XqaZuh0bT5fx3
PEUhwgxoz/YubDzvFIISB2UaCt+cL84PShskLdCiwmu/y6R/Y2Gj29KpNunaAqcBuCylSoe/7YiO
Nw5lAk3FlyhGpm5zSTnvjea/E26Tgr4hgEKMQoD8Smk91A3aefuv268quQQZBxs1qj9uQzvZOHfW
4dcp3iOOWU4/AWakNxAKY439rI87MNxoGZIRClqjZr/7r+hjQQjRKHey8YkVTafviU/0Esmi+lrV
ZzjHd1SztJV8o1dEwfbCIoxnuCQPTtgNId9/Oexd0cIyU06XM5hM/4UCKz5T/vfowYwmMQBLJMjJ
xxjIscSrXambxzvVrwwhrAd29x3PYc12pupVpIBwk1ev6PfUd3uJa2p/JSzvih8+XBczdqkSO9yq
BGZZxQJizlkaO0AdDlw1l3OURCSaMAZ0WqQ9QgIq4Au4qlBfNE2vU6V7PIjk2dAL25LGRAM4pk+K
EFKJuAdNYxo5RcmlW5e/NAQs7/Yu1niNE34tjiUVYEvBY3OO8+OZo+P/09xOs+x+9y5N7I8ZPjfC
KW019ieVHd5Zb6GOx5R13HrePx0BaivXx0D83bJ4pnRM+Ln54YlSqS7VCbTu20Q1PVWQVAFJmLcC
+AueG4efHf2eG8M0esbV6hnKw8T2j5zzEQENORJolvG7lZoLdwiq18dv+HiaFNeVz7BW0Fi8kRxJ
nPN/F+h9Z8F7Of24nGgdCbgxjEsXsTwkSR8vRevkeGTbZ3IY2V5lrANWrwKkZr7wCpEkmRopgSb2
JBeVfWlvi06w2S/LqQEgVPHv2dqKcEYiBCIV937JHzm2tSDpW6zCTdW+aywKmLUX3MYkXM2e8uXg
aanG49Hs+09mjdkRTAeMgo1OIr4gx0uHcxlDSW6K98tL72kyDr/A4tFH/73kYr444E5l5Ggs5pF7
x8IRyKPZUNGHmRAfZort9jt3D4FwmUMjVu7Un4i11w5sTtZLs6yVi0rwLBj1mq365ZLQKWai+3lu
ao4Z1UsTUtwFy2uOYDH2ZtahPVkC451BpOld4tVVI5emaHXH8lrQSY5HrRsA2+5Gsd2fp0jOEKVe
LecHxZGU41/CfXwwrtWm3s+GXrP2BXYZURuinkbEV61pEjeOpTfPYSouMzPjI+tQG/1ICLpe2DYr
20K8+MG/ggulsgPODfFdPmzejMxoNIqtWGTFtoOg/Rp/jkfEioBzUFomODvTHeRgu7qDvMlS4sHT
b3mbJIX9t1xmPdrPMpFEDXM4rlUrHDqFuNpfdpjvmUZ0HuiFUnBYUr+FVy72OdG0FRDVtn1nVS/2
peWTi4xPiDBdowPH78W2Zp15xSbvfZH0EPnUu+xmDhgfyKDKaN9PgCc/0Z6+JZ5+nmakYcf8volP
MhqTmN3LnpJwrwRzXv8wamWZRvjGWX84RqPp2ZqkgirHQkf9o2dwb9h+JPtRenEIoceDGRe8X29o
IDLUYNIIfEyw4yxgdNWKBQx2Ic1H5ONPnBi8w6E4HCyFzkotNSbLlgxC2DtEp9evpf/VuPBBNhor
xN4lCm09Y+ZLd+8hhul8wSDfERjfd8ZI8k6PJhKCXcR2LAIT0zCeWnp1L6LJNnmAeF34BXfb+MH4
QGrOLuEumfPRqq8Sm14HO0Ege3KmO3B9Xscisn1VZ0JLZ999C4jIetn3bOxPhPBfHLnRBohSyb8b
jSJ8TViYwKG9/kfV9oZQnAVAa+CtM3qQVTsLPo0huKl9kkS3I5+j2XtsFKexn2YnTXsLXhXXuPil
/rzAVJYzGZJ/vf7AqSBu+NNTY5YnNixksgKgwqqKpDsk7X8/oDbpdEkXutj0P50LBWZJZFzPC5KZ
2gVWvPh98XLRQToLoK0g6KyNMeV9KeCmes2k1MzuCjNwAOutUG5WSTqEY+u6xVb7pamx9ZrgCsWC
ZTbrNWWIE6pmNSbpkaFtofoE7IaGdeEqtOlWcXFcdO73Jc4lJf5g2BP6Mcc1FOGaeCQev/sCrySg
R4jExrEC+nXBS16r3H1bS2/XmlDpzONo18sOQjlXPOabayZ6ngr8y1YsVgrJeAyrmqus6sV6hxGV
alHpAOIxBqooOLY6wwgS8MkBEhhZRZ9HaD0eBxdSHeEiftorr/KyKzfIkEct27xiAC+03KXoC/og
ZNym18MOJ62cTT7+oOwuJ3YeAF0zSXntzcX8WpQVmjAiiao1EoeDDfvnImFuGHJ+RbT9pFQDRva2
yFxn3g+hsFAuH10IjnmW6UVgKFBNIMEh677f5QXzd9nV0wOzMCTda9Wcfsfng/JVN2xhYS9+bxmK
lRhtuRz0X4AprhgcnYGowPbqhhGWUbyqgvxY+CgF7xjMMK8gOfHskRW0B+seG03UJbVfbTgos9Bg
h+h/BqCL0pStNiXtKaLVIMj+jE2hVYWr8JhTy/JSrsAjH/Qzj8GCTLxobcx50ArIk1IXJe5gk+B1
pvFnzS/wQWkDPGLWZXYXKsWM3wifu5RlJXPbOkCs+hallTGJPhp77TyRWcEXG8MJnvmbZTIIfgU/
WXa86pU8UIqho/4hDqAAq7sGVCplLhBx3mdCs0EgiKVjSyxLqN9y64w+/tbbAVZzA8iAIkbIeXdV
gmv9ob9VROQLdALjxXNwAjK5A/llOFnn28ctK3d0dtmupppZC6EkX7EnSdlok6HEOQ88CE6rBMXJ
zCk2YvDmS6HUI4H7XsmnbbuyRhM8jNG+Wo5XXA0w2kml7LFy2IxrvSKSHzt+0MCFDW0UnoT5EMyu
E+hX7kzz3MBwAnqjlOo9HmRCuXS2Q8ewqYg//4GtvX4YrSXodtsnNyheomc7a3V/1yeuT3hv+bMA
6GyxfRtZwmzyYgF9IR8tfmB+Zw9pnby+QA1g6YZS/mnSbMlw8DJ3Qt9LEgNbT9uJx2PcHmib4k3e
H/6B12VtKkBh563iWXOgH1ZMWg4ymT/CT7bCgrt30eCfLxZ+wr1Vc67VzZGjW+IEZwShtjT//AJd
tCojGGG8MUOWYBgdxNvf/5dtRQCOUTQC++1nvWlFbZP/nsP4/cITs4gmJy3Y33+OcrT/BZlEu5aG
c3eVGwHisYTnjlI+6QcMh+cSJnb2MVd7hcJ9ui0oR4siO8XfHVogy3inH/tLdE5nGJdxqV5vqHeE
7zgyuAbOv16eouCG9heQ+BO5voa6CdZ6oHmpUB8224CxjQxHtjGoDOtIOWb7ddZVE0RdG2ah6APb
TzxgJ98oRiOYIUgFrwUIQKDpWXcwj3Uy7XFfpRi0/wRGrap9WefIisbuJsusgilqjzaRosHuzc0I
Umh7Yz65uT20FWqZUUdoMlzQrxDbVc/gdIB7yZuugC2eotUXHG2EJq1iJ02s9/R9wHOCuH6Gqtp4
plBNuUjnECDAFW59U9leMszdbytqkqoLf57c3fe0uYdswqQtd1Foe3QDJdXXVWMU2q9TZ6FB7Emj
5acrpSrAJTBfYYMcKNh8r7fQewxu8AlBp+ON78vear4gc1RFymWcBIW1+dZZ/knZcO0/jQBZkGcs
gThKMeon41BefGkmRs2/KRewEEW73typfmi3qcF/9A9+8eZ6hQkDbpAILIwSN5KCKOkIfJA2CJeB
qiIo4CkH3GpOPKtmZNth+1VWmA4XI1tcAdJDH/Pn9JtK0rjpSAoKIHfAF1U8TFPuVqddMwbBGaMb
rI85J+UjUVkugfep9CRl//kVfZgPPRROboTxyc4zD4xPivEq7SNoK5ilWRwl0+I3mOp4dHs8MLns
1cOYmbb48kwze1YNJZOX7GdOMnO2Yju5ReYV1J4BIfhQurEdiHAWMiIAd+rrM8EziiXwUEO79wOq
AGFVx7Yke8gckTPIA9YkZBrNH/njU7OFui+vxn/LGrCoQjLSmxgboJne6KsL3/D7L5JZaaDjkk32
1/wtBXafQAezcf3mw6vzwbbE2BS0xW4cd6/7406KyX1gFycfhJcjxGdHMaNa1OYUg1jzEXPMvRUi
EaB1BSI7MRY+Z5qVXDFD7y6VPiQUN1Qls4JBgZTl4ApoeoSdLTD52otX1TMt1bCf8HwprRY1XUmJ
WHAf72Nr5keuzpPEkkVYy8Nmoi5xHICoGRLu/PF6Gz2JBE09NKQrJGxVLAW8ouE7s5HClmuHqCie
bjvVe2CqjRJkMYo2Xo3zgkrisIe0KO3TH/tI1byWT/ymnHRaU4/ZL99mwp9Nmf/5uWbOJ44b9eFY
kqLB2DTRGP0ymNe92WzMOA+198fpye2TjasUDZ+OzkiSdH1j8SseFLMeFFeX+UQgDm7tRtSSIwLU
e/O4kf7kirB5QEDd6MscTJZ46yr5ly4HjobVw6keDwn2xWZVQK1qmrtOJrcl7d56EF9BP3crkzZN
6rOGtzvHjXoFDGxIXpu8qcqt94kX3C3KQ9FGipdkFDuMUgPH5AyYU5vbCcSgcWE0xAlv+my67XqV
9HT0DhlXS8skh42D8tLeAo0iXdvwvG9JEg9CmRinW6hnW8AqtD04SDly7SYgQ9dJ4yUNzF7qa/sO
3p1mxS6VjdUxoW4XxJPADRW3RZasVhE9MVZpTovicN0xs7o2TD4Inw2CkCSvIPgvwF/3eFeGaAfo
abaX1G30ht4947JT4SDcKB5eBAVuOUUfye4QKbARek0yiOfhUh3xbzO8t0Fi1/Gzf4aPRvoP19N3
gGS5fcmARhbSOibDVGSKvCMYVGV61DQJzBRaI4kxaLgFlHde6Uafa7gh/cCZm5lIFf3QQmVVxGKP
Ju6Fxwt4zJske/0hxzFh65SfxVA0ESD5XDTLTPnuMdydOduApOdOsEHVsxlKIWR7Dxqy1ImDLl2M
UsPRTFDlVauec3xELRsmb9HTfhaeZHZnZd4gSg8DrmPcqz51zTGCsl2aahHapYq7SfPpint5chrR
texC3RCTXbgFlRHePkviNfG3BEPlhuegXjSQiO7t9tmPtyWx3Dx91ijjtTJXF79Pd2aa1BD70WuC
DD+hC7az1yavn+9v+Y/K+7S91G/3M+hZv0vVI94XYiwyIqRVGrNTx7uICEQjYIz2kPeZs8n6hpH5
JWUABQN4wFkd8l8wYwG2/TkkBVpzq9nLxCDkgEuMKWEVUi4sLv1Wxo31RvjaF0niIN/7aEdIxlw/
QVKjOqxk8sP+htFuVt06q2jJ7qDLlTA8dWmH3SJTeBHxQw96UyID2hSj2/yAKC7H2mdV34q6rQgy
1ffMQQDDHWgtB4NG60rOYJt/5nGAjrmR9FwxmYmPv6kglcPMZAnE0yRJGT2A3QPlQH4zz9Citt7Q
N0MDf49+yVa1pJT6usk3qFGkxRmxLXYuR/VEU74BeSa0ELHCAXs5s0tz9cIBcNso+eisWmjvdIcr
VyZ0EIgAYtbbYNViV+dGw68oybzDcGQa538rvx2REK9oBazJ78xbbvZ1laJlFdKLqSHJwNrnRrU9
6yPJMqhMLPnfZyyMYIP5NSDdPzHHnqZshe4jCHeteCV8DY6YH9A3TPw/OWv1LJWJ/VfJbyMBRzPJ
sSztFYCwLHacZDb9P0pavIQ3Lf0vx2kIoeHUTVmX2if5B5CXbbYVEig8/oWgJQI1dyvKk7ojZcoh
Vtx5srOrAdo5grgHQLG2LTIMg2hMruNxqVv4Mn8/buZr1i5BslEWRYHzC8YxVDHZS6bs0SJ9Sy8H
2jAYV/yVA2yJ/unqRA4Y9Tr3F9r5P6DYc6nJxtZzZ8UQawBbuomi+YR0/CHLj39ewXtM2wkoj/CA
Zk36wGSJ4JocaFRM1yxoyafED6xWA/JWMo+ZnhMINR27A6EOS56R4Twl
`pragma protect end_protected
