`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10176)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5Aw0DkeWO3TFNRVsnQu50ECCcSDdTLIjGaDjWcFUDTGUEQPHW6DtE4Y4
z2mQ9TW8FM5GEQ3zYCZ+vC5ThoTEFPsiY+7cOgQ9jIarB0mt5w70Tvg/UIzR4QJXXhM4KILMYd5b
prnNwnsM7vPQZ/FLRqdPMNttpRm6kJE+NdeqkTZyVh/0a8SRxf1HVEqp31LjoBVmEWBbCtEj0XJ4
K0Vm/BJKTOZ5GsgVmooxWdbh9Qz1Uplt4VVJ0pfxAAPOQIiPChOrciS1601R0IYvpwCowS/ixXTz
qJVxOwGNQIemSB8QBV2y9DQ+rPVKsKZkqyRO79aSlfQo2LwIf8QN44nV2W7fDIp1WsSxdlDAf2rw
zXne8tzmRqcak66WIAW1s/ZKw8t8AuaIli/sht/TIJQQIRMftVrgAdFAtKMqd9pxRF5x5fj8l0JH
QsxKjy7aRY96+Ulot5IwyrMrWBmgK9GuhhoXujAEh4SiQ7Ae8mszNDqjxIIA3Q9Q8nj6wu+U62Io
9NtZop6zjtWkvfr47CZ4MOcUP2E6MsDt4Gii8055CuTbQZcVqrFAwsF6Ygqc1Oks/Veizc9a4hay
90Ky9dW85kTNyVStoyFReRVp6zB76Gw1Xxh1FTQqIbj+IzDzwbijsvEXH/5CwrkpFoGBHhNWXi6i
MWQNz31ydj7iKYYpkh0NRJEItaPrX72Sc9WyVP1wIwdOhxM6AJmPggk0LlKJOfvNPmdS7UVTXvOL
BcoP9GJmF6+FzSJPfORz4TSHDew4jCO+f8UiCAmDwJPcpdtY1sQ+1Ryb2YE1T/WUw0IK7AjYjaD4
PdzLL1OmjffkyK35Z9wrFCbVFcZfqzBrRPiVjr7U/GePA5mR72cKwe+OZwDOhlGy5N9K2VRs2bIe
zzTfbuAugfaK9BXIXLpHcXV7Yr75kdcCCw7M721PGXbGZ3rzhI37xrFvp9fYvrf1ILl9/EraYjFw
0IXtiZs+1sotI11wgohm8zJf40YI2BPffIVhPfU4pd5sQpvwbuyZo+E7HLVi8WqzBR3zNvdWAPR1
aM5O41GwquJQiDAv229Z0HcVi86rgZ8YpQq2lrCFLD7jbDDkTih0K4XgCx+d0bsASSIurkVI2W6V
GJWW2TNSavlAGWX/aNs4W4/n+WpxzUlGu06Ud6VG6j6Xsj5N/WZZmVsxdybfc1CkFaMoVA0URjR3
XRk79kzdeeOggL6YoKvkxQ1FrNRlPC2HImoO+7BztGTfid2Ogb6iWngx2bIb4alRJwtqQhgVOmMl
Zn/ZPCkdyP6BI4dd6BOF1Adv/tXRntumMrJwC0qq+SPe9wzEf5mSYYtWSrMtS+125KFiaIJMIZdO
qJOxftcVr4Hlh9XLBgs1RspxxlNJAOefosBOzGEbkOdfmDHps2R2BB7WQ+KLtLzomz0ILzLymAcm
3cmJQoeo/sXp+oebgyb/fv00n6diW8wDC5yOdcAwfniNBL8Osz8LE0Leg4Del4eCUnXHgYkdEK2o
dS6ZyqIpE/FcK722fvqx3nsvMX3Vh2Q9pbbzZWLzjsQNQ6gYeC9GFy0mATNrAYhDk8HsTn/MkXD5
qYSXP6XKC5dSStWizaH4Gt28EugfbFF4DHkztq8FSiwAowiuZNskOqhbPRcbpZcs0pZ9N2ngbimn
II9bwkcCpfMTHeGDpnT5/Wj78BhaULypQIQwQwz8uigqOPCqauiGX8+J2L9Sfv4DViVwTLieiDBb
udO4OGDaHWM5y+0a+QvYQ2KWj9YeHcd+6oBMN2hHtICzcWUSp2TKxeq1jt7PEQkf2LGTFM8vpiYL
Mw7hEgIotFp70f3NuJBuPQUfZBCb4TJg8eFRNMOIWLtMabxHH/cJRuwQEczls2FuuP2gHj5C3LcJ
ohED3NQkDNSRPDD3F0zNQkcPAIUgUHMqjpA7kf8UwDpcVWEDA3aV9LzDuVaEF82lV/bzqZ5NMBPc
+9bZq+V1YHSP40fXXXZU3HT7+ybHnG5Qnz3FFRjiuy977HjEHmlnkuRYVtRxihtpZ218uIRSeVb7
Z3JRip8eKFGAIqwH79gQVga1bPMm2UQzGlWz/2cYjBCZdN86sa244Zl30WKcIYAD6D9hxHHvg9DA
sY1lr/TKqVXWhRPnPUhHiUH9U5uoOENVs4Bf6kYEr8xyQ8eiR37/iiAnOtmkOlW6KFVet8K6lwfN
Oq8guhAz3T83m9gXetMWT/p7OgMhNT+l62JmH0xGqy7ShDHJRLUH1xVeST9vrXj42RnVWRQOIZ14
PAIfni+AE9N44T84WZW72gM3E3mvelZEMBW5rSwjcQ3tzXRanjPU5M06qGL2BLmRtb/q5gtr9rVy
eOXjNZcXuOeROz1UEApuPXOCKn7bs2DGbgNL7PnJOp3DAaffzohgUkWmX1f4Dme4CF+GcERj6pnG
9uOloVwPLyW9e2U28u1BcWvh3mXxFM48YPH8SmSRW5SVgdipsL/Q2Zwcfkkrv4j+ADprJBagdOkR
bAersrqtkSyHaamfoVQOrg+ubpjEbFDpRjm9wlsDuXYZ+i+keMps67knsW+W+QjqoLA6YadlHIhn
tIoaLTPHkJhMvjdeVyMEUJxmcyIdGhP03lgjd5a5Boxw0Uv//GpCbRxPil5ptkVsxVPgWMwJJpy/
mw/OxvCTFgPMSP7yRymMsfNryl1L4ZY4XQXD2VEDakQgxsj2nD5yT5cvr6NPEGYjH3qFOIYmSnz2
tDAd7eqxbdgqH4uYWWKEUUBa4gwUPsiJKQaVIkK2nf1TTtqEIroMliFzUCMYZ54+IQR4Q4UQITf6
ssIz/tuG3l0iHJFnOZHA1KMsSCHYj8dyZ0sj6p99of8K1M98SVMTNyrm5sXAkSnVyQX7A0A8yOnS
wIyPDJBmCVeQpP7oPpAWX+I7pUaXO/42IBeFKlyOYh2oSZKMWvMeJ+1QMPJRtVNpilhXBwgPDfOr
nenoDpSdafivoh+dPG6uDXcpaITZz3Rj8qHvf6mU4/Wea+t9wOmNoV+y+so8dhJTngFioy3YuT73
9O1B4T55hBdepBFwvPdC8Vanm+ApfZNrGEccsJQXfJVzK3wQ//NP2nSTkI/80yL5lz6q91YDFtgm
sUXOFRw3z7dqKTc5wwhqWcPotSLh+Ae83fs1eH8pLCG8Ohy5jJWA96Y2iofWThYW++4cknfpeMEJ
U+jfDsSS0tYYl0T9mRZ/4hsAQL0mN4rxjrffirNn63CJSOgFOO0TYji2wYmRydulXSyjROIWlx4z
AbIfuTDXdBbXMtUnX36dYhG8pzaEcmetnvBVo8FdU4C3tI2GmKXTqqJSTNn4URRMOYa5AZnHO0ep
7WY+kbKbCyZrVhybk84G+SC9ArmGoeRQS+Zy6FYO+Qwrx6QAi8RgUGWlzJUiavPIWpMef8mPIpaI
tlion3LrPJ9byMBPxxqfsj5M5BrmE4QwYW+tS1CfPzxgfez9JXTPHFmxFoRNDn5+jM+0AugkfcA3
hv6M4jCzdKC+IZpgDf6bUf3nb0AUVjy+iJf1u/rrSmcC4tbZcshHyDhMe2/vFOKextwq3JadrvpQ
wjrNOW3zCtiE1xWTxOOXvQ3cDRTqYs5cdjjfLnZC+nnDL8SLqTN7NClvcPZ/coflG04Fw84IMra6
RFbE4E22YO5yYQP9/NsEKbue7DSWkfN1CQEWcPAK+zZcIfWh3ufku/PBIjEmKh741Cn+cK1mZOxj
xph6xHPFFmIMefhXWcEC4pXh5ZyI5n/f4UERZfTGQQWQIGqVBnfSchJG1yvrN1MpZhgIwGuHz9sI
wO6kwLeiIsUkSFgUbURfX69gfWX0N5pYqZitER0DxudPGRxaOVYaDN93IoVnTtJMF7Csp+96eu5+
W1WhJEmwD0BUZWMEpDGV+wnHf3ZR7bH6B8nCkgdoMg6WNlYgkTvO6txi/IT/S+spTGXk8QyQfmqo
/kusbCqfAqk6G8ZEb1YZH4peuUEo2jek3JlXBwt8Kw4FK87tVNK3HmFk+nmsUVf/F6+mrX7lExky
U96G3gwTh+VCfbyF6YkS/Frjo6Zg4O3IdFsUnPUgzP8dHqXf8Z20LmpRQ9LYnOzmbogHYkh42/wq
xZu85vcfpLO9diOMmg0p/SfJZW43c88tZbLZEB+DDfwz3bVBGNpPNx8bKoH9AkjcONu7a3GL//Tg
j3S5PgV/gdfcQtx9XNj0KBefSwiqnBSoraqKoHq9M7me8fvC78jGOqcOh69cGtGaJ5+YL8SXO35J
4vgW+WwIvl9GUe9T6t2rirsm+Ic8K4JpySg+LHM5E2RV2NANTg87UVJ6wwgplJ6Ysxtu7xEEcEOf
xBN5yUjLIBcHu1zzMNFRYqvI0sKkNPsTkyrTLd8+7ribq5PW+6hXaCMhtoraQvWgmi7LIiagNtv1
Vc/53CzFwA0Imktdk70spbAeA64Q7kubHzH1dLK73UUq1St2l5Tkh9UYEoK04MqSW0DL1qW3FCzc
S3g1dBsCAiBgsavh3HjOwNYMTvYy/z4qRM8GcCGNFa5t7zwJI2Mai2DpTgrIyj9/wBBVZZTWNUvQ
HeiRcRSVXA/M4xdx61NBQnNO7EaXFcOKphe1Iv6SgBop7QZEDT2pdp2R4JVNN/d7r7/dp+BohNse
cqcJkMozbpOXhh1Ph+gWkDbhDwNl0kFWpGqGhqdYBz+vjUQHboGPsAWMIVr0vMbLVhaXdtBZTHs4
oSgurHaU+3mtjvT9xl1oAgx4IOZ+FVQQAQtfdxwv0RDri2SDpM79FymitpQtU8xa32DMZxvCxbbw
Gn9ueqhy0BHmgxOpA8U+kl2e78sXBH9l0dkAKOyUSlYgeCk+0nQls7domIrGCRcsbsZFdry3Mjap
vEvnaHrQdp+491Y6o6EHTj1paNbJTGg41KVHpmYSTuP40dsaY0QK+Yob6U1ZEMZvIQD9pEM1kFUH
5gTnO5OFIDz1OyVXdqEP9bKuIzJpXwYu/0FgTFdAvvwS8QrQ6zGYeB4ycfE0PjmD8EKMJ+wjruWQ
2StP6TykG7wjK6gd05xH5LOkJf9gZR4LjDaNVql05UOdWHuNO3qHsszM4s0hK/33EBGtw5UJiYM8
rlKKsiPeBE23X7rCXuhV3xlV+meon13g4Fli205Fy8Ofq4NIExaa9/ikwzvcDk3XSSdyedYKZZvE
/pawwGIG8Y5DYsF76loVs68/K3Sk4b6E/V4QdthP1q5qw0tqDeyej69Xsj5onAV5XitBdyn+55d6
wlYXz5uir8QdE1rGpzjSNUn/SLhfhhRU8+d1xndYtH33tHwvDqBfouaaNk873zRI+qd51vZNNly3
A2z0tvEMV9drAe0IfcRSXNJss9/CYmmZgkipxU/spybS/hsx4qK4++hkSWjIbzFFvDrA9XE2Ilvx
uUrv76uKAsyQBS7VUKQilfmP5r5eDRFTV4UONwqzCHmSUP9Fmh1An55mdTEToF2oSUqSDp4RoaRV
uvxx8wzo94zwqlLVZyjXlbDBNruWIH3JlZDx/PRcsbhguRxLTNtc9P1+2UsmfTj16YY8GGCZ7dnM
ttXMW14HOULU9+UFKoi5BQ68Ynz+Q6Ql5dCtFKrPvO6Lb2F8V7S0v39b8/57/Ha7L+EZx/AI0B2G
V9X9D0wAJxFfptatbIGNg+RqACqHwu8fJfWl9qJO62HWNpdllMOdR61zBCwjtO/iCs2wcOe+Ni03
bXsc/w9hLrj+9PWbPYyOPqPm0WsBjXHXWfwWqdA9s2xipSbK357xqC0L3nohS1MoeROj8D0KFGBq
FFLPD/VJ+YqUDwPx8lP5rrBLmb/9VSYNa7rcgzMG3EqrSrvItBZmqbSqHc3Ie3qrHbyk6D4CBRKF
43yuO/bRJolQP3WUJzR7MkjUg0wb+5wOkFLklyPPqEXURcPeyVHSsm4MXthpStIdHgthU4OCQplD
/BKGDmXLVcxsM4jT641L3QPy3F+iL02PCwEF5tUhjEo09+KLR45OYzbiEh5Y7WwuQSFExswttWph
1LRfH5I3sDStVzVoqHb4c0L8HNVr2N6ObiHFrWlKD0aFU7W6X3Z5qzNAqaFpOZu0seW49zfHRnxT
rXmWFLh9grO+GeGIxn/N0TdV4VrXsj6ipIMGs0sAnsJy62NjoooENtgfZ9xyMfAWjuiuY/YkXFtE
zZuKCuFNVlM3tVCkGKIhMBqR1Myr8LNdVtiFiHexIpaB6xGVTFMd471fm1/wMSwCnLT/MQz8xUq6
CiZ7W3JOsZxmBt21LWIeDzzsUPNvwkzqJjKc+e0VmjhHO5+1CW4ShLHSto0g+zYxj0O9BiZLmyFB
H87CB8nuhdnoRUT6KyHL1uVVpOxxuXF2BR7o/3qG9G7Zb1kQBaEmEd8RvC+0aJSdkEz3bMyMD6TC
diQqw56L3n5ltt5DQ5WyVeKIQqmhkKgr43I/J8Fp/3JwLEpJXgPLJimL2VKGB0cFgPcEXky/0n8T
UcPS2DJCysXxJvYstbBt5Qn35+doPFZNl9WH2An22KEs/8QtyHg+oNT+Yhyxol7jKkvBmJcn4rVT
isJTSXQfeoJERRx2wz+wXEXVoALoxIh7P5jXH9a9x6wn3AhcyWbbFfyo6K4kUhk+zOGeIngM/9o7
B6igszNZdL1NybRJeiBmFicFm2bt1D0NVBZCZPcK2mDPRk50IDdhMNSpn6H/8yWlzCnsgpaDawLF
EL6g5GRtSPthx5e50SEwPxQWpOCrzDEkyUQD7SSQLQRYA9+g3C0hurPvU8oHgNUembbYKUl7sngK
MaUEaIOwhUI/GVPlIDJS7Ze+BPNXOG/1KFQ2tQYqaHyZ+PY67QooLnyGB5agSNFl0r1gnk+gXYMu
JAdQIAaTdn4FhEX3I2bZWTCRi/bd8aiwlpKhlZZMx4uLDl3c+6igRqZpeI24xG9EkgQ7ERwK2zSZ
fy9FalflmjpzJyV+PjqGXl7+crz6/FloQ+GMwsoeCCMnw4B8un+aAMvWOL0KFXERvuJTCw4a+4PA
DyTB+7MoKvY9MzVJ5l90/fn3ExfxjITixiRk4Zmyqcl+UicGOIwi0FnTYdWYvW8FccTOxCEMJwaS
krBTCf0YxH4pZffLZJwlyRpp7ttpDgksXAyIHqyV+pXgb31Ts35g6oRBxyLCcEbqh/B0ZT0483ri
gX1dzbFNby2AOn5+hIiJAnJFC2Nko87VQAOgdqjEn8tFlNW2Wk2lvdXNIiJ/d18FxkFiFkIvUV1+
Nhe7woTyIU+hI1h41fbFyHFZdLQ24+rbfXz/ObX45BEeeiH3f0rJyb4R1Bgkkf8TqrD/lyh2XmaV
iygumrxn0Xl++0rEt7gk8nQjJe0OwrxiqGPPLTexc/646qeILWyxmCjJoItk5RedHzdR4JG8iHI5
2pktKw3mikUaRVc+7C3rGt0bicCnv68XP6ryNf1UwhIyr2LJhbJn4Hm2a6iUK+ks5wnp0NbRx4mb
B+sBXXAaTJ68ALBiJv4ohyKbxnLsenITLweyvbKYoUaUMadyUPwDaaOTUWNE0cFZ7x6EQ02DE7eC
Sa5tMnRjOTLIOfdx/2YK2HxxLCVoECaXTeXNGdDRZErUIzp/cUxVx10L9afv75WuayJYBQe8kLtB
iKpl4OJXJMlCIEjR1k3p6/Q/2QoeJifyXsynV2LTNAVMgF2QZlxCLNubIK5NMGQL1CJ8jJd0+iap
UEz1udxApgNXOWVBqmq1CtRB7kzYsG1afMkOyfWHnrRtgomMatPc3kJ+dzdmlwzWh3oucaEpmp1w
x0NIPo4W+pH3HaQVTYezPy7oWUG1TQQSYRH9fQXntKtU0TtHgiZRJrfvRICsnMN+/iw2119XNwTh
9VFLVKvRcNJOeSYAj/iomNZbMOSzDwCvjkEsjYM4CINgV80/yKcRH/1FZjMKPbv1RHZd0+Y0eQtn
npqszPqf2uynV95b3L8wITzuf+peeYI2XL2+teXClQ0q3wq0XxLzKNy6WOFK/elYZSiCCzEl/xkX
FW936ZIjQB6sncLJsT46q0A+5WbhHMXAyCinfdLBgke0WKNn+elceEm0YdUZLaAMozOfX3ln5M1C
HbklWpGm1qK5ZLpF6DSFNWNd4E2MHBLlT7zYhMTdoxtJvWV0fNMRQYiC4o5MjWSHLj0RQJCSLDhy
I/C78uDN6h7a79Si4voxxqyvopyBk+Jrzdc+18F1xYYanZUyneNOthSoOiz3uqqIfnDHFATfVMhk
6Hs+ciWxmtagDaxBNaUp3H5VVePerx5zJ6S/QMdDyoIcTHmBMxH6RNXKk/4O2pOEE762hMxJoZWN
pUJiewuHnb09d79YEGGHkExNPShU1ZfLH6Wn6bkYSNpx9mSC3rWpdbHbCURgS2HPCeLxVuzAyn7E
xFMhraRW2edElalTXMqyQOfOfikVK7J+L5w7g5rijAla6PGfEvFVGuBZYaWgX1lXcF3Mna7558T6
P20hl90OHoLtux+y4eOOgykdYCbkyqKPVQCNaNl2emAUCE35F/yt2nY8isH7NIOA2UtM0lG2pQ++
yTQFPAlRvYYhqddt4d0E13uZ8sD3tgkqIiSGLpC8QG/n05OwNy3UTZrdwvgTwUwCZJ2TTVrBMazl
tXhkHWYfWuhi47kjBcxqfKke3FY3i2/DdsIjmC7pSL/oldo2WcH+bTva+p2WLe42nubxC0C3PxZP
KtomASg383IXa5CPMtuW3KNEP50zngQgvLpPQJtZOa6mgBlhB9GRznnURitTtWtbgnYnDR+Dmwo5
s+jDIke1Vt3SgFycAEtofvSnmk0adwQRWyGHiCkctJgufJ+xxBB7mm4t5ZhWV3hxsYvrFnY2w6zS
i2VbYiGeTpjC52sN85XTBrW2wPPXFak8tsgJShYKwPyCUT3HoJpCaHwPy6Xpt/GzwuGYZuu9ZglN
j5iVqoBHvtofNio5Fz7tQ2vUafyYWg9zU+sJlhN53tmSd5D/DeiXLLi+JD0KVhcG+MTMVu3yt8tl
+OKoavXiQB5kd/j540fWnBBzDsa96xlAt8qlNOIkALo0bblhXyX5MZLKQxLy/THUsyCWInfJ0xCy
f8XCCD0KbNzIR8EevO/tknh5PHEBDSdx+17hoe1B0w9j9WUjLyIBG/zNq6JykqU8ODKHN0irYupw
c3Sb7zzFs9TzAHUZsiNxwdfGqWHmCQBHzurmCpilqy06ZsAkwSpNwzwY6P10lYJj6ADGdyXoqus8
HlloDWHr4JNvjhO7DjmmhRhK+5gq4k4THlmNsDo3M0VH77AMgNKDhkNQ7KwL8CjY7Yf0wYnQ5oQI
UMNYmwOp6t7/CUyOQaAfpOAjAFwu4a1ZEDSbB872MvW8cmbNb2qhZgL778AXavHUa98BVFVGezip
udBXllOfiDGVCoW92L26xEAU3BDlw06umjfzFImV7FxlhT0YZJC4gMABMxQCgdtXD85nUW2JtGqh
QfoRC7bXeIcq/7NMGh99HiBFMYt/e4Gz4tF91OaItBmmtaoWAYvJ8rZMNnRbAXzSexTAEinnrI5G
jCxpRqd0c6Ig8PVe4i+Hb0KVC0ZMSq+svMwu4jLrtFFMil6bgbNuwedz+RFP9sCpIOFV43lgihRB
MtgAnPOQpMjbmktm3N5+g74fXBz+taABhrVB0Ehw/vcFHFxDGysiFgoskN3cL0l6FrG4jQ69L1Re
fQhSmccaQ8W4DKwuXPcMNx67sJJNQuYUDmNZDqSDVIwXbRbwgpRgLfigEcx55hKadQgM349EtKKw
r43PrwjHu9DNGe6Vukcr8fbiTLt3Sy/2idV07s0XUsKMXkvC1rLSN0uRVWU7tHjiGRJbPHK+ExVm
GRMnbVPUC46utHGrGyIE1HCMU0SzLKVmX3WSXYGizVUmul+rVVMdSHSS7oMP9WphvCsWNA8PXfvF
1I5+xft+kgDJ7na+bqq0GB1D0f1+yg4QI0pp8UkKJ3F5YmMxWCim1AKjlrMKbhFG6wctRDFAnP0F
D/t3twDJBjiEWCsr9konxF42ALYzVXVJoCCqb3A7aMrmu0DI926/bXqcZnYzXooZpGkd8sv3o0xo
RfWHAYaFIlQhEXwyl2PqhbMgqecD52JakDo8aKC6JRACXzAQZazSc9o2bwy9QI9e4leWqyKbco90
Jcoe36MydygGzlE+KBPCUOd6J0xPplJmj/5GmO3pF+svJ+aAAG0gog76P7odfU0P8lim8sQYiPoM
ZHrdaJ6TM1eRq8JbU7FZW8GIRb4olq78iEbTCCI1kl/eLGU0RVh8UUONBWsfZ/jxJg4pYAlqCv5x
/x5JNmEvUs7gkxNl0rhjRSMXvYXcNZd8cDxTXWQjnoaSlzCYArAltNhGxOc0sRdbQjZn+hdC5wBh
W2GC29ushrpj5N9rhPGposLxNV2zt9Fy8XdrFsyqs/qBVS3iZM0AJGgVn+64B08XEKYn4QkdmjDt
z0uL2XGQvPngABuZvGWq9Ay2DJeXdk9FbX/ajY2i1AQdpEhlxswnUXSWwF8NkY24YBxUGlQWsHy4
5SDoAzOYkgScwUnLhqUVEecV3Mpo6Zi3/oJuqpEi+RgpCgZkRRaIlW2NdX+vB9x+ih3918HRI/Lj
WeJacUtAIurjwidIoeOF0CctopSg5ZhsIQ8rYjkA/OjNObq/tNbWQ2r8nEugfWavKrGo/eJh2VVH
VJhcm7flWkR/YtBUZH5QjBphgklnsEdzLOsdItXT0dOLMZmZh3c8mi/jsnU7hlkweT3ZW6q0sIDd
ykUpfJSHf2agBEV5LatFnsEyZkF0rs2pY9TbufSkKsdgIrXKK8Sd84E9oxUxX0Fz/v4OQ+Lgsane
LSpvB1x1mhG+dQj7wAWzsCNoIS3j2uMwKEbsMY1exGQIH/BGuE3p8qI4fQkIG9r4NgDqzE6lErXz
2tm3hubafZ9vGwVRpIm4bbRuelT/zlrQfdemUvqXycdGCXnvsDdmaBj/U5QwbRT7YshfqTCmYBra
fvIWG2FbBzy+HnmE9i5aXM4tzsFLow0e5nq3JukuC5IyQ5KvshlhYNyMaMoFnjkPcePIuU0Kl1sj
jDtGg8DtL0ul5RmAnkxYFrJue8bC/CN6/HCzco/uB6Tqt+gpWEj2hNKD9kbLEkpTVjL4GFNqn15n
1ZTsTArA168vkmv0AA/VqMt5H4sE2MAZnw3xCzz3gQ7YlUy77q4EBAhf07b2jESkI929YA9Z5Bac
yp5HsHrLUH5BvPPwqtqQvRECMkJyJhqLFaoexhFECque30YKlBlMvO00oWbJGIFbFBaPApplR0Jn
tOWSZJbQnjg2zhvx0WGUMg5rWl9lHDA94T0XouYwUOHSvij23gaziFwODwQdEBCUigVHlT8rwjyM
+IDIZ4H4idf5qrgJ1v8e4UZG1P+MHEFdtBVRBHUejhwkjf0ePAvuDzU5YQyCBu6w3Mn7dIus4b8u
kwDtiof9oleoIGs3jX1SvXLLYnNRwbFdZWEwTmF2p8mXX8RUX7O6O2o+oQO34gycXYkDdsPR+0H0
Ii0fokE1ROOa53p1FgbiyMaD3LKwuyNXmciUei1v4Ln39PvFHcTAHdw1PF9TUUUMkuaN90SGzy9T
xdLaF2hqndBfwwqUedsOxdPuF+LLoImCz174HPE65zY88ipBDeDMODOWugHcyKlXjIb2U+QKcyri
D57c0RQa8DnoSi+gpWZYT9cwlssfearzzGVPj9Mgw10d7oaJEFBT0wHlYA8aAuuI9d9GeYJA8zaO
Pb24EWmTugufEEN0ExqQTl/YNf6f9CUrp6tpexiC1WyAia76d0cnZQ/vV4wdNJP5MW/xGLA5+Vdo
eL1CXI3nAG4mAGRaE/N40MAU3u60ouDaM9D9mqW98AxcwfBmLmoN/tuYd3MStI7xKNLS9vUWnWZO
MhY7RiwuYnClqP9nVZAKz5U2C7kw9T+EomwiWOD3NwMyG3f7O0iOITyvKRytklfjhd6Z0y+koOmz
uZcwn58ig3jHO28ZNvIrpwW8Bwr9DMgbgEw9NIICS+9zifk07fSTMak//MoGNNWmMA/O2L+zkZZN
AlutYFAO2l6K6YYkK0T2VaMirG5cRYrWRrhXMg3c2LwN7ioMbkzViLdfC1Id4LGZ59BmjAHZvSaU
ow89PX6Pc79JJ9zCE43tB2DVKmirevvh/u9CF3o563j2aQbFA/vis17kJPpF/LdGpCV7fEag3kge
U30w42LeTilgPyvokLl82BZ3757Pbt+Xyw2N3utZ287IRxpU8KyhbDbxMkjz7/kcA82QThadjKVr
sarbfOQMxBjjFLYrb+pfp9c3r3cDyqereUpTl/N9tGfUsKBC3oKK5LbPbC+zCeSKSQwArjVuTy7a
dCuWiaWMfG73s3q3oCKKb+qyictovq6rYuuhaXLQapMh1XDicbm9KQaNDH4ASTSuiJkcBxA9vIhF
zdh8OhqsertwZyRs4Q6IuY5OBaBWknyqpgzyYTTVAyNHzFVIsOZEb6P0sG8EerlJoPVOY+CeliRW
0wGvVEJfVGm7KSkAQ40xuPCVM5lcc/uvi4aXQsjIkfmMmCKmG4FK2bhkmIMMRHh7MbAwlC5GCLCS
K5gCLPR+1LYw74cTbc4jXroAH7qysQrDkeVJ5I4W5tVe44jOrCrhLE4IHeCj5nXZVcW8r9zhpEOT
1bBWtcJPI/3aTG3ZoQQ0GkjfNsbVXH9HIqGxXd5h0QtNXi7cWflWipBBp8cb7GK1wdae36fg4mvI
v5Bh1CED6llUV9PKQw257MHLbbfaPzqJRLKXh5QThn4hERFVQsI4VZmuzYXsFkkZSeH/czaSXCTS
rSQOuQF4++1I7w7dl5nOvx1X7DG8CrS8+mU0r/iLErHr7aRX3Fq56jdGHU5BL/wgnOT3Mp3Zl+UP
zl6904H9/GL9iRFoVOhDuq1cvGmh8JOq4+xpSsup2Dl3fu81nILeDuQxcVNVJZiaUVtRdlKpntE+
YKiTLdZlWsi0PpPI9kAysLvkSBUdfZMweruEa0gaxKom/oCJnhHLGvHwAWu5/FYUnhfxWs0fceKq
4uBwK7rulXUOCqX6SUbvUbEwiMM9sMJLvA7l+KfLRlvJ7C62YyIS/TwwFArvgPzL4lLUcV7Gd1Qd
21Q3ZTepCnpEH38gAXJ04S1mfWeYnbSfBzNWgfXWt+4CSAqen53kLjQuL315YWMHoN7kmZn0S8Ie
jReUFj0FOsfUVrND2vYQfESlgRty7Z+JhZFu4zJph2vzPzdenzngCKpdrSuX3WKWFEeT4ytfTC7L
g9LjVvySNJ2ORk7VO1ZdiuJTuHzcr6c+pBEu1DGLY9xyDMDAR+zbs5eRwzv/VAL1LQch90sVZIt5
JnEqTOUNPiDsHSMSLAamR24iSgjdD1ivnvXSA+BgCfgroFwKAwclitGgmb1ggLttIVSs6/gSWL3V
KkOxzMG7CfghrOiKcOoPWS/bGjccBJSRgHQXunKx3YpbuKrZ07UZvhWV4lS6xSgczXawdnn3RceT
L2UqyvmM/2g5Z915flKJ94Vv0O0Bb1Y7L3WfBm1YOENtHPR31a/MXLxt62FgpAnkxEsw1iO+gyuN
bT4jJvlRMNGLabMrMXAq7rSyRNZi56JC3HSNo21o
`pragma protect end_protected
