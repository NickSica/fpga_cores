`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
V82h/mp8FbHcv3//3zVZ5VW10Mue/LSt5dvjsUkiSGtG5WaH8H9Fv7j37k+xy+3/pQvfXcpqBF/k
iaz4/vETUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n4WSOWV3uUjyMD/l4IGcKD1bHONRRplCKgax9lu4YRYlORLHEpckVBvOD9geZHtnlLIjTLNUcuHS
rc4oO2K5x66eEf5+m+hNzaPYWCrVKWQI7/tyX0imMAsD4JQXzU2CP3ATsQoldRyYOQZmggmbIMiB
stLQ3uoRuVc4t0kXI7U=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zgo3FUzRcS1G0FRTCr4C/JBs44dp3dv5CUvkYU2vM2fDyGtu9ekJcjDXnFGi3Qx2X0BV1gEyWxsJ
xqQkFlu/f/1mutspkUjOMtKZNCgPGDHkGfwBEPN/xT22fOBwQJUR+Oj5KSeDWe2U4t5UJ4XXcGMb
ZV9syPFreDWYOTWkkl85cAKcf/WXC6oz+tOUowqV4nSLA1PaSrK4ohf8oaOGNVX+4Ji/w6ViTIJJ
OqmPJQ151npm7Kbt4RW80tp1OmABkNI+o6h4rwtTS1IHzM6bJ1Krrp0V+2aEmmqoZkuKINjX5Pw3
P4Vi6iUmJI0uMpdsCPr3MEC8HH4v95WCnjh0Qg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A45QQ9IEoKpoNXpmniz3AuFZmGAAZIhtA2hP4/pi+Iwurx8nPI4ZkKpYXPnn4DfH42bSsec35aiS
Ve+A8f1Q00bmFgtclspinRe4YgFesk40ftn1mzy6g6sLCNXhUm/IIjCSNk+ie6jVQS7STfOdio+z
cvSm8QQePoJjzlJz/jkNhsD110PhDAevJWb+C5fforY6kT0k7ZmJmE7btahod6wU3o7t2HM6+XGU
DDNZ5E+RLS+IiJYVCOwsdqQFDuRaWwS0k8Mk4UuDiVWtU0+QLFZ/8UGJhy2ZDSYlL/8TrrsWcD/1
Vku2N+fkWCj38RSMWEEe5TmUHSSzP7uBI6QwVQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b+wEsHDGMmVXUM545W/2toIjDItLsHFsIOyFDid8Fv6KhzBePVZlc9t2c1LfdAa6UEpdqcx5kgIr
+oVEglJG3R/fb6dRp2mvlu6+x0AYh7FK0My5t84q7uKZ6EPBxHnDds9FLGQdMDUFv8E10WtGrG31
lkto5q+L5WLAzYgiD3//MgdbP+aqLc/75XWIRhw/PfRn4OqyBU7xSBeoK9TDxBwOscUv0cQ+dauJ
dUQ0W2ZCXwF6cP5c47k76Ikfu69J0/IO+FTLKMkjAB7Wzsyqbpl6RMVdJ/iYscNROh1xxo2k+52w
4l9VnVKN7wTWZdW75B3V/MsNTrKb2I6dBdveDg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyn/owx08GdB/M0CwlYM5XwpK1DLRGgNdNGvCa53fvz5ftb1LM2R7yhWTTXlm8iqXlg1S70wvPmw
WVO2ZNZ0csmDdQcX4HNMiokrI2gpR08Dk8n3nzdOhqyFyh79/eVJzQItyKMQmJZNCvFfww0mtX5K
FbNe2x6ria5jEBEBp3U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J8WwILioFJtk4e6vNsFHYZhWTjvAMbsqHcnvhYKYzsY6fpaoYuWnjTNNNxS6JYZj7bKOFgPjdnBA
rKaGPLghV6UU9fx6UcBVLjNOj95AU3CZPEjWGC/GqjGRPxOkhGtDka91PZuOBRTBqJT8F+5qIgQR
vO7WJHaKezpaUm2zbeC7+ShM5p4Wm9L4dzJ1OuUGZNm39p9FbORAZNzAWa35wpfJ6PPOgATFMi7Z
sN0Hg00oxMFCKSg1bxvN3p4iC3rVT+wV6yuzOecq97B7Fu+tfvP+shqnUhodTpF0WYfGWHeK9ocM
Mg7nt62XJybi4Tm5rgYGMIIM0i67934etK5Aig==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AF8EDKLpUnsf5U27caIfzjHsL1dKCT4FvrlOxjBwD3ZJ9vsXwbWO+EJTOJOFymKnoSSFnuslr7C8
ZCAbkJJLJrLXJwfvC9hiPRksxuYzuxWrtwsjJd+5KWtue3gL5kHClD8Tbo/V+Dnr3gvKzMRNdFRz
i+4p8dC6/32xR0/NITJMYT1uOYu0oBFDHGLR02Wn4PqghcTR3gQMVeL0RsDhJibeNnf4Q0NsKqCF
7OscDpis6r9ZAFao+mdpLGI93rreTlZvJBUPh2RcpqOjL/8IUv0iM922KOCZ6j1LtvD0igXehvHa
5hOx0DDcMjOoejqJiwIqLij0FB13lDBsu+fjWw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37408)
`pragma protect data_block
BMP9G5RAk03qFRu5UmzfhEwWXVNssrcytF3IPfT2D1b7tUYr1en2c/ryOoInkpHLJ7gkfkFoI6da
9K4zPon95G0vM8LQxEgNKQ+B1MEk4gLJZbUKSdlMXCo8aKkZCNF2n/6+aTouyl8C3/+Q2hdjqk48
QJWyQEYvDNz4o6pvOcPz7iayyvQ4Gc9KibtMYABuKUao93N/JazXUUb8ZnbGgnd8wWU/rNs8aVvZ
mQlk9rmnPLQPmtaV6sRJmChYlf/c5Qv3XU5vruLumW41uJDUYlv1AHz6kKOgqbVrsmpFH95v8Ymv
fYLXolzHJBvZW/+vENs93y7R8WM0Mgo6BddojDZWYZ875wPtrFUiijrVAekEzhsOey+b7l93t/GP
Qo+kL+S4EXGdl1W4OlXZkzu8J/tyquRWlcs8rIVZ9TM3m7apNY8AvPtbmPbMCEYiKURNT3woAriD
8zZRbbyq24gX9yLeN3pGgYsAqUaXz5AzGDJ/qjp7sEcJFVxsNOoHqAvsAxgpdOxls+l+SHvJtNck
tMW+mI91AuddNf1fEWMKDD4cHhrX4L03yYJibVDNB5UWKn0NL8t8LMHZSozi1krxht9EPehGewpg
yDQ+af/MZyTfYj2pJ91UcW8R1qpGrMZ95ihQ6eDj8NPwvgUBzSOZycg2Rdrcxg+jRJzpOhCxiyXt
YGPVrwCf/1lo9+wvbSFF7po7SsXA3pVK36HDnGdwfV9sWePgfU4uootCXtrS/bFn/TVIVh2I3NGG
Xalc+e/X8Y4r69Yc8C87ZVf8V/p1RfAVrQqvgwijRJ1mDpW+oMDVIJzBbV0HDvJ++OXP5e8AVt3A
WMGxV99EURcjC7kIGqpXqbYyge7KZ7GqTPcn33oxUMxkNqI0x6TvsBsMc0u1J3Qlyn6MovGCYNka
baEwNOFsJyJaWrKgVglQvfegaGM9KhuTze1uvt+ob8MOM+2sbqpAYZlseQWG3+LttSLre2k5vv0y
paa2UGPshgdY+aQBS0ChZmrjsyVU/IJlgtphc6GgDnbpQN+RxewE+Lr7+gpcZXAW2GVFNsM/IUXA
6D/N98DQo9iAFWeaELRUtEC+oeCYZkn5dkvND1euyRIIpw+JXG7WiKgkwY2wWKVnOsTVy8gxGIIp
dkcGN3M3rQJeR2W7IwKP8yrKPZ1GMCh3GgrZyKAKk0wsui4ezPzQI1w0zQvJk4qtHuOARb0Gx6fv
TWdCxiiyrATM0TRLXszRocKn4PXgbOkLOWb9r4pg990vhdW4MxQeaPXIiCKyIoV99X07JpEhF0SQ
6xK4CrbsBtIW4nL9qI+mmnHWpx1GydImxwkPMhOB81T12SX6ci7tyj62FRpBvGME6c3fdUjjlRPm
eFHOejMTwvCpmcEI/EBmDYD9FcZDnJ+Hf6ixcTZHruX8uSuooScyw52l5XFh+lBlg+je7zpGGipn
ObcSau2OnDdP4lymsVOCbxQ21m7BiUIjS84iau1iV08c7qH/hwofK95UL99Cu3yTbm+BRr8jerFW
ssY56TCewbOb63nUfZ24UzamY/O2WojQHdI4dbLHE8BF426Dk+/dSVrbCQ9+XxYYy82UJGTKUym1
B4/imuOzcdFMAWpE//iX0+a7QB/Ef+bx8n/tg4O2ZW1KW14Z4ZGb1uRIg2ZIe2isJsaXbuoTOz0o
6/J+GZKA7ehguLy7uqHnW17faZpXROm9nPdt8WyqeszSmeC0CRrmpSAnSZDnsc2sGb7B28xzBAfA
flVuTS+2nuMS4SPao8SRFZ6/ZcJvkNQJ6xM6mTKkgqMgrR3CvwdAHkOU85U13OYPXTYnl+oePfi1
Gd3blD050Y3IyHPkJOcENgKax0kF3wlQOuYgA7hLN+jB3HyCzOyCI8I6z4lzyGKtC3/LEogET6Qh
0eP4ECwln2tHzpNv1qpoEqLijwV1R5v2cX8tVVtPKUla8o5uAdBLqol3B7EK7GNUFdZRm2EnWsvo
eRJWVOYSaH8nGPTOjnl/2Xs4ibBTVHZVloN8tTfiduoM/p94KxrsTu6YHJZhXz38KevAdhp7ygf7
vopOnzkCcBIkVFG+M2dbMSjMqMJDS24qg3YdG/70OorsAFqW3Fk+YTtgspBhgudWnor9vOKTAqhU
jhJyeOXy/GPZNrNMhNanKvbP/Qm+dBhHTSotXGFzZaXeoJ/QtfdCQz5Dn9PkUEsOtAfIt9HwRXhM
+Qt++qorCTO/uwm3Tt8U200PX89hw/vAvHrJlZ2Sp9RE2rw1BeRRig/UUswbHfpHuA3W4naP+D5p
J2J7EJ/IqXZJGSS3H85iYXBhf7Umci+FrpluTquXLzcN1B0anCL9MHK1zqP98deKLKZdcpb3G5Ox
rsQBcjqyepaO/oi82XqNQ/PPOdeaOTjrkTntjMqEFO8NVBbtXq1yphIrbZzo/JZVTY3giL/xbIr7
KaujKsj+r1m14z6rnVfFP0j8lCyTSphsfHwBQC3VjsqU0yHiYe2zlNCkE2bkc8NvtBpecTZBBpJX
MEKmoJThed6vye9gMKCyAhSkVB2fkOiPzBJ9iMQxbz5vr3VSjlG+KRlO58lNzmKBO+7uUghFLKhY
3df5HyyhTINXTkwJm2jTII7DJ4kxQT+j4meGEqofud3o90SnO1KGig43T/Cn6W+QEuFx503VxIZG
0s9DMQYmDYwxzlOzg3eOy5hl+RMGAGrat2BzlJgfzrfPw/PmJwvJIshZ/EB2e0K8eJdWMjYkUBnO
aiXiEfueLqAwsOfiGH4dNA7pbhqb/qPVNjInXk8CsUSif0a0Awh/fWgjb8MbyrsfzIeMl3UkAyW9
ojgK7c5g08vWxk/7kXmxQIG6pJCO6MZYu4z5qOaMK97Oyqb9N1TeI4hF4Sp73IyAs+hXzKlmzZ4j
GXTmI/UiIusPD8QmCD5ZuDY056+582MMkkkrhXyb0/zaGedRib6aS9pHF8BRGplSkltgL313iCJR
qgn+6ZR2ExK7pzkyzIvxbJv0ZNxGf8E/qV8t2PaZ8rEzC4/cmmysc3a0pktzjLyaN32hKVy6gqjf
Ld93VQ+8KkvA7ntQdMuTc68nVkGr+WYkhiAkXA1c/+5ncFI41gad9HAwSjAsC03meLfL/MdOarfO
lnq/QqknuMEmOAxP7pqI0zwOdzqZ7FCvCZgRxc7w6KPpw2EySN0xq8DnviZ0d/nfDREc9W0dOfy1
csyVv/mo5skEQKhlhOc0+1yqW9lYj/qJPr41rhbyJ/rbIWlQyRNn8tkzJWPyS0rXRB+HhZlIEZtE
itwJjd75ZmVNUGvgYaOIYY/4PlHE827mkRwfSHBY3i7ei1cp5X5l7vfBr21UlV2DmgiILV10VAcI
iIgSAjDgwLY81Zov4obxJ/AO61ZFdLJPXL9Je6wMhehNrUalDfB+fIB2FqxAtQLPEbKzY+UQ6lKP
yjMLUiXONrehfUlej+yJ8XCmjPSvGcP3m7zRqrohokt/MI+PKcg0kzz2+NZBi4RqdbwSJG6Fmq82
loe1h2ANYs2ALEZfLBnvDJ1ZP54lV1SIKnTzXIU8PpqW1l5X38lhECQ3L5LZl3IpoMPZd/+a1HeE
kO27SPFO4l8W9hK2uuCuUOwhq09m7CHhK7fIf45jNXXTQ8VTA1zHrymRpBhAHQCQTh282PYVEd65
XlLkvUK8RI7b0B3SrhN/taGHtP8jHOpWkf6u2ylJCsDlXDzifn4fBOf0pJguzgQbKENOT0ZXHjZG
5RAVb4j1UV/28r4t6iunOeIgtG/4cO4tqQkLvtLIxNbJlgp4Itz4ooB1oWNORIXsQUKYNIlluC9D
jWudeM45Y5JNkpr/hdLupDxB+v/vP8sw2gaM7qpt6mzELvgBTiW28WI5R0SjGiQXugyZbLsiUWim
jJiMem9AxKlrvrbvsCxGQJEj6xWjVAOcUKJ7qqNuxBTvT1RYbaDf6d1rI2MMPAycMJvg78AXPmkC
GanYk76aRSMFV2sAyy1/1hQrmJYFD2MR5loiyas5HHvE0w1xd0pA3zWFdWeuRzUg/zXfMPsZT4xI
OXjxeBWpfvCqtm/WlsARA5e71nax1if747/2mwyBR4S5Xk80PECbL/BNJWbbpfR2EbL5/F2wncE7
RrOAPBOe4nRJ0WZuQM3KdoZYZkJfA5UJdonND6gKdMtx1pjNo650+9WWPeRIy0F17+j2lN1HaAID
cDfuGlNiu9MF1/TSXjpAj7wiPmnAUvnDwJeoPBemfISVmOY+bFB8OLDronuB11A0517ziCbXk0qI
5ZQnYfA1UDePnTAJAOEK75cBW84g4iBzGFMKk6gqHond8opMzq+5R9A6JCPUSWupkdx+o0Wwog7J
Ig+KnmHElFYep9IoV88NvE3WzJXc2uKx7XLMg7M9N6Vtbxvvp14ejlZP2geW2rY5efT/f6dOwjZ3
Xb/4G+yTlUCLAgiE8iUrFnXaPip07eo5RgATF0lgjPHr7aq2Q0pkkmStQdEQ4cBGDdvbsCO2WH7s
IpzfBXYwWrAlv41N0oFYt2c6X9DSg3GDVl0I77UXQpkQ64qjsZWAqzQkr5iw7nia40iFh4Gw7v3y
kh5A+KJr6/aJBaoIrlTkok63rUOPlulxklaow64vT0jb7JeIFjHJm3HJhwdX89OnADJBGqHB/x2f
H+Ukqs8COvwj1t6dfN6Ihh+pfaY7DGSjAU2qp36jI7a5TDKabmbcXhutYCKDLBVzEKu5AQDLeBdd
yd7t10qnDxrKJ8+EqpVPvR8TBqWphoocbFa0TCXODLx45Ad41u0y3QAT8RpJMZaqMDskhQ3dFI5C
VA/WBwGBWowSalpfaLeK0Pv9h6SeYrJOu3MX2wpBCnWgREFg4ckxcYkhOy1xGRbdL812eAp3iePf
iROGBgV3o42fPtNK9/SMvw4H3U1kLIjfyoZatXSjLvbJTEUWOm0H75qhvpJ57ulsdtUc+S7Wmd7k
nh+XrqPAVVOvt2D/11nnCFKc1Y6jEsr5ABd6GkfLw3ZLRZJLLRRIWAsH3/kgWzRXv7L2PA/CLl+D
inwBxd3uAOlIq95O0603qOVxceDph6KrJ+vTNgFTUhASdVe3VdfcIJx8VmGC+cEpj7J8nTyWxluy
kGWeIhCv+w1ek3NoTeEKZPoGppwsMR22ec8jIsS3/NoxfZLhS6/l2FiI20CLrZu0EvXfur6jiuqc
BmLItI4rPFxoPqHtYb6rOJVx5KehuCqLJuh6tP2J7nf3vSalqJdkzILqQWQ6lb3TFI7HSVA/9tjG
qm/Wces+dxQug9xNIAhW6/nJX+mceJ7on6PhSjih+U5IsvT1+9xpYdgdzjME0IQ03kbAaIo7dGwY
fvemjMAGA2g/WvLTijXB60Q0x1N/VDd5Y5R010LfVIRR7Q1Xc1WoAwFtPy8GnuKw4lBohwoEGVw3
FuVzpBSWhzVwlV+1OiwyEii0cqE4f09D85My8PMxQh8FG+X2b0DTCc6X5BvoCWpwebYRiL/MpgoS
CVf077lsjtVTUihunHtzWT/7ayQ2bKA5rvh5owHyiFhhtnil9xkFaA6kEcXQyrBVtYeHLT2uxZMC
XDlHp/j2v+njmxubSOzI85tqg5Ci+3JCv4it5YL3k3oBTquxTrhGowFtiYOHkMS4lRIpLh/jaQiT
MCuGljbN8tmapnITrKEJ9tfUzFp0t/azOcdFul42xM7o5s587oxUlIjnrb3h10eHbEz0K0RNwPOg
rloIdihx9nj2hnWCXCkVllxVPuU3XpWxhxQlElWuwxEF/7Kq1u69T2zxmYzkApkon/77bm6D161m
evRQ8q/ijGnAqVScT/RFpKceWfmkP6hjLFCBkQ/Niz97NPEqomeFFt1lNUsOuzcNmzrIH1C7c+HU
HGJq0p9Plz3rE2uudbxFiCO8PJow0SkP2Q7UkAyfJ7UkaThqNHGwLHZA2d6IhewFaKDbNKTKoq3W
8XRIjLJeWkl+snhQBUCJ0cSC7zxpiXBnMhlioREnXXvMJkJ1bu8ojhJTU6uMKpwxHjHqTsKsUWdR
x8pv+cCDaMjNM6sOmp1CcNjwNg3c2Mq2z0P3Z0ekEuFnqIbG6D7CDEaOkXKrNWRKvXCZKAWQqaMx
gSPQM7hpdFFYKzb1Oh4XDjIEGst5vQsxSHauswzvpuf1oTN01qMpEUlnkonWxHRdlXrtomvq4L58
mLqpdKyx8rQVy3isxEf/2m5gB2NtemwfvPyUXSgqvL8di1vX6bdrcI+V1Rid4WMJUqk8u8+i5TW0
ZwGpvuSdFp9fN48AfFwmZauKpIw4USueGQxKXEr2lJFb8JUdtYTkZqZ+SV9lKvCvOSnKi+8RhHXl
TI3OhaKBxXLJ+o+eZxjKaKMWAjKGRTlSNpZhckoC6KXRpCTo9j/49HYjyHs8FkUv1m71NJvEWozG
+yL1Qs+HdB00QM+uzChtQ3mX79lSN4aioSUBUH90pTYMcLpJjYVP3za/M069K78v/vNsLjy/nnng
YNyXuciOX2dP8pJmx7FrgNIPbsRNTiHrQofmwDax3IxJFJweYwVIwVdy2ODd5hQaIE1XhsEoP8SQ
Mt2fH2RIaJU5WvOUjnRdbpu6tvpgyYASDaEEy3+ec/VfmGSjQyEqZY/QZ9rPMI0ez4QqfTiWfqiZ
nbKlMPtNffbLw2zPli3PlrJMCuGG2NOvvhhW5ELUmcQ4/Qi1CVoomy7MvgoKnuaLsDb48uyXKrWn
4yWiQyT+jpG5d9gakNE2AqkBEBCJjZ4BX25t5N/2ht57sh9oEdiXIjGPKGMYZG94xQzWqqobVI4c
rIIEy9MceqZj5Ip5PSv5L1FKU9yaLSSA1gcGLqk5QehgSu3JSN4i1n0S3OM8zDvhuVPkcZ9aDbxT
mFwGuY6AN95lbJORk0gf/56SxxJcNxdUOZDrTl6wmv7Wv7Ip/22VPu6ePd9VnI3umzBqEG6W9Hyv
Kyr3DgdxYHzBwRBucYSUSUHbS3F1HbDnDipTFGrLq9V7vUi6q6GpgJJxPAouvPIHHu4dJbPlfaX0
Iv1Oi7Q73l0Px4TwoAKLeNw3VYNVLlDE2moakTEkF3Fzn5HOmqx+vuP6JFxowED8FBZzbspTC21N
Z28Hmqc9404IYbRRLHNOUIKde55p5szQElPjz5gl7XqORZ3MO6dHDa8EnumLExHlm/M8W7u6FIoW
+KyajKvRYHp6E738yAfllBfGl0lqostNEn6LFDiY6tpUacAimo48K/GspIEUmQzCGNJwxuh74xSh
n9RD5yYrkdPCtC32Aq//WeNUv9vlKymVpbKV7DxHkL2AKhdIsjAuy1oQA/228dKN8g11GD1W75qw
WJ0m5Huk0m8QsqCAKckqz9zW2tnA9Ys3t+swGiKRFkgp0LgLgey6vIKZ8KdlV+itkyDEcxCFlctU
o9yGDyNaVkySW3RI+Bhkxk1TN69x9SsWFCLDfITO0JUMjmF/K/b59RuMVHHNZIPMRS+3eS7oKZ18
quDNOwyH9VCVKJh8j6VSGaT9XcY/vDyZ+ouwyMGA46NZ9NuSvzJcxOfgWu979ScyxyJcpmU90o+K
J49sF2wh3ZGU0udFnfpWvGGawRIlf9Dym+nwmVuGHVLTZGOOtyEQmsLtQZci3Z3aNv/isEKORnJ/
coEOV+vWYdyK6mrDBtGGWgPUlUUxxUiMpqQaUe8Sum0UAIiJ+AfSz6tiEnB/ObL2q4CZZD/ol286
4UIzhjR2fJPg09f1ywOC0XyfEgfeynwjTkgrcNPONW0+mo0iLz997znxGL7PUQDmLHh8IAfTPJlE
I6+uCSqS5KNFxUkKP3+XPOo5KIkecJVOdSGJUbV/M0UHJW3adMjYpNTIW875sipbMtAaIA8frzzD
Hdh4wqpU+qoCy9jsl9n7oxxRAGMUijlkYWnLV/+NzMIWeD0Gj8EvjTvO1VPFqF/9vA0kt+AqmNrp
ws5IucrjrUblQoeV2UjplSdhKaRkePb39TApay5sUDi5bEv6JSq56TMm5Bz0HrFh3WpXsGq/IuHi
adliRpRw8ZsfOw9ZZrv+Y82b0KM83YOi0j8VYgtN+v0tQJL0ve32vlzhasM28ahmg8JaqhlXAITY
zDD3bw21E0QlDeJfxGYXjzyEPZPLVqXsrq8AWQXfQ8vy2jt6ICt1sQjlJ2eo/9kgzaprsah3sXUO
EX+P6uMcudh/veFD2Df5CEuBjP7QZifqZLZwO4Z81QWbkyKm7FapmPnIc8SuVolVby11/DImN+6o
KcNiCAUr4yRYWXj2heitIT/UwXT7r2QseyBeWL1Opq/5BoSNgmvJbeg8wTejY3x3KZRA7u57JYip
w7tnH1Pt2rMewVDpz/NNLw7sKOvcYJw6+/rWpBbw3RAjgRRXNo/pPyVz00l0dSLiIi7UPOwCymK1
8qiLnOk0lzwVJay2YAfDs2TeGJW84S23Rwl0JPXKShz+5Z7aalfuW5sgcN3r9EP6Md/qHl9xH0OK
UhVlr8/udS2Zlnln/U0sfnxFIVKFcnGqWk5UB1Q8ZTGd0Atdx4XE4q4+YPB1wUMM4JsvLDt3CmSQ
iVkZaE3fW5m4toqOBwFJGHBVMqFq2t5HVEahMST6yvj4FSxBH1u6vwW9EGvmiUKnDF+z85v5ma/5
/4s9D5RVu5loLE4t97DfCEBV9ALkc7w0EifNpf+b6EeGvJl0HZbXhtIm2A2jSI6Br+mUm0wAVsSQ
roQQNr17V/fl7Pcy+1w2pdK9MN2OZ82Nq6SAAqKu7+kQHz7pYu7wgL0b6LRiIN4GVe3GJy5r3fnP
1WSMH/vjh52tyq3mJXX8iSJ/u29ClYlpmGxq09oM3GKfIahNPYaax9cjwXMsd3NMjW4TfOfpZuAU
jdvwgdRkJqmjmjeeJX4dN6NA3EnlMsyjVRgYFBoc5Myn0wPpz2qV+IpK2bFJA+/PpXHVrnG+zGP0
KnlkQHRZPRUr02cn9JhWUGYCks/aBCgMX1EGYMmG771NJkTuXM7Tt0vTCC5k+MtNoKA6Lb7UutjS
sm8w4jUMn1nDF1eFxNmTUkwWLslAK7nHUtn4jmQlLZF8BIBV9Po0gn7tyOnZrzW6PnQy76pnvcrY
l4teKtIZ8PHqXGxg/NBC777cQpekWyP/LCtwUSzSMrePJ03tjQIrmCcI6eqEqA8qcffZffTpJMoR
EP3yI5WkhaAACie+nHdtd2KC4ToBr7WrNNI2/ySzjTaypYwDid8E10U6Z4AuPLWccpDVtwzrmTRU
o/PFpk6UY/sT4tcEbFjnEKvM/qonPDV1LcyA7mz/+glCKU816FeRwy8Siv83TqaS6japj2GmOK6B
oqzTnWP9LMYysYokfT/kpHjo9FQgxc3WTQ1y46nZJDgNlfkxUOfh+sViKb2JBCqBlcS5HEPTBu4o
Ua7noXUwQT5tz8xOSURsrSNRJECXKD82UFq5jnbi6/mlzaXQW0BbS4X3LZD8YFCJt8bfvbx1hKCL
MEIgbkb/Y1bZdW+H3Lfc3z3nJcMgBQ2/RmGmuhGeyb0NxGW4sFscrlxriJXwLMNC4iGj0GILk26R
ycDP3IroudeiH2m9IbPEtAJjXscbgJiqPxf+phEofwk5YThakQe/fEJJcgb5uiVZUmkKiquzoypB
73aKC53mXJh5eQSkih7yDxsWqVJb2L3Hm1+ru3plu+JIYW2cQNTPVDqqL3vgiiQvpVoLxHzeR720
BP+e0wSMpVAWDYK7rscQzUFg6bu+KOqADo/JoRXrn3Y7YWOBZiKbk4iw8YjemoTibDf7cK5VHKiC
d7FDFYKOgvcTUH9K2Ad14zZCqD8nWkHsFTdBx/uX5kUcyHTrlLfZTmtMzxWjtkcO1xLLPwaVCORM
zCEV3jb+6XSMZ+5UWBT9YzqAwQyOiKar2QMA5P70N4AC5JUhK253O2mr1QypudgtkhQtpS6uJS0f
x/gbA/+HQldm7blJ7Cq3KN+Q25YXL1x1CNeblZ9MTIS8sCYqRjakvJBEOO5ZvxPnFrQNeA5HYH9N
9dv+b8yjx5pwfLug0Tm6ALNP8ybK6YhwQEfIbnXQVhvUo7LL8GNUmitzRkQh4RwYG0MerMaNFmUw
SJQ2vwynOhs2nikiFg4cGt4QdUGfgPDMurFJShwKTvhMYFbamihEn5OQZqj8qtRyzqVePDco0yiU
SIorAkkVfdTYdWLfbAGH2SYs7PKAQ6EJ0qwYCrY7GP+Mp4zviIPOvpCKhe4oPFiAAXgIe5hNYB0K
MhkRd7sdUPeTkxzKhC3kd+d2utHDT9eUcZz4NaTWORdN7Hba4X9M7Lm8E+ixRy7E1fgMV6Z6zoa8
InMlyBknqnFn8zQ78YddRrgrOQZpjuVbGaWPF1S7sutLoS7ybLiozK+NA8uMa0+xHi7IZoQPe8ow
5QIJJctOzRWuYJFsSZ7MevMj/fgQr4LONrpGVYgWEihpjRdF+XnbkCRcveMqjXF5swn7NmE9HJ8W
IkxDifsMTbtYpQ5UzLmm82ksStGeIZdjt7nwC7kG1iL0Odx09Pb+hy42PNjIgIhjhrEzuB8cRVR0
/ymIEXcf4t1x5Gx/C2QJSst8JA1AZX+O540SYunrGBmxiB0cYNQbV+pZGTdth8aCitEjK2wEP0qJ
TnMAgZ2Ag/sUdCW8cHXUs4ow41VkTehsn+FceKBQ/lZyvlqygHahegNhgQIGn5vUZVdOfi2vIxpS
QRXf7pqBzBBXId2skfqPTYwLUJWHWnsuKMRAwSF5/wAjhJxek+dIBEwiDPhpiv0XRi/+YadXvvvC
CJYwcAZW23mjmZZ8Zj/KYJYhk0ZTWGhGY39Flt9b8iqqMILkJVcqXTH19Yjssvh4y89tHkmRAkKr
PQw6YdtVUowfUHgCaLvq/wF/TXWYd+o4kKLb4zTS5wxeCfl+R1efNzRPYrZ/35uzKmXsQO8NcJLJ
Lo2RhunPVhcvT3xZkzt0ts1Xg9t53iU4XhbeyRSUplVO5yWonyDMdQDkHi+sjzl8nd99I3fBS9Mp
Qw8jiXdcwfsYq4QoKUea3M8wGHiX73wMlQ2ogk+r3GzOxzQMW3fR4GAFZcogpKJxBrEx+NyN9S9t
S3yqpK9UIvohG77vRdmpZh02q9+Ym/cI+38q9OcKoNSJeqxKSTWtR8FL9tIUMn3zcPmer01JKscm
UWXKZmTeQXaNgxzE7tbkyZeed8vY2k1JAo+/WED1m4+FJNq4eZo1/EB+QrIOrCSiuawS1iqAFbnU
hbo6TD0L/Z+EZRTEBkNbRA6WJ41j35tNV3H+FGuDWjHCUU8qnmWJffEuSf/KaiUPMjODWXU1Htdj
b9L3CbrfDTooA8e4u1CrZBkyGZR/LO3M3/B3gSooPLO8Sd2JhMXlg+9Xx1DXulbzwsar+Fp4lb6G
RuCqb+++qO8XO4eLkA+eIT0i/orXVnYksWXaK9nP4gBvQeM2fK8PbFTJ7c1WshhsSIj+8cYCgrnf
JC2hbtDsnmiESpO1sB2yOPf7ie1bZHUj2g9x1SN1+n1qA6Q63r+k6pCF/kUsUICMPW5JCCVDmHhq
e0wvy2H4+sa8vuyRvuJ1v7bSdNHEOtAg8C6fU5NSHemUzvt+60JMOSAanvIHraSgufAR2R5VKHtn
utkEO2HmWul3i8utPlNx2PpxV+asZpzf4x5GcRYvEVJfPN8phYcC9l3bZ8DL0VmD86hDPtJOtvQb
MRixUcgfqo5F/7AJ7aXLQc2ZkQvrr6Z5ZoZmLIDSlUEUFo14uc34/X0U0F4eARPfXtpzo5LuNPr/
2t6OZ69O5nt5YOOu7if6EALAgluahhMLVNkGPZBnYK9cXgRtjXebxYSa8/iKzVgJAfVokDKROmuJ
/lenener7ULMlTewNtAYRUK4LYIeRnHXIqBD4jgwA4fmuCq8YnOhCMgbg1XfnIPg6XIzuuHL5bjU
eQKSkgKFiFjHFx6mD16fDuG7X/ZAXO6+iFgNzGau0ceehrZVOWU6wcbMrqkMj2hAUhn/IvgxDnQj
4cVg5Qr/xzRI6UZpaTgZyJ7rYvipNEJUjvgdcpC3WbCSl8zrHiEAgQB6a5xe7ltwChPn+TbVzQqK
ttSRX6rDqfgBle07KmH3UfJ0YBmT12jjn03gd5Ed+o4HhO4L0NSFAcuN27RhbPyhDxj3V8bein/f
enDd39evrzSGWx6J9hHLei+C56KrKdPyngtj4BYgz5ItDTUUhh/Qss/MVx3wZCBNiOCsK0Y4igI2
j0bTmyy+YtTZD1qXgnx5YaLOjqfsIFC2S77WkKhYKuceC0qkcYy+GC5/Ra2NZsUaC/EcazQKMjAI
bKQUauGsxtBzTLLsgPyLhJiYKCJxF5TYijK3X37XVOKwv7BP4/tP9OSCKc+O81YNakiYwS0G5flA
NiiqGqZU33A2KGw2CTEFPbySZqlmhz9rmXKu/GKWKVQtAmd3tg/vyuwlJ7rezE1uLr0kzrizv7Rx
0lhbqwHYLjauvfrcDatElSZ6SJHQMR1OuzSIioXS80c/S6h6UZmDYwz3W/AF3lMW3d4zsxWcMRJX
WWPry4r6SLiZvl5tgsGihDb9LgNU7v/ce0D21lI2ZDvLMa+D1CUViyBg2EzXKX1FFIE70rXi8YWg
FQkNOJl++c51Kpk0L/a4tQB/+kVdt+RsZFrT5B/jRn3rmafaW/9Nt+Zk81AS+trz597fe8g1wwcA
smjlLHWz9O3cWmlVypv5XocVlLuR4lHTmV5PLUP8K0mLNipglPgCpzlvVn9qpgyO8Y1xjz+PC3bY
SAYugeGrXDjHNedEOGn4972ymStOCBIXuSRfbw4ajuV5IEOfVxpL0hYRISW/0BOMhmjdAFhaJ7ZB
654OwZL0iOA3/3C+wg3pyV4+NkWlp/AagN33uEOHyrxwFhHTt2JnPzkrUp20Y5C3M1LLimggaUpO
BRgbIiJPsNzVRdbVGtLbdyzcoo0IPz8QlIdAWQ+jkmeuUQm/42s9EhtsvlmQrbdUy7YgZendiwhs
pIItRe5z+3StTsmJcU2gdwH+Xw32rCqumxGjgLxjL3Fbiv7hx17Eg40r0A9RnoSG2cy4oPtHG+2A
tvppEuhbM/dy42DHwVPmjnQkmlkWFRbDs82Hr/B47CQO1yx5p0XXPYVB1ran4nHGmT26USSVqEOv
rQPTI7OSQIDUsK6HqLQU0bZcYG6QG+Xk1c1AGGjVdsr99PeVvNv9ZyitoRJiOlTyb34pBBuNWcpG
lhwzvKtrNWMJnoCl+7sv0OWQbOtx9qs8nnVhcAsmGWpnkk6/Oih1GIHCs9+96zebWPTWS81Gwv79
9okvzchV7M/XyTke1qjRoP47/CiMCh3bkdmedBGEisQ+kx8fXVqqr4uzq1Hc40JbmWvxdPDib2jl
yFPcBctXmWbufpndfWLLXgSG6oWFCYFt19Em/qFIilkd9lqlcpNV13KLh0yGi5/CstZm/MIpddmF
BeKif6vohdZLG8vNlxIu3tXfAStkAtH49QDZPmVUzTA2bx0Kj6Dc+0HkecLBRlLT0rK3+9tuQWMR
OSqWkKjFxQD693M6Nt/h2HDuZPrgjHgJApRTOdJO+luW1wu3p0Pihq3JH+Syx4ekPSjtXrkUvzL0
q73ImVg4KDNahRDxc+wE6xFCjwWjOz9GpSPEoOKf9CyFebQ4PJVjuBt/oGGOesX5UkeepDU+FL46
OW+KLHa6PonzL3/nWd3HKLXh2zUMe93Klb9/VsHbFf5OEAZAvKT3vxVPiMf2JLFjibG6MTP+suNV
p2H/Ls3RXMg4/HAiY4sFK4oI7aujw//xQyaoDptmB+NWE3gGiXvOwBwknC6p/1Z9Ds4+vG5Gj4bg
oQGzCLUkUJR5J1Fe3QAKlFjfpj4ynpBI8Y212eNIpPkZLJxCE+qD8uBIuuywWkPxZIHWeu6ozChM
QivPxSRUE7uXgy7qukZC83v9GfGBaXQjoSq/g93PPzDIt5txvE/p534cl4wQKYDj0WtNRr7riPFE
D0v9HceT4jW/dE9SvRORZtC9kPiN0ZxdclvGJoz9dOQVzbCNajIU0TfS2Pk+Q8q6gG5nHJVprDFL
C8gCT35ED/7GSRoiEHdj7g1mv5N9Ma/1s00qdgTy34IQjgZSqzl9tTHWkgK+OG7BDkBYm7Yei0cW
DiBUpC7D51CwF1BMv9FIKkG1jF41sCD6CupP6Kd3Qor+CXc3Rb29pZ0KGJY4tKfOkiD03eRvGZA8
XTy8nbwnZa9itOzaa+msLooNQTdJPyq98mPFDF0rGW9lCxiz7iGO8EYuM/Qc8jnErZtEC+xfWuNm
6YuFE7i0A6D2wCgRybE4cqCNSCLqAfw2AL/88xsfcJrUeyfxA2VRu3hvVk7Q8NvsZcYUD3Xtkd38
mcY04IbmiO5tfga1SzI+FUSZvgGxN0w5Z4HKkokbfkEjowCZjD1TyzmVRRGHsrq5bxYndnwoOiMQ
PZTyqGEqPqmXBqBNt6dP/sIdOUX7B4anXwclhHsB6WuKLcnrksVRRwDDTGAHLsM8balrM7V/7zY/
lab+v5ovYrooxpOOKsI0VyhAbGx3wJQYBVEVSG2Pz0l/A5i7SlljF45/cIqRC0yAq/me349pZU5m
kL5NI49exIictiD/kVrThOSUhMr0Ldp4PcBtGlNUm47KPJC3xgmuDL9ACtoqwRfqjDx4siJ1cSW6
Ps0K3DZEeY8j121KLlrN6KNV5DbvBoNOBZMlnTx4IQapBOsq81giumbetYtFt9WZOkoFKTvtGA6h
hb0IEzRmoBkFmxLfTlcVRVqSvmoaf03f4pHHk1yZvwvdjMFHCGRegjSJWntdRONe65w3EXuAd/p3
ZjxfbSu1e9ZDyrn/3KjHD2hXZ+vkhE0Z1Ft9sQe0Zg7j1qQW5Vf60Vs19Kt2pPcFeUEmRNawnuow
YbgyDdj+EC5vGgjPm00d/a2FKmplQP24EIhuJbstaIoVRFjMnblCx2aj2/R4e6SFR+5FUduwyivm
PnswwafVA5OFnlK9QjB1S8ff9fWKP3j0nq1+Nb+ufRsRBJdbxAPnAEAJQ8IgzdqSJW1vsIVJYWMp
9G7X3haVgGxbVtNn+4AQ9AMLDTEWp1cPSL2wikPc1T9UUA8q8BZisCtqUKKssgKpb29mqd0vY95R
3L2qdU+eV5p+WQ082bCDGDwdqG7IjpDWErpiWcwhwnS1dJ6Iky24Yv4DhDUZAS7MN4q90pKHYrgV
nYO5gXDoDDRNg7dVN//IN3lA18vQWXZgCtkjlgEsKn7j/FhVHWQ3GVQHKLjypW6Fuc3sqJTFO/He
BFnfFCf2U40DiS1/PG8ssQ6tOa8Mi7OWO0tH6aZhmP065mom6gnvssOmJAExLc8u05DonvwyJT+2
je6xr8OxWr7qB6jDV91OlSTNffsEGTa2Y3np6t/eRtwsqYB0ksfmYRaCcStsBM0aBR2Lnk/f75vD
Nqesqv/4XeI19qr+sucu2oxvVgJ3cvhSdyjt3snE2ca3CKHCl4r35fsGMdcKDQpOhODdYItEVwfg
d3mR3r/iBxwROqlAvoJU5EBx3LZsj1mP5vROh5nB6uv2tMw7Vuz48ZacZvo3MfAhCIggu/ClQF01
v4a9O2rVj1BNlJa7jaDlm19YqBmPf9RNhl9Um7RHW5vDXU4qdApHELLFcpM0c0Yv5ETaaiaUVUL/
MLMyw0dteBLngo8It67jmIhjoT1cn3cOEPMlxwIRudtu1VtHa1J152yqqtod3+vA/8UuQ4gbnFax
tTqS7CD5sLhpstmNf6EotMSab0wuxq198tTJ7Hdq/wfH2M9pJhmYn/WtQrpb0PVWj09AiC/djnqR
zbnRYxCLHKuuDDXQtouY8mKC3ev9pweO3liLa7uMtjeDrhYwe7tCoffV9QypbLOeEI+DViHqmgSz
ryCfbTXTVb4WtrLNZdEUpaatmybF6mSoddJm/OsIi3X01sNWlZq9fXcMv2WtjjCiutRG76qRij1F
t2KPpkJUatuYL1Fc5FKxr7blKuSpNZk5oU9AhcRAp+DTmN9cJ9g+CamUb145IwSD/E92tWjuAZ4P
wzWu1CYQ4yNKLJHtkFtDgOdVryRViavOGB7z8YgHOzfwVCstYlLmOWFwLUy6IgmF9A2+ZEtBkX8/
0s4fuuxoJM43CWb5GYLoJh7nIciP6sPA5qL5NYQydTFfcHlaom2HmR4/HevNxRwrFxepC+TLBCmq
9twQQiKlQgRXpuab/6RgGNTxhzzSYEBGDTzInZyQRO+5AETARDxVmENQBnCZbwNzmcIcbzgcDCuV
bI0oo7aIhj4Swkb7s6OaeekbHamRI6kitvJ1ZJ6d+hbsJYbAKvU2AXmBgQaMVscWUsccQyCuulA+
kZeRmskzxa7VTp0daovTgjheKXuHIv5fbkRsN8DlQXavb4cbCnTELmSopoZv45NBIprtM4SzZ4WD
40mZsbxu7c+9zVDSz97eWrGmGdDNJRlDB+irBR1tRSGOzxai0rRGwIQVx5ED+SfAiB1rE5nvQxVh
EueHwP86uJnij8wxIwbqJCMrj4YyMlUUJX+68fdqrQt5NuYASgFHQEmuL5vkz7RBE59/jM9eMrN9
sRWrLadsIQsA9hMQQ5qvOMi5ycOGBySotXGoIubAQc+J9tESPk2PK+GVWzwYSvxR29/3h7oA3yNb
/wdvatSeFFrqoeKdKyORpylv3naGD9J4/74XH7eXfNW+AC4gxNtZ1PQk7yVI0vDRcSISg+dpJrLI
Nw3AYDE40o059FMVfWUYLXyEEEuXWy51VDzUxk7oC5NscYS9mL3aC4CYiXScmKhpVKfw4N/7KIpf
w78sjkz6hIBzlrgKCFSpNwg4AlFz/7gameniD8S8A9dUYnn7IPrKQyN4wUXBljwtvXEf+2dWTxRt
JSmlXUwhkBaEBVEI33peONClX21nBoldWTF2L3vG8/bY02oH4cytP41YzRAOc7WVrdpOGJZWRKr8
IWhzWrEwm5k3GKci9ap6dpIE+Af66FVQa58srIlNwzLqPZAU+EDlHOoHayAVeXVq++Ic4qmKjvZ7
mfsGtbG6NBhVvtYxGMRPxVAg0ugtWKdDlyk4Ke8aoRBRBF0G2zY0/VlVMez3x2kRyFF4thkXxNDY
9EUIp37PUcjx6ALGR9L+S1DJzEihdE/ukbiauMwD6G4NFMuRRfLT6XYRIsuVjyflEXWbrpYGtQvR
r4zD4mKh+3lmW+kyb7/k2kRagGZNq8BmjcOmVO7+GVf4fnIPkbtuehaTGhWXOVI3KUxUatVC2hIn
TRDBcXW9mOWxhQRxLxO3ktJgwqxBhfVUC4ftxorEbc7ivlBj2UOjPkc32EkBUJM57/Z44DKyRlEr
GJyi0mHpcHnfbb348MXgmIEKgRU5+TTVwfKCwhbM4H+ZQg+fx3InjwwKsgGMczznhQ0tBSSlrsDP
/e5ge5C+FKPXvhD2BbqTSmnpw8R6Xmvfhrpe1igDQPlWqm39Gks6ZsGi3d6leHGPyypmM4SuMz8D
0fL7g4aoG9SISM+H2FcKmobTYoMK9es44ekZwy/N4HTCyiCTfKNcjwMPIYeRVMoi82QLbNb0fkeG
Nn/2gHtmojhML2Zsc6QMUc7g+29evU5aVbKO7LnUI+hOq45sYz/bGg0OzSdQfBdl0uKpi8z52Cs4
CVrFcwKcMJn9a5zWtXGqAr5BUYyS+mDzbsUq9TS826KWjPrHiLjgG6JAOcA40HlSqLOYtqrjW0sZ
5mWF+tajnWJQsSElOY1a1NGZzvdiba6q6u5x8fFLj98OPABpwvnMoCij/UvsoHHKYxBOu1hk+VVq
KU83EiRFzayfJLatPB5+m0pz0AYQy/LBosIUqZjuLSLLWbdctsf4fcA8TuGXDg+64gVbD3JY/iCy
8+befBOXqweeNWne43nQipNRQgL71wnwnfCmi5tEi83gP8/Xw8WcAf7Evj5ejas/cf+fmZWhLdsv
iPMzUOEnwNYB5xgZ5YOHdn5womeJNbzNR0pYt0S8wRtE3zXuOYuGniE/T5kNCZ4lQjciru2+Jeyr
bP8ngMtWaz59pDsD1wX3R1UiXnxqNCl+pozhyDQy0TsmP5d45FCw8NYe7w9IyPo6wBqfStGprOV5
PZLRfCt+PGu7O/bDHjOzDEw8eHmwD9B2R325OmRN0CZ54x2AU6DveskHC4y7vxA372gElcAo2Ox6
x0LDfwvTOOSJxy94Fd7gOpGYR43TlVqeBcMVXvQVhtSr3FJ4uJB1QqYAgu+U3E4tNvvXQ0hTxk8M
DUfPxMbtmoMVyut0QJ/Fq95yXMvaCdELGSMHkDM5AS/zdNsw1RLdBM6StUZbI5GYlsHSMIdy/AI5
jVWRae85Xe34xQR8hPa4S2xT++W+TkleDoWejyxhCPhxH+ILTlyk3m89exwPnERXrmBm9kRFiHGi
m16BKq4ujTj3RD8qPH/YHMRO3LB5DbMasTkoD5tq46SyRDjuPUQBCc2+J3VyD+/8nY95q3mmrs8l
l8RANehSUiLpcewucQuWNIY9M6lsXwaJEHP7CjkWbiMQPeXObxY+i1f/BA1KM7azpzihipxhpImk
MK/ManBjT+tjU8aEiWgq+ScVeNSTvGmQeDU2gFOjQiex4bEq2kbh6Bv9V2tOp9MfobFwFay7Hwwp
w/UsYLRkpAWphy6bt8LRpmg/hhmIFr7ZY57AcIXYlO+niUVbsv4UAgMQzxlxcgmBnNmlonggRJNP
x9t+mcIBSpkw6ruHSRgEjFqllDgM6bj9BCuHwkWqvWiZUqMabO7HYnazkWJv6eeusBE/RAd3jf6K
Z78bR6CG/dBZcToIZeC6HlX4qc6TegPWvAe58MrdWScipnFymyGJ0duvBklAIAFlxdJXZ7aAUfQk
TCRTY29YoJRGm29Y1Bqodki1eZeGo/qv2JUH3fh5Ll/dRHF+Ymriyp//SdIL/tn5GSmM4kn7Np0X
gUO2qu+u5i1+bN8R6FFSYStSSkr0GWHMuTgHPKM1qwWZJwvk7FV2/wxdoskOe4e92vCkAG5B0tEK
1hsviyHH1Gc68ZMkFpDtiNDnUN9HZgu9IDdS3v37kJXRIxb5uvTg9VufT4BezhNV2AdDwbZVYBgJ
a6SCNU6Z5vspWxPq9MljmbJ9Rz7PRbuiZok9vlTTcDbIM979FtYSVV1RbCHiYpUMuZu6iKaomsdM
wRiv7YenwfFkxym9KAfiAhiCTzVg8L5iZ0+7YBpLRxV6uxQnaH+f+HWggTeO6myn+0HVYno3r+qI
2ibVb3E52x7pzUvSKXeZKzLZ2chj1Z7GY+YzwuwZMFJGcxTTeqkcJzxStFWSKE8y7bORdfpC2FQn
nTK7WPWXv6BsM9vao0a0Ro/LCDRh+oQvyCOArDsRYPfOy0ldjtOAn0sXkSIlgPUfOX8kid8PgbIb
HDtxf300+i+Tp/3mKwSuvBc5rsDLYoUE0knhrAoi1vIqzIpdwae/lVkaxHq8wcfG9JO6qEsUFvII
1X1S4/0gSRaKd9vVlHJJ3W1HDsMrFXje0S1ODJkkHvzHcEgep6vx+cSx6ompi6MvuLZ8hXIAqdff
Y4ZQ3so/YTreINNnLmYe1AnG9Aaqv6EDJSxzDNQdC1tR6SxKUWlcAUKA67LbmIcoaQVKsiH3QS04
mpFon7k0TOOxFmwarc/pTw4Gtie2BVElJXOzjvlTDyMqu+YIo71VD1m3aTe7do4+VIxMLTmVJ1fc
ac7N//MIz7HbJlDJJBXy9D039TfQ2/9B+nhqtRFuJupnK7Mr4vbA0L7lrS+56DafaOgU6kMDuGxn
gNPfSwn9LrmXxdyOhD56UsW8TtSlusu+Nqaea2guJZExVcem+4luP71q504lTE+wYXmsK8yVrrSD
LnsI+i8nJSiuLkG5U1BxF5ol/FFfCKnzitM6b9MFVg1TQkKvjj942z87oYtk5ifh3RpEPauQJPNN
y2srCo8JHjAYb5GjovuMgy/5Gc2ImTrBtW6z4TSh+TNyl0seRViIccnosApy01cyxIxAUjPJAELE
aVSoVA8SS5nbbtO2vN54hH/qTMj0xmpD3Ftto6XZB4wAaSsFGauMeoEtN4R8utKwFbH5l+ViqDfE
9XVLcU6eWaCCcOGCoAjqbq/E8afDXp8QuHBzwfzBXwLDnKrgeFff+3ydhNpZvwUzT+sineL0F3er
Tol+jYOLCTgLW2Sh38ZrkXV+K+9+BsC1v6idQPDcYdgNOuMZXkF9u99vPlamqlsdABTjzIbVkP/q
D2G0z8nSq8V+CPjWJx5MmZnESISpNbsaoBnVuPdJBhIL87FtYXNudVbFTXibK2MdnpWmnzqq+c1x
NORECKSwnb0O6EQaPHuVX1LzsHznWfmjMMaVBIHvdFJV+sbzsUpUT1iXR3p5OLY3QKs1+fzjGqyw
TDPZLEN8RlJBaUGXJIMqbiSiheN+E8WpEqX11QMu+gZgwXkei/9Bz8eMPjkYnUmOYM+a4AKmoHqz
PirG5MSyotBpWe3A3pPDA9E70TjAmT3+7C1Q1i7I55yyPxiH8RN+ys4x63Wv6oP9vqtZJ7QkDCr8
DqsqhXaJsPkCNZu1nn7jJT/ilkn9tH9mVFODIqEWJY3ROiPuwkWRgvuaD7UPEhS2d0nEIHpAmnC/
7nWJXufMIGc6P2s0BCy4hoRRM3rbLW28tbPKImO0pm5dkomDf+JZB0Q3JYhPhS8iIsln3sTLWmoo
1Yrpg2wF9TE7DTXgBr66dz3qrTK8iAfkkWbuOCAmGHLPSwUVo83zxWCxDK6yTelERnKWQ072PvlR
Bqs7PdbeylqzqLKoyegegPyBjpPnlNty+1EGD7lHzJqmU2vgjH1CBUJQyR75pMJkIyxE5w26sCi4
1m79xqpRemAGzRCpLHvIxsEXDmqgDJclr4X0o0t707g/fZ/hPoXz+GWQQ2Q3d2msij46sX8Qu8bR
ZwbLZeAJbIqUHhNAhpdYgYH35hKkWUjeUCB7rdltuhjmAJveWgo2y4Wvulakavb1MXvhIzI8hORp
Q/zUd8V7kfOLbwa4f0ej1W2sWFaP0AM0BG5U3jatgpINORQpCGLrvXXQ8z/bbgL1FnN9JtLDQnnj
eeKzqG9xS9iZjhDW2ZbjtsHc09GWVmw0HDAc3G8LLndbGMH3+61zekGkvxX/fdlThNSSXpQ52k0g
Xers05PrfOLdlxu7+d01VF2OuOSwBqlgLrjxu6azQN9dUweR4QwfWVqJvosvDQWv/uzicxf/tk20
Xc9/tBbFtonX0s+e3nsLrYo4ih2LBG++jFawsHu/N8QofWT1N/ZefLAZ1c2FMb0tacPCBWPKKyw/
Hea8tUD7XIVPiV8WyiyvRqAJ3oHYjOwgvjOwOKGkhgUwKwdI+cD8D7QPDSH5idJ/InCFiRpSZU6J
UrCknGICEEYK7/1GD4aV36xqItwaFZtSBStnwnUWPxNb0y6m5wi/2dUJAGc1rP189t0dR9MDIIsD
9I1i/RqoRnFXEDRphLhqJ+TXrvdXg1esgp0W4mkt+23tH+8fgT+hSexslEkzu6DwDo7dGjwgnBgk
3MremE+pfLcdq6Hrv3bzip+6V0oYUwK4Q7wLqP8dc3vCMpCdHsu83HDuIVKV4xZCk9UrOWUdkEA7
fL/CSC18JIw07u5vocvQaeUO5iiSwiWvAPbLhh5zzS/8Suxt8rZpnRK++fDQF595On7ALX94/MnC
N1KEgT3BeLYrKRbxsBcyukoNTFDwIhyxreyrI0I9ou7WQ2FM4orVSxJDUhhWCcaghnHNN5TPLExC
KgjGjWnNJRPkGNORobl3seo1np1scSBthu3GqqIzYOGBfYM0vYlRajKKf1NQB2ff37XpjfFf5/1F
MV9HJl4u8AuMzyAS41qkYu/YK9gP6qz29gSOmZwi+TWr+XgHb50Jghyd7pvpn8RvDqV5OO46P72J
CeiSW1ijuL8/9G/K9aB01N75n7KXc4P6AJWNTqjIWBLo26rJ0ncDX1q3oRkZ2FkR2OBGK48f6PQS
waFuiB2lMO/JQC0pZWzg2jpITsb0vQ4EZAx7soWxe0qflMBhb4uHBsU/ptFpwYsmu12MVcFES95u
s58SOUhdxgdore4x3DOKImA+05+FAXZ0XPIM5CF0TzAJ2gROI5GCGKmcGUNcAXx8+LlpkyckeUqo
X0nWXLCdJYqEM2UVKMSGYqk+w4bOaa+zQvSbbyPhqDJLIDziYufCXKlhAAjipqr2EdWDddiYytlB
8vVJRaez5SnerHWUl09kp6zA/OkjAJ+F1q/aRfBmzaRCGx0Jif9ltzNgcWEjJc8meBZkMhbhiSG6
9JYgJWKGhLU74jGEtHgHgOJ4DuHeyUIu6uexFJc6ePiBtu/QAcL0/CqyoRvCdI0rR2cV4Py2G6/N
AaKUrvczPb3z7CQAzYbFv/MGEdu4G9rOxDgcU6ucT/zjWoNM71iazdhu5I6TMEOuTggGmkusrmz7
jq5eJJWBGD8FSTiVq0rILHWKRELCWhJ6hu4VRC/8rei+O4qepfYkUFRtSmmTb0Fn2NT6J9HQOc3z
LeFpkkOJPZqqX3bCkSifE+dXouMruA4wpM9dTGUi7WklGAYhVDpXR58PgY0RtqeP5CcC06ZXfDEw
KdXUDP4I8Q3iASz6NgBfgrKV9+3PdQug+v9iKzeaKItzoOkA9rfd86/dr8RX5fmHMo7uAPZWwEy/
K9oBOHwTwVYdi7jt6BAQSy7Hya1fmLk8oA4+0UwvXo2TXfJsTSjG4KGIUJYX0SSNQ/oLKY5E0vtk
85JHc7kpuQRlHLUfPze8VApXIUX/KKDgj2/luPqCawyuGAPtJNQqW4VHccnRsON13b5iph1IgGeu
KR6kjWbZQnlaUYvLq9RVdDEpgzbEL7CKEbv+nQW2h4sI2yR5F/jo4AQPF65O2LAzv503XuuvZ7R9
DoTJXIpDb4r4h33k9y1RBO1DwWrhFbwsAJBxymP03MfIv2hl+gV4BnWWDpFhAv7GGzSLH4iw+hGA
lwaQZm95xXOtgIWTWlVJWSbjHYvZfqGA7rat4DgKPC7vLcwg8kaD0t+CfZ8GPTGx0kBhNtqYy9GA
POWMMOcLQ/sOkQL/iTfzKa7OfsbPIYMeALEnBJ8X9UvtRnmwgGACJnVAKQRyaN8t9O/9ZGlAHgyZ
55+bXsyhmZdpzHwYNj672OEit2/DmwfBImGrpItu6HgzRztyqL+RxI5zyvV4Mkpzpg4mnVMwO2/I
aRH3M/7B/XOYaogiymN4K8nDTxJDOOl0veAKlNLK2cd1nxMmnsT/ecRGbMYO04typDQ1uDq8RF6l
B7wW2Q3chyvDa99oPlwKtWT+WGJDsCfMnF2KHRaLWUcswio3Vc180rawDoVPNoDLTcaIQQIFvHyy
fdCQ4bWO794eNNoHUr5Pdfw3MRuWAYJhDchP4oVOFvOP/W5ezZbZ4nGM1O0XPcfXQOUd1MtnPBL0
NlaoI5KOCMLfbk5LanIwTjAJmpC3027Bv3Sqt0Ujt29UcIwx3uuvzEzTItA3XTZdbPgB1eEhAcOw
lygDnqN7I1ilDmiYekL+xQ7Xl2CUu3PoAXdLz3x+LuihOmcktAyM/tGy2YqDJbJVqNRzhBGKLVB0
gF+TkcXXJmcun268ZMkR9bMkwLwF5kxP1fwGb02LXWcvdI3eSpdznwNQcfbBHDGpTi4IYtwKm7hp
cVnJPQbiCVC/k7VLPNAOa1qzI5NpPpmSHr9d1OVNj7Ce3NxYUi0rMb+SDnqeLT4Pu0noqDuCCqXZ
77b6FWW/IZD37nHpPVNSFraYy1/qnT5iw+g7NajbOKtce0hnMxMHuyHQ6w8wTOOSss3y3sV13rYa
SQKjN9FXZtoJxoyaKa8BygC+9oFN603ZegC48S1IuausT7/1erYc8ollei/y3IEuaJFTPpDnT///
2WRhtq9E2ilUN0Xl1TDCLYypHdsA5HEKzggCKiIaaBhnmcV/5Klj/5kGmkafXntN1uBT6s+OtS1j
eBrm5i0AnTgJaD+ic5CnE0sfp3BIilADcOoUN24wnVI1A2az6RYfdMcORGGbDH9g+Cyn3hY3Yvuc
Tp7YdtlabFUXb94eUkE4BgJTkwqNexMTfJHaSNZbgXkl3oPfgzAmL1MR8sbE7MYe1N92P5LyZ8rc
P7ldUrOKSaMDLp1YqCQxcrcP4F8/r9Hldrc+o4fFAvngVvizB92rzAqyc6hONgk6S+51eXhnlQUw
+7XD/r6eN1UFFKei6F6Qs3KTXJ1+vIKswmWIS/PCCmfC3fnf2ZZNU4+aw5ROz7EZ9ZzMzab065Xq
EpMMIxMddj0pqUM+B2sLVMFlv18LBUlUcv0ao0UATItCuXGvHTC0Uu2Vx84TehZqm4tRbgtAKny2
u6y3dJo8tzrx2IoqfDiPZBHlS30PRKJFocdDWdQPXxkee1DTf1hlT2NjtpXRx4Li6JwvcpnhhgBq
err6OyiRiec5OzdRQFxMSdOHyVUWfeh6jIjHBNDOG81qoQsf4BkBgtT2uVyflrQxaIf8rdf90iS1
b3SKee6vqLEWfar/xSJTrlf3tFez/I1vdzopQZRY6C0mQvF0ZbyEv0e+ddsbLaZjHlchPmy5DWn8
b191m3jH5+nOkBN85oXAW6aG/a55ujaAZbzTe7yCSe33eTC2oECpau4KDL6/mLljbo+0qyiTxAfV
o/JUQ2xMgRdrlNdk2qVdFbWbb4+MDr6INfVpE/bExhlXax3eXqdVYO4yfLhGRnc+3+ecVfSR1Vgg
u9KUtNYabenbe5eWMTCeoaME+rNv8HArhHRefcnk4tqp75nPNvmvkcj9t8oKgA6ark8kg1KT/Zbt
UOuc6b7H4Rk1IUU1vTYiCSdwM1sjRmQ/wOvlTtnbF5NSuGDOi5pScm8J8udfLR2K/UYOc4q9RX8M
7cz55zMAV/89wslWvXAt54xYUT49keqNsx6ZLiherwZIgPidxLJZoiPFU5KRYIntfOVFCB04ZIkr
SUGBmKy3RXjqaJwG6jsbNNYceX+91BmPBtXG7+hIhCkaWmKQ/U+41hPL+g8EWTG77td0eye8B6eF
K/ani6aEyNWNMXPIkPxCSmGKf+xGUlt5pvMBMF7iyEH1E5i2fYX8aenVmpFQr5K6abxKpNmgla05
6ea9v/9rutSGHwQrtZw831obrEdQ0foTXU2Ofyjsu2bIfln/qspe826nORmClvJn3PhIq0PxaGSQ
U+HycI+rBmsgUJrKGI6G+LYcoCOKF7YT2MjrNdIs6NJuVkZSqbXXRQfMNQCWGoOtGKKPFG9xZJzW
E8OTUnX1E+HkTmQLbp4KWdQLKv5LbJtCdskYaJZ5hdl6OTR28MDpASprx0LBYP4thG/KJeSnCZ04
8gCvJNMh8luNXTLKDVmnaoyJw+KXB2u+BVZITSBUoAsA2d6LyDRocTiok5X7RuD4gP2HB0UdJiQV
rkttaFWwTfQUAE8S9Y4UQKV81A45e9miZ+VuQYbd+yyzZAEwRNuh6+w5BLcuOkQo3O6k7GWzRavH
uzwhH8rAErlDI6MvNfK2umn7gFzwlwcEBhGewSas6pOJzPEAz1pLIP0Am3pD3tnCpT9p+H6wlXA/
hUUXwhfRxBHxAPPh3wVIl04Fx5a3VkTd+Lkt76TimocpnH8o4ezhLfclftoCspOyv5iS41UhRPlN
f1Xn0wvyw3WuLMQ20+CklLZQt4wuJXBeLN6ahEy7ctY3ADctc8d4ax6G+uJAm2ACNbMn/ZusIcWa
Ub3CjM/1HZBNHhj6BIIKwKUSfNzVo+Rb04BL7iwO0q6HIun6QreDepUiHxUFZBMLXc3rcqOozfkW
NSi1Q/HnKtIbGGUVtrpa0h0NYZ+yMkPWS6dXFi4d6iP1sp6h5D35dYLmnHRWz82GHZBxMosFVoox
TN/8Qj7ASN0jDHAiWyN2bVFWby6WzzT8QWZ3AcSiKvETmHKYqLinc1VW4ApmiHZf5K2abmc4y5tn
ZhLuo7xI0NgwyUygoi2zgUaPib6my4vOP/WrqfJ8RnSSkg8FZ0DpVdOodM5lpOnZns6vZJqDyMVV
/x0hgWBPtezSRTNwWu/UEaPcrv+8H4/97liemIZzh7YXHd7SK/KqUVIglVSatJx5SufdJFtYJ1pv
MmATcHmPcJJjcF7YyNSruwyECNTSsskuVzXgHEDreM1ZcaONdlrqsfQA/OLD9MuT2CqN/4a8jTtJ
stTU7V1tZCxJR8lQ6h+uUjiV806JbNpwmmK2awJm4hjW2ZoAY7+CSKTUxbfJsQjrZ/z9yOJaBbDO
t6KN1KpOUayUB1QhPkUR5a6e27JlC6mp8kcD50E+UsLYGISswYbkydGSMB1jgiFl4gowVCbPkaoe
S2fQb8JFfUPI7HsuPWBFybj20a6qd6FxRi4c6gSLxiVPt6eFFIZM7L8XoiWzR0/SlxuMLonz78S5
7PcNxdKVpJF2VZ0HILbzcfK/1FwFQjVTSyq7xWdFIAHTUq5jGf0Y+h9vNsUy+qK2TkJtfBDUuORr
kfF2R/IJj3+vcoS3oBNV3sxl0HMvzMLYTbWCBAJFGCLrinOk9Boe8DtoA7ClP7CC/d0LHid9Gl8j
YS5b01mRwgPZKWCghToavcb5TuOiuIS6iam/dkv4OiEBDekQBw+umcv+hYtezgAojscKy9m77rtv
M6G6jHgNrWIWuZbI5yJb8dG/4cTu9FS3QsstPjbx2Chcs5EpNjNDv5DtPzcfPv7sJs7BVXfOnEaN
dZzrdCeycoOfQFfAX3Tm7mQef7lJ0hsGW5Dup5MqbQ33TONBTUpBa+goHDAumTS1vM4lnrF+bz1l
Aj1BxhPUid8P8SjQxBRIiflo0d8RPVLErSk1sxCmUDSRL5c+lHg9lbAv2tqHRp76+oHFSmeXJB/A
qs9Nnrj7UDgZqyGHJBThAfZZ02PEJZyjoRbez+B2ew9vHArPOX+5PpxhAeRDasMpwq9ZkM3omX/6
IfKRLjeoxquXgIdQ5bjnwB4xK5058Gsz2RzKatEQ4V/D6POD2AdDBhivPtN92wuO+BbeU2GQfOXY
URhFUDW9gd1tNnP+0jW7RaCxM5ROWUgtIHZdiXrTE/oiXb7Nt+n3oBKUM+FQrHVJAcXjEbsv2LIN
noZznnLJfOCxhkaDN2q3M+adMttMcvzKibjKl6LrKCU9vMViGR77dF+QrRuwMB/JlXF2R0V2tX+Z
sMEXbCnOqrLP36PkuL/Ct4toCWmNyeh9ad7Y3BNKu2ZKT3gJZtmoDnUc6YVeN8ZMax+l9MrGOb7c
twMg0Q/1gczRmyeHUQyuPksGSUOJbdlnq/NhZAS4s72sH4ZtEVvd2T2A7rwSxMLyDvKUU70Hz8dw
NxUM6nxnu84tse0itvqqPhru6pWV7T7OLt2cwQ9uG/x67A6KbPsh7sF/nrfLkxFoqnN4KIbj6P48
X7/OwiCBd0+df0izUn6ltTEjugAETcHFppENAWBlqjKlV9/yORl73h+gZuSedYazhY/VufDWaEby
ieHG9qnTrPvgvZ3HtmcJniTIID2fpe/CItO0h0vNJu+MVnih/HzLzcDmhlqAlKGyujzQGzWOpgX2
c34iQQgyj6aoRnyc1NKL0yTg4BB32EZlnL+uem0gx24/RMVLumjpR6K23LLrzi0W+ojSwLUPlsIn
XNkgYJPKlGG4QZqAB0i++pLe3Vo+NzaRmmlO9KAeARFkOLbGhlNJQ2g4Yz5+rdZ1LfAYdfm+1jka
VggIUL5UDSdOW9pzHz+UucwYPCH5vgzMkpow1DMwi5CWVMVr1CHewSdwnSE/QpfQL8DhzBhmKQam
9EIxtwPnu/+ECiqO/7IRxN3m9AgKb6pcYRBVWQomctF4eB5K8FEqP2T/vdq7afGgqfos/k4zNygA
qWc+2JTmasU1iS6ekmsm7DCDTxBjnnpW4NXvCNsETEZgG5ZwNsWJv5Y+HxLuUkkff7SALGbXWgBz
NW+6jNZSk5VaV8SEL+ofAJ+tOIgZOaSMyyBNgrOQGfz9uFQuspxLu3bW3WGz2CdtbYdVh3Kz+sYS
zNlAdPKtvom1vs8/BnGLg2fHRxFEcN3x39boE9IA86wDEdrh0ZtXHNIkk4lFHxrP0u7IDfGWDNOy
3IXOcJbbbRblCK8LTb2MjAYVyOy9NBU5jQM2ebeTF3G8YTW2JWUbGSFQPjVYI2XgXIjBZS/Qo9o2
n2nShAJnyP7wbchLqYXGvvSz721BQhMse1gGcxqALPBGpvTx4F7Az9ykxyNkI3OT7d6mvOKI7f8e
d7VafGddQh5PCvFps6bMV/arIK0HI2p18S+fZEFSLzqFePD43pp8bpVQvugu9VI4VrQU8zfRIdNA
Vcol+kDfLmVy162fdqRPCp3FKhs5WqDf07shagOIzEsogcdbB0dGtNSv3EIxpmfyn4ojr4X8B7fl
h6SYvA2o6LItz0nbOq0dZA11ZVYWRBjUpcE04OXstQu8ZvCPgKJNToApDVA3dtX2LUckCONiy1KI
zKGntJqGuRL4xKfWv07rRGDPMCn0+xxLWqRdengZRJPjLkHBmVtgTh7KqsRXPiHYPcoeY9qPoWa9
0iLzDy70q8/MEKbWSnj2dxa/laNRK3Ewy8peJ/NvhztY1RJMVWRSrq1uzmdB5udTvFv5+1UUzLji
AZnf6+sPWePveDkHGQC50GL5h18jChbvdsn/Ldh6ylgPrpLpW346eRhREWLwwzKIrVb9p+O9GYsP
mp21Asrj5BTyabbBvFO01C3ufObC8NNMy4IOQsgd+IPUeAYoqzTuDovmDe7oRzBrqp/bU8//MK7N
unj5jkuWmyc1tZu4Oiw06QgcZwZMepPY3F3nboJ0/9dVWvuvv6wBiJBG9vlIBhvBp1zTKMOM37cP
8jfazZkO3DSUyUiRQo94BKeYSG9yNHMuPz/zOC4ogNd6jP4LYhVGq5UZhvP96wNRGptco0rV0obU
Jig3ZtO77DbcNAwzGzrPy0IdKmSX+bJFbNP0/AIuqE65Frbu3R8OT0ijrZb8mKcREUWQKb24rLXD
zVnw4Rm0cAe0W1GBi+NUiIq5dMtVQRDETV49A+OgaUNCcLfFg75VqqLYCfX6KwV8jGYOtYcdrpUA
sx254XwNcl5jpDEp0U0F2PTADGMpWNLXwzm3wThfSwKASwoj7+/CM1JFBnBV4f/w6pVlM1tp+ViY
uqM8IEoq3U+eT3nP6uitgTOtehkjRSZwdlB+wqqcCAlJgc+XRy0Uh+0J+qqYrBPSaJakt9+1BH5c
hj+JWtMKN0AztV8m458R65XgqM+LY1KWhOcMBnn+gKbhP7WD9y5+5SGZL5t6OS6D9SFTW4JWI1Ds
zfbGyu4V/SzPVGkbPEGKS4UP0fy1moR+Vp9BgLY0fSHhufztQUs9zt3RH8eTqjCF8IeRVktqbjjK
JTxKzvhTRzKRq0H8v+GBz5sbkYwbL5ukjFPwDNKS6skSn0Ldl3nsg92GjDCY7nT+nH7okWw0RH+n
6iQJwI35aII4NOVMnm7PCIornE9Nl3j9VDXqxL46bUQKBeKnQp/2MaTrM01WbwgOZMNY7ugnvca3
CBVTb1XTRBYS+4KkGk+uqQA0PMU3+UgvB6dnOZ3cwKRGp8JKkYnSC2QpYMZ4aZ5yh0OsSCvIQh0i
OzubDpEeWweD+7TIZeei6hDpLx/sk7XYFLw7t0fRkE1/lge2fLjtmvI+niKJLDASowuu/RN/xB/Q
3G0uZj3QgHxz5OUadSrl1pmpdHRP8Cp4iEXPiEVNRX4SJICUtyKKZ0bXAMEEb3CIQIz8LwvaSF94
EH1VNvxn8YVuUPGL3bqfYIdKCOHEncXvbe+sK/4JofV7E2GwAF9Vi+OGbHgpgi0+FTzg5bWgLMSW
0RSNjNHqUH8/S5S1TZSxmpkgvd4/7POsRHWSgjnVvSQGUSen9DkDGVP3lUMmZRXBEjAHycQJTnsG
46RvOMhptUs9uDOpEqYHjXdWomHrMpBnME2vG9iDNye1aO/aMPZQFoDw6RywwUHkbovKrmSGy/h1
CsGocPXv6DyHpEoifnMi87pDdzPpZms12x8Qq2bkzk91w8yPI6saM3T7U4DhPS/Sa6gpYbnjKVr0
TZpH9UBPP8TJC1AHoJEthjASXVCRd0qhwEWJkvCsD6ltvc0APONg0DoeRzRG/hF3VcEOmwwbWgBw
LGPN5ImLuSLKsEcPNobH1QHjP6NgystrAkgIOQCEAylbjpkaGPHR/Bs34/RswFGih51oJ705ZlT2
89cvcxLl3QYU9xU/LR//h5JhvGuBozSp39L3I91r0ffeOLbihZKo63GqRWQ/UfYS84M+sHe29zqs
//WFReqrf5L8kQtTiDof9cLnEaWAxsogXblN/l9uoCIsA2h3jEDyOuSRSf6Wn90Rb9Yn27ya8tEb
Nri2BEkDmgNfyAEqwcRNhz4kZrOjzOwuzttG5WBcUaSMVKfBOnFV6y7Nf3tQnE56YR+YDkPKhHii
FZl3zHlSe708OUS70Y02kKSGgyUEV/kbcjd1QsSkGSz1WaPR9/XVQoeJlKY5V/YgZneDVDq2Lv0e
RIctnJKC71XI7zgC3xFBjIG0YD45yYoRthl3m9XjJnpwxKkgBYDXazIbjgSArPGlL1Om8X/KMNd/
/wC0DpZYl7FWi3l3QZj/8l9axsGcqeESjNY0okJ06RpAV7Ic9QcDnK3UtlaXo++7YOs3VuvAZM1W
Z5iqE5AT9qb9KUoK7JfDPlsgF1S1q4BKTeVwvs1pHHexHeS9h6YwFzefl2jb8rMuIH+mnkUa2Z7o
xeW2tz8SvUVEwd+CsAwhoUq6yPDEw9xXLDCsEGs/znG83vHk1e3Frsl4QsDZtpQ57Do1C60To+kD
7SzPmhKJ23EyCb/iPAE5W1bb6TmL3RfN2bIS8axL8jDj5ixLW9vB1bWvOKPuLfBQuUgzLfmbf8JC
31NHEuGJ+GxJEle+47M+MdJFJc8xzQIVtDvsHLxjToOeBSMTMRmqwNVL/AMpbOg0QIPGVhFlYAIr
dYIg/su4S3z2fiYJ38Fq3QdalkpTiZ4oFgXYXW/d8/2fHDtwWMIuO4P5uwOuE9+FihiDKV2M3c4H
TMO0fvMofuJSa+4wQt68aljCYaAiFumuNmWU7FHaVq4gl14/0j23/Y2CWUdFtLHnEJLZHV48FJFo
xHxGFOBR6r4ODQbh44/RfrNnBdSRwdZeG9SRXvCRNN0Q/GZ3nOfFOnCNf4bRlstxRuIadHjsw070
2v+2dZe1P8FO5VR/czSo2b1uLsVp9rIUB8oj88Iq95anAeqgFXVmjnowjwVQ3YV5BWupV59mEbcx
4sgnq/tThaXYKHIfs5ZyzmletgV3tMsgIvNfQiksNr/LiuR5kBxY6vdPufjM3t40yJcv5QsV20uK
tr611+YDbU6S0u14sjSduosEwqjiPKgWjy/3yzkZinUzVJe04HB1oa4H5yiy/KPzvJMd8KE15u43
2xkcZPdxrTyCfLv3HELEoEpxs6vxoTW7BO0Olf04C3rfcDob3uNs05ZpzFJApjoF+fJaWg8S6O5s
WHsF/9PjH/Szhw4b/phwrR9obCuwouL+tDTqQ5yhkDNQe1bI00bSHwQILr9c21gSnu1z1qeRxJ2S
WRLU2dr0HNoFIzYZKSjvHZfPng4ajkrLJ4GAscIN8alMN6nu6p+IYpgUbzl1TWrMUHDewBZnBfpa
dvhWHE6o+VFEIK+XWs/mAas71YpDtnk4nTb4gctJUujNBCINabx80GWgCwwGOa/isCmcT9VSVNmO
5VUAqyUsbTsWMdpo2btp3ZGnxppVDA3JKX+/A2u+5DjL9GXxayqrzWAg/DkImAiEjTwwqV5oTIG/
M4sOPOM/k6vkKH67stvs1wHqZvm0GPLln+F0RloS/9BKJJXE1+cS1KTtt9eQUfIu/gF6IWeJOwSO
JbMg/IWBryXa+djAy84v1OUmJFY2RgX87ppzJQl6KiK8rkqFP3Rs9rVz4C2Wffi5dQvD4TshRfsY
GwlbSI9Vi5OhKqee4aYRTgXtbfyOF3Mwts64+kzsODJfx7KJszBgbu3KnPOiey/rdRlvW1z34yLW
xcRlQmGZVJaskTCMO0ItaQn5Wqk4HbUFWDs4LDQme/jF8pqdGPGgc5HbgpiYu5jPbZ1KJXNhtUtB
ijzzsYjqgMv3s3WODv6yt1m9oVGTwx6TNVSNK3Pe9kllwFCeBNehXfuOOoTEgJlyLleWCsxPoBZD
rwp+SUSv0tOkYKBpt+l1bKDhxT3S7AD63tJjBJzZjllZlPRnyyNauReNCS/nVZ/RQRGo++QAcBDz
3jps2TFZ+N4FYfRYMFNHJ73B2erW8IWnZRCPjAN7GmmJvVbAETtvclsnN14VD83IdMe9Ual8AiEp
+KvoQwkqNKVP42aPwbatlthU1u8QtCPz+6p5cRNKdRC8icVE57iqHITad9fMQDCYWGUZFC0UgX7c
ykWeX5SqB0+N4U8cIZl+F+oeseNZWaFoYBt2ZWUh0mYZWbBkY8jr3NB1J0eOvJTNzZxQnvfNg+bD
39N6AT+yPiDoPN+Cu/YiShwO1f4OZlGsjg1dS25NXqNph3YiWdmzu/QP8CBeulZRNPlPrQRz16rA
oEwNcKk7zKvmxbXqU/v8PMIlfMaFr+oBhFNYJETrVAmJ/4kl8JCUJg+O9TxjOsGscTE6l2gcllLc
OOs9yyvgOhSnk8uI0YC84o/eY6X31pTgi90doM/1utTe013vTatz7WL4E38zJQc80qGM7Y5F41G8
3hCsGCoKunefCcI4HjFIm1ivgadAVg7z6iWQHjtgIN6DZiZlSQK8tDi4cv5lo2qDFyrgJ1KWAKcP
XssC1JeKl222Yq0NusulIlqo6K+4A4b4iBW4g/uoLunEmnu/1h+XkPKjFN7eQ4N6bfceqjPum/l0
TqD8wZpuOC94hY3E+oArFHVWRq/4yM4YdufVsiciakWwdNb5tDa9n/46YQCxTuGH+P80cOcwgb4p
3nkg0AbR2u7v7FIfRy6vLKcc452N7R5KrxBn0fOJWvD2pmud10f9F9ak5A3+AQtfPZ7Zy6uBRJ1R
Dzri4e4lDpQr2E560CWx6IUeE0OVTIr6IbOhRaTOPE2PzhJKRflDeu1ETUmfnIYzoKjq4L3UorSs
tbvGee7HiPt9Cw0TssXP/Q5x2nwr+W0IpaecamzaEbN5sBj708ps8R1JrKP515bcJEB0K9zQCcc+
noAEHmqgxJHUBmDVG9FLsAbclHEURj6SXTGZoZCo8LHoUy2S78tm8MnWqt5VcJJEMRT2+xKcVQ+S
cdiP5AlZ9M2ZGWStXXmXCL+0h4aQxJqJbusDMolurT/h9tupQt1lyHIKUmFXQiYYxwi8PqUlOaDa
+MFiMSd1F6kAOJrL/GW7fkUQ+9kY19i+XrO/GSgMSLywMg2lgWwrUWIPd+5/yscRr6t+MHGIWTY2
ZPN5fDu1lFWmAhPStEzAqYIcBWqSUzsmbYuT1yNuLZPLDefAVSDv7Qc/GwPfCAc8GGWtCLsuTQ9o
wLys86a7qfeNVHYBKN8vzXFjjuaKtJwa69c2jQVrlnf2HRonLicycfMpmVioxaXo01VSMtwobV1c
uwa7Ea1eSxU7ZOwUJYuzdzUaLBO8doPF558vmbe8nMQVayVKPID4O6rLS7XFtj+BH1H1tPIzrArD
1d9g0EuIGMkeQzDftCnuVtSW2YJnknQ8Zo9+Pjlbgf//nE0R3Ai46C2N9Ff+iNAf1EBAPDNMLGT8
juyom1BXXk8TpiT9Dlv+kTiS0htiQdb9SDECAkI8zcj/K24rg0PbO1Jj743gjiqLI/1z418+6a0Q
UhVlJAyGzH7R2DZ5OT5Js2SC0DxSWBciZNf2aDQXVUWeDxPrxk4iIccCiqoVE9KtdHl5MDqjHaHE
DQGH9MxMPsMH/tYGR6BXhvszI/ToBRL6gNpu8sUyeqbrlO7JDwL+rK9/GPIL+ay/A+ESgfUEKoNw
r2PMBDas6B6aBHPkWRXJdqZwg+Vu5aNbHFnIv99moUgHpa+BHzMOJjZiq0/1gBDDB7/HRN+qkhv1
B4jw5Be8PHDUQGiT4uCZinoh/BdeXGJsuTDoGpndpDtFGPvwrxiFALdcwl3139gdJnsoMmH2JNTr
pOucm2PJzqNkDNEp0IyizNRLn2A3/Zyz1M9aDurmFALmkDLWJcM+KDEgB5R1tNs3GzuOvYwPfvvs
P/d7U7wGgG+h64LMRfAbtRr1W7Ohz/SC//wd2nlarhXzOc//Lr7DNx4EybtJh12BD/aXtVO3zGeL
FbmejTkSGebaa8pc5xrhEZ2+TfpxMQrz9D+8mhM+mLpe6FcH9qWDooEZyT3j2ysfXslgq6uM8BFP
A+erFoUp6kbSkJ3/5/fDOzUYBEUXtAZSZaPkkA0vVRoqAAfSZxyuKUfUA/CXJwpUmtyaxyFdvx2r
LpFY15bLed1fV3m5FWuQNiKM9kr6mpnd3jLcGFpv7rIuurNydG6fsW+kdZIBnJqHCerWjRCGiCAX
zUOjeMxgbBIYSEBHzFqB0y++z+fyTCF+RXn2L+kl/TxV15n8OF3CuQjHqVcPnPR7q6z7DH6GfuIP
1nl5HGyqCFfsvXdKJleKE/8ljRHNZB1TaZIDBuY1nLoXcOxu9gZfMzve4YzDoSRtPkuaL4x/Tz0O
jhoid9v9JDbIm8szlr7GCGFjOmlq+sX7UDO4b08LDyuUnaoTDi1bhuQvtBfJs3KmW9elPXs5syOn
PdEOEMx8qs7Gr9q2b5YMBKLn3R1zabM3DqND3caSoMqm4FJy2ooVotbwHgP/PkfGGyRTjJ1Sszub
iWi265XZvcgGsA1U4uLxCXTCCvf2tFEpJcfIbHfyZZ1HSUe0uVx9DguzxVFJxrkf0LYuICKqfrdO
3pvmttanC3F12pkB0OdOWFnRMLLtqR9Fr/4eYCM+/SKKs+DRgEGHk/YFIGUoz2CZAs6iaZ5F0GQ4
6qP+gAE3ZtrEDil6e9hW/hhN1fK4LSn3ASSgw9Jj5RdHeRijJeOIQXFRKeHzP9I8ibXiL69S0ivz
DKi21TaEl6WuVVMF1F/ztEgC9q7dvLiG7Rh5Rls21l3QTIdaJrtFejJM5w1oY6MzIde5hVg1lREb
JeaGFr+R/QU0nlMIIMRKb1PKOijhdtMOjC3OgxGBT/8aHTdUgfxkeIEe0aP5hUzrVMWkx8wyYngr
uGtt0gbzgVnmcQV2Zje3DkDSjyXvZVuLKDbn4MuSEmN9l0BPYCE+uMAnUq+mhLleH5SRL49eF0xx
FOUpN+a4wAWIcMxrYMEPn/g5L5eXd1cX/4i9E23pnaRYv+7IXAmg7ga8o+pjeKwNwMmXtQFgOWIE
MDSKJYpHkJawFj/vg6SHIywgUFPGLFVf+KaAKb+3ZE2PDxAwrP5jEY5aXbSb91sTRE3yJ8YVDgZx
G25qUSOOGT4IuCelDfNxDFI+AVIo0eWDe9ETm0jxy9+Un1KGKgkaV5ZWJroVSvRDosP+jfbkKGtN
7UEvf0Kmez8ZKXMKJD3lzGpn5e+/xML6kqqObohASQVILdRghrgdsavle9FvsuHc++ZBOzyUkzwC
5kH8+Je2M3Ut6/tHynvsng9y8o+cY06bObTFVFkhxvHrelMImtkj2194PtPc7yukYsmPPLcDmK4S
dn6f+3jA4BiS7PMdRekSslquHGIHpT7Et1ivXsE3hz0YmoaCxCNDdhmm6Z2dnCISt8hkeR6nHxVo
EFat820uRnPE/FpmEVk0AJbm2FeAAqRzBGykxxKVBPOhQVOezLno2Opgt7GfB/gY5NvUoDYYFE1y
p549AATJNrQ9KbDi6lBS/Dmwh09Zy4GYtyMw5siG2QY3zPo0f8uxLO3nNKFoufhuXkgg2jfWSAL1
7JQ0OqNH/Ao3SGmLuL2rF6NdTWM9TydZTWnV8j+Tzsq9/LTnZE9a2A2cbfkaEQMHkNdt0dLfAEti
NZZWjGvVpG3DkoCNGECBncbX0TGt0lQz/tiPsd6Rzfl3V3bN/Kc+6vVVlm8iK1bqjk6Yhi+ClrrV
VG7ydbTHdRKiW0NUURot73SB18j8qRja3FgEXmp56ZXhU9Kz8LLvHDXo3RxVQnkl9rrYSHf3ZwLH
Br//kMs/Y4Wkt9mgogC3ALK/SVLFbNuiHHSLlaD/3kMB4u6l9p7cWPIzSPD75ST6y6JhAJ3a9g3I
RLkRyVOR8ty6ibwqH+KkJr4SZO0P8AiJFS7n6M87MV5X+LuRLofZJwfBgt46qFvM5xREy3QF4fqb
bbw66qMnEGFGWP67QYJzZ9/bdAAoyZTboWMZE0m0VWwnIWL1ygMqRedTIkvblzIE1DdvKhql3J/a
iJX0MfgkSD6gGAUZ2ceEMLShde4GmfhJg9kJ2p6iPEq35by7jR/8qn9L/wbQXBzQy+Pt3SLSIKHF
UV8GhAg9EluDBW9XurP5zDEoc38RCPSGLQvSNjKCYT16/XyNaFQTLvW1rCxT6gtaYdHFSnD4xOen
S77CsQNbvvTY8C7l2BNl0V/C48D/eyRXg8Yw/ODQxOFos2n0IGnbMZW8jazA2CTLm/Ik8i1EOvXE
0wSOABLlnGs5Pm5nDrLIUBdTO9Z/v31cdJ1k7lq4FIZsiDr2LKd1UNhJh57UWNgRnj6WqM8ru8hX
afiS2bVGHVVnzU+9Vh7/3lFq430d4vVepG+A0UwLN8eM+QJMOn+SQZ5OKbz4cJmhC6DHRLjVUIPg
/lV+PXA3AnA4B10Wyjudunlcac31atCS73vwv2bxTS9uBsaGCuhDm21FZBxBsv6NTcd+grYN03Lm
+CrmrOn6rHIPPkSuMc66VyEbTx6o2/0Rj8rfkpIp4o8N/EgAZzq9TyJwS0PMKLLdZrl97lTSXVHs
FeI4XGhv+fXN4AtisRup2mNKq5odYz6TCW3kZaFH7Dx5lgPv78wTwzFD8odETxEk1/ZojHAGgAsE
SGyjf7t33SfcJ97jAUVUvm+6309fO+Te32N96CtR3KjWM2rFyAfUCUp/CrGS1DM06biUZGqYURBA
9O9GkLPz6Ea7eAGsrjl494JMSTD/MMjcU78/9jyzID+kPAik+QSE+CzvN2wMdtNwhRey2w73i4JB
7rumSEmW8Rr5YKBeTCh+IxZVe8001MLFs/h+pN/htt4hC2pQJjPeqdZh0J1rPZEh+7uYMqIhlL/P
SsEYG2brBysW9GMZhMC3YYxbEfw/KCoeULEHDquE/HT45AqYviIzLFG6T+yxddmDNtBRSyXxr/oR
GB6O0nbv8LsnjPlNjvaT6igp3xP+W6D9jd2Gs/0af/57y2r/fRqTIwg9VdahiAhO3XpampHFeLva
+6CpBERm9sPAlPcZ7gDcM+6bdXxqIC7T63a7WLHO2YV1dQanYcUqJYGzSQEsUX7yDLDMnegNky8A
pGSqus1A0glr4DQng0itmtkby2p8p3Q8mJ8b3wd1yt2odjxVKbnreSIAZFUaS1B/Gyfw7xfPlBbw
4pwrTicriNOFiW4z1kldwOpzJdZ2vJgM1rLXknwVbwLIgpx/VH3rCJjFqIVKvSOXrN/HCpECM+sW
1D+49Vbglxi8gZEVzMUmzKkoEJo9zDSehqs1/bV57EPbk3ngBR/FiHBFO+vE/GBKmGA5bibxEpb6
xF7VTlWLJZndBL/TrXjx6YWM30PK5QAFVTDCcKzKlDGGlJkfqzLCpXGAuelkZq8LQ44I/Wem74uF
eY/bBIaQWWKMHcbQG3c8ocmvBRqlIfsC8AnKfdv5sEUp+w6BSQe3fNC8ETii/1ahkINopnPY/DQv
3mc+/TpGier7bYddzJ6+GcihSDZGXB5rqf3sNFcsEmp4Mo76RlVvpLfpuLCOI+KQhIeENTCh1E0h
k0x+FNbqdrYbBtfq3r7DtmW4sbj1cm8WYIYbxzWY9zKwaL9zdR6iGuBvLHyDthsd6KX0NcF1tjnV
xVqO6q5WHLqQqkyRDUUNyjI+4RdA+zVeLawQXqJuh7Ps7W15fuiBELurpEWwraOdfSK/Fi6f9QhO
2UaYkXF/XMaP8TSkpNG311A26CFE+dEK+POiAxqxcx0q8RxD9Lxmm1Fr+c5gH4eKwAZM/Xo8OVVz
MfgwoROVro+L3ZalXsX2trAu+68L7muwRhs2teySOlDC0hgKQnIKbrEotQt/jIJochU88ZUxiJa2
B9GGGVQf9wQQNNhhiywEl4pB7c6DkeYIMKgaHfxJWv3PVn/4JMSRm9czS7qktgXr1+BUMmu2Da25
70lBelyppMSDjetuCtolMaPWoHcHBw2EvYYGj+y/Ecvgc10kgJQITDpNtTIaa16Rz4XfP5FzblQM
yK1yWaXKeRCm4NBU/k/qR7R79ZQXVCaiRIUSy4ToiE17Udq81M+NKr1cCrqDN3s5K+JmnWN7xe34
IGdffHUFG4bjVGwNyKFnuTWDXq9mu/7AjzmUI1cAIygXKOw1sLf4iVxtMcVNvyLNhO5efLC3cTWc
XG7aJdsvp3SFKFH2HU3j1r+7q0jbEab61nVRBbCsMsZYY1sJw7RkqvLo/EG1vK6+DHbUagK51pwV
NzHeJ4WpYAHTETGwiP4R0en/7WR1ledR453lM3lAxOiuTLOR5g8SzetaeaoLl5SJ7UUC5Qc0P4Ns
izk5tG7o4FjOnYNEljShCONMJJ5X5mPTAiXwh4dbmtHu1ZZaOX7N+vfHImI1RF0Ex7IL2xJpW+Cp
Cm8fmZWA8g5zOwVq7qOFU8ahhnJi1zC8+MER9A/UcFVjCT2OEch0j6h0cIUXsA6bkWUpL7jD6ROP
Mr8EdCuaYjdoRp50tPqQYKfY0v+aIT2glFX56SvnQ6l/f3JxIY1WgcBtbl2LCeKQlRuHC9pwEAW3
z8rIEOD3YgDAlSk9O9Rwc/a/tew1CM3yBLX2VAAK0qfQhRrkYrkHM+qUwfwmDvg5s5x5eOo8WZI5
BdQ2BN7mevaqs8Bm+WcrK/0GWQuh4JOqeOCjYY/rozdwtCAZwQ00LyQ8a6JBbeyg/8jubn5+uUtJ
9pgaAQAZvrOu1krMh2QsXIimnV8LJ2Cb7v3DUbCRIg3SzHiqTy0b6jjTGCCZnMp7LyzA/iR2H5kQ
GOQWNJhNf5FTgnJiZxHO7Ph71NQ4T6keU6E6Krr59r5SY2cID/3HOw3tT+G2XAtZNDsBb9ZQ5idZ
CwIVvXLSrFCjF5B4YTAdXO2J8H6gUCguOhrc1AFSiX9onPh69JnI315RGn/NmfpUIlZSRWg4KMYo
bS1uhVkX4mL/qW14laxkPRb3n+bNLdCQ0/UjSinqbLoGEEIpz6/MIJepvXeMeistefBPEh8iIZhL
X3el9/4mvyvjhP6cTDBqrT1cKez7pPN72ErNb3uTmtudVRb+PQAKVynS3FRRPEO679yirOt0TnVj
ZrNBJAdArMNoNJvxZF3KRS6S9QuV7DOXKvGjiK0vNMnJtps5f2dAWlNBngu5pETUeQgQPd4FCVnp
lPP46QapGI9fSr1bjw8MD3W8XbX5W1toEAL/dT8435O7l06uUpIJK8HFDQrVteSO4kVBVcHKzKfZ
witbAsqwe94Dk+PlE+I0In1souFa8MJ+GOfRsvhCcmjzsCFYbKS4bsAz1NqtBsORT94UO28VuZ22
nN7yUJBQ/qwOWS1UtRuEKp8tHRYOXKlmZhUZr9b7g5bfAVgTPHgRzzFKuT6oj3I3RhbL1EmCrGhM
FMPncNRGslbKtvhZFs9bBLR0/giAeIYiwZG1NLiEy7qbP5gpz2bZJlTBuxdQV4dd0aosKS3IDtT8
VXerGBDKzUdQESIGQkaI9fpuMEHChbDs1B9VrSq7TlSDepyGRkjCxP2edCUJDNkulRE8sJkb0Nm4
l5U2sOh4tF1WYWOey6oQp9iPlsfG7pUSi3Vk2auRG99xa5dLGPgWosVxP/7zN3QoVK63B5JshkgQ
L+ETmVO0Ei0e1QkHs15en2YhA2EZZzD2b/COW5517mqf3EyBObfXsbIof2PF+n/ooJZc4kqUhnoD
U1cDfEm8/tNfge6vTSae2DVhuDCw72gYQDuzosEGHMLqFBq4Nj/MtKtkrIxkvXJHWHQK3dwQ8BUE
/qIvsrbd7BSseMKoRMQmx5yzALntleOZstRVXXkxwT2h41AjCUpfz7xah5Ny77YtO7VXB31EOnWQ
0Q+giFZQJlywFzYmsSIdrd296h8gh99G+HZQY2QoSsOje6tbx2Fv5B859mOcP1hDwu+GZOBvR8/u
lsbPRI+4xl6XfB6o2TpIOSKJRtSTnZqSll8lVfoeeKj73dT9+sgqhJ1f5D4VAebtYxsgHyRTp8Q8
Ist5rPhIZ/a/7zBecqQvA1tiUHVc4I2ST8ftOuZTRLebZOZ473jwEkfemE7DceqKWUiCS8ivsVrJ
/Z6wsXQuSriUQRSG3Hf/BD2GPwKOv2zjW80jcQlK6InuZKS5H2Glxdz29NxhmGO0HJ/3TimazoRp
w35KzsF7nrPM8Y6nO2eTx2OtvjG+82xLuZzkxRuts0xj8b7+h92w55xJIL3U6z22K+PawqeMCTdE
P5vHrXfML3hFqPKL00jjt2IlxL7rWqGS4En0ro9gi9150A00FU8G7oE91r/4smy1pWu/D7EgAU3O
bGdv+4C4N/fQSqaxggYV0i1H4TK4n7CTYRIzWqwvpnfX3Cnm9ihXKOXdbhOV7JHix+gWjyfHnfVZ
62ulXuRhR8yMNzKoWuVIPhJbhj+y6nH4KV53AGRpboKL+S8d021aKugfYzb1BZkf6x4kNkmU4TVx
EWJ6mvodLuO5NiffgZJyz5dp7o8fka7Pigak18qERy0tmtLyyo9e6XmOxM089ujy2H+AVB1WZfPh
Gr9SEyr5v1hkLL0NM5yxSDsU5ndwr+Hids4WLkCVOTG8HmQrOb0rQmWI6DpAZ6Q6m3/t2X6c5gkF
M3QmbMZvdcP7fPo3XUVuJF1k/ZaWDVlWKSfCIoVX7gAenaqFbKjsMz0HPPBmr290mbb1peQ22N/1
hsMSgBKJtupuyicFZRw2lBw+IF3LRmCkI+BYf2Ooj3A+zQok6Z1isQ3iZRIYncrj7LwKvTycurG9
Yt8F9hJNHXfOBeAbUMlStYifLfMALrnu3fPKhom5ykASJGkk1BO9WzH5ALpXEVkvbj3fl+zUh74L
D6ncvhhvD4Fum0P9jGV1XNtBqwOhdBNuO7yGVzbao1AV8gbRZt7yIs/TlQl49/MUEY5mLQgaJ3lp
WiLyRftW7uarWyFZGNN/sMT5ogHO8g05W0vUdsZMwIALNt2K+zYKOsY4ffNlbCiGl9wgCqheJuBe
cDSJU9kQV2/XbBDEtqHpiZrA1gpBZL4MZJMRVb7Yt8ux2V4es4z1QL8Ku6PzHAh4rJWgxZ8yeIuk
dpV4YN1MTgxP5afRpdGAiGCeCNywa/SsxG1S5TQxKmHOvxsexlm/CTXxE3G8Pdg6qjgF5BC9S6YA
qT2cOI3MwxIX+zXDOCl4bGWgXKNI9fr/zDog3yK8bPIu6hqXdIQvPd/40Wk1eptI+PH5Dg6O9fxR
En0iv8vPEf3NM18bATZIg1sRTjvVTe5lJiBhkqICJynyAQ6ppcnxlRtpwX+63YcR4q0+IuWX1qwV
ggo21ghlkQR3+tDn2Oqw929v11sRuJzMh+DYDt+kU0HnadWQWzbn1Wa8eQCOwqX9GTsV8mxQSKyE
gCLiqipLCQJ3jh9msngAZG++oHvo34xL5oQz2G8Pro/HD55d79Y42D3BEwVo4ylt2fYc0g0h6kGU
UUjyOtHotCpvZrCqaMyNUMcC2qvG+zNdlP/o8ERUrmfG8DMM7KsBCXTGI18Wli2mb/lQus0sB7Qt
3vu6y70Vgn/JfuIcD5sPs0c7PgDizOfiwqaP/9oSrICSe7NNbCaKrYp/ENaxz9BcYOSe+Ep9pZXt
2aOsjV+AdHc+N8BNEx21Byks2AbOZjsnUL+mVsjFIVpjIu5nHl2R3S6cY/HwmpJvIzjzlhES4J7u
isdeYzTOZiPfEWE2esbcOYsA9txU3IZ+H+blhksFDVdBfuv4+nG9N28oSX/EbMoDJPzBtj0mmGgZ
9aW2mYoNx8wBxu+tAne+3nnGvyVWuvHVYcYBotuItxB1CshDDfVYR9nX7rIm/bfLLHBFBio6WOJj
e5uTNZWbbH0DtGrFg9XtJ+fsNDhv2wcPc3u97i51PMliO8MzIGNcK9yipBhtVHAy8otCJVZPWmEc
p70bNWSuI3mmiXUQmMJCakiRVNFu9iDcIUx9LKNQmixKeBmvJRR4uj0/V8TVFOIIOmkBPQCXfQXn
EYPc2JOYTMTOzEvCimEFIlzLLIC1G6kYKcFYf/T7oMptwj/8kYmTs+KAV9xtjVILs8myZnnnM/Fq
HGfL5j723MzTKZRQjk4jHW96QJRIayC9PYerqm7VIPJTeym1BDbmT+IgpnW2ga6UVfuv9sD2nqom
IWDaLwnzwHtY+3RdgWCzop1Dd9HjT2uqNJzn1c/pcFk53AM8tAmZiEaob9t0FZ8yJb8KA9IWEk5+
KTmqfrnHyjjIETc7xEjfjQUwCj+wnsqsxImj0fyZ67xSc5IO5Y7HoN57ZCZj36iA48JgoxOOmhbB
R0Dv/M2O2dQSdggi5/OxKUX245XT9T3LCWMAfis775o6Y4LTosMhGQ5yuh1Bl9ZtZbIlRkq7BG5S
9kO6xjMeUp2gR+rJwfQOscqfHGxittPJVLHfJXYUzIejyO2hOPzaAtLwgZfqkq1AHnYPsPujd0SV
94hrTSq+o40SypBz+8GT8oVFjSS1MksnapBs5yrtY6APbJSUKztSRGSIS+uZx70NX510hj4s1TnO
GFGnh7z+aEjS4vUE7bfvo30Z0we5HPXIaDYOfghU65x11PjuBPW459AarT99MXz1BufF+38YPanj
95fAtJPBdgfjXZxXYCHYtCXpwS3eEuVzbkcP1o948bQuTyhgyhqcUx/bxlfvwHSrDpKsm+SkSYdc
kczJghrHF9WKaIMevhUQ9aYuDBz9QYUAOJPXwmjxDEKFV/GjVsvCqGLoBwCgAjKhGBYfbQLjNHwb
nVdVH9LWEcN5H+hUOTh04r15qUU5fuE2lKD51te8LrQHGwS3D1LgI92AnjPvvKEFSlWm0Fja5bsz
IjuYsxClv2lApKwCzgzFO1G45CQtX71A8NXY7JSJlSdg/apNwpFpKkftoQFCDg4UnIJyMhKSTH4R
/yg6U/Ty19qzvN6H8CN7QdkWzeLz/rFCV3mrLUjIu2w75rfYlMc1WWBdW6ryd+afJt6t9l2wctlB
bsxN4GIR9Oo8SreJm6h57/dR26z7aLxf03BYGGHWyYTRtikeuB3rVVhCRC+uPHzbNwMP8RawEvvt
98mtjLoMAzOaF+lYktq1ad4g36FgSwGQk1GPeUuiItZL5qZ1YgQLmxhmPeyIew0o4iYj+VzAkCcZ
ZFSwRW7YkJ6MS6by8XjTaavFAPIdhXDEWrADXe6PuOP2YsM9bJcI5mDHoG78PL/VIfC6qewA3B6h
/lSfni8FWWqEWF8ocugOAA1/yHl1FVlBQ/ZlX+Y8lY1JSo+vdN9JRv2VQtit4r1QU/3b1xeap5KP
OUUM5L0AOlsDXQo9vJajj36/+HuRj7czt3F9tXVSA2MA8Wo5vYINwmr5BMHmIVk6AHyXdK4E3xO/
1L3BXyoM3JnHLw7WgoWnCKzVOT50MkoRqEyteH81rRZvVO02k2oqt93E9gObUf/k65nlewBmAKF2
trOvgBO/3P95JYXHnWwhs7TlnnnkRvI8XhdIQdEl4dq/Wc1eBY8rFPR9qCNlxjkjo7D5AE8aum9p
IDOd9f/mHa8u/i4HoaPfmWf8Sx5RePp61rZDf/LicWm9XECdCoTr683BW2NAkAeqftK5EF38nn25
aYrC/lK+BzE13hMmlyHFYXjf68osakiLgehYll/eTLEj1fKf3i7W9bW/G0IpDDCs5i65asITpwWH
ErVLctyqVZUWt/s2QR0gymr7ieE7SZdrODzU87Wydf0S/s4YKxjXpFOvk6VRX/7P8U+4BLqSyj7m
v+NnDL0IT9F8zAyX/ELiE473ff4B7IKQwGNyhIzEIi5919QvlGUtekPDlWZBL3hsMnDVfCgUxE5k
BRys9PvmEvOrND/0zFuWjubfEce2T5eADfdZcPonELJrhL5sa4psgX7J06qH26dMhJsDbExhbpwg
l+y5xO/XQRnA/0YLNjFIRW7b2e+HWd7ubGHDSW5vYApcmUTvlODkFcPXHlAQ0wV+qO82V726+g3D
x0c6YmUphzHtYZ1crCVl5nQBeC1RAGBfIxAxravp3q6rPuK0u8YnOeEPTLK6hcOKtJ/wL/3YLdG1
0Q+t/78ruXvB+kp2r3Iyq0G+mhIsai2HUUGmVg3rXbm5g5hqtqnI0tlSO7r8om7QShfjtN5ZIoEN
M2tyvll5On7IcmpznZDuEOyvg/862wl9a/PVOFkSKpcGRrT0J8r+vjrFVZyYIWGh3XE5ZwIAFCLm
6EwIPyPNWSFYEaUiR7DUWPX4HFM5IhkYOKHUI1CQFoET00y7CxrYyUOzCUtsF3YByGGgJB1UmNEZ
/9evrY3GTHYmMAAWbVH7FstMpjoDbandHP/UV012u/KF+8QOFzU5pXMe3lb7q9nVm5NPHsJFcGmQ
kt7Zw9JnYp9afQiMge1kU7LI2RXKxjDvbTegLC+rTkxGtHeb28cVIVmldnrBk72hknM7lUQ7e+gy
+Zear5nlc8xPZe8MyUsnYW72CEF9atecco4XRgBOTgmSWxhGveZ/076NIDRVloVALnhVvKxQSY/d
K0stFPCtPl9gwklskGxg79Qqx4jtoCt4jeZ81XDlhgZO801tjhEmvA0wGgVJB0jP6b7WGzegDDtv
I5INsilJ6YexxXz1FnPqQG5VQYmqbHQcGsdq9b+O7DRRbRtRTMYUVSbgjytCIBaL9kekeMrR5Ank
1/FkhFGUfxDpPSXr8Va5w2olHxB+HtEbGOo4ZaoC+T3ZjEbHE+oYaoGqxpoWFma1GvvP/oTAFHJM
3g3QtGAmJ6xt7YtCDXRJ/hHltr83rrjaXC672Drp23ZLGAmuJHAG/YLC9it+gVx0XoQJoFrO9GTU
AzjszJaqwvSdns2wMfoSy9DwN4/c3j+khZ000bVsH0T2hhtIS5rr0tg2kGlk3811AdJ7x7NyW08R
cAZD+aPtsT+0Uh1DLVJJZ6+JBwiHY+TOH4k8WBKa7DR/oGyIa+DxcOm760DszJkH6ue1hEWNtN3/
T6BXgjADXjLFGsL3kIaXops4OKlm7X/+RG2YX9s/87KMSDvnczkuFHgnlCKbQclOkWO3ohpVAeN7
l3UMoAEkMW/Y5IISegxdgDeTYT4dx/vYYx1j/4dqYbhT//4VYcZcs6OAzWGh+a3gPiQF8DYavfsB
PZcAM92F7RwOEnG0b+jE3wmstO+NTzQ3jkqYwczk1XYL6yRkeOvDhgeenRBpYwnmn6wH4eT5KRSk
6GTXLpgf+OqZWN4ckLiYdy2q5z4LnUZeOczosCthcbJiU7IRDzq4Txx2kP77G1LWx+WMTH+NlR6L
iB1rmBApwKq7xolPXlJ8Dz84bOhVn6lls0diAQZOTIYlvjCUha8lrWUKJTG7BYQMb71yBzw44T9t
rwdVkrRpseqVlN87je4sbBn/QHE/vCrhsU/rp7ZyHLdM5SUrg/ZGAqho241FKoIj7+sKSnCgLSoK
G/FU8V/4JfHYEPIPTHX4iz94qehFCKPlepdf0lRwUwlEAzNKLgbYEcqF8gDAHsLiQm6KHS1KQjlc
zhth5Rr+b5Vf5wJU7kcKVz042iTF3OafN5hAl1UgG/foT5Cdp0lPFvZVkuJZfYn3YpsTJVlq5Mxc
AxINIGJHyfA/r+8ahHHjiTQEegq/bKvy1R4GgJ3+lJ3PCJlHGUnzBw7F3ZMoziixOU5Wcc3AUcla
/0QNkZMp3axcs/NWZxP46l1vPhwd1WLDfuB7VMSdZVcAGoa8WzxVWn1pQF0TQvgoz4G7xMrSHSsE
3uuroQf464W0OfVWwP8ixe2ZkvlyWaX33InxUBcy8h9c4aopPF1vIT5VXweLXD/ZGSGpRMegSPce
GdXtgsT8JyuL8z48QpqiXIQDSweKNPUEFl0SbWFgVa3aN6VOJMeiFB5wKN5TToVmsgjkHAS0FF/2
KGreqNsLI8u98u4KiETMWXicksx4x0KQqUwB1f3mmDeVDG18DZH5FzX63mm141xQ+hWiHLQEvcaB
9mgWtfPxoggYztZ/6IDNdoo9GtzTOHEHYJRIpp01jU50iFNhF8SXFQnXHYRFSKE55dVkZlZ/OVIz
w7tnslYGwmuoGFuZ4V0U3/ATdQLIz/umBN7lrPZahl0oveLN13fapKrvu+8u+4R7RymE1Ix7fvfK
wogAJnnLMsMqnLvvBwISOhhcVqCoBIaI650tfyqq/3nKrzmCWj3PUvvxriv7B9zkna+yscqnfESS
5w0vFQkwJ2m1brYb5cpe6ZZoDbw414Jn003UnZFwyJwf+763tgPfzoH6lbNVUmwrmgXc3Rwk2MxR
CkzsL8yNYfYY+1lONz6udaP2XAx1uafm1AJYeYquGRt6m/XFMONEftNH4x2wfcVByiBznz9zfbn2
lg9sdog+We5fLBdfrTZ+eIQyCk8b4CsC3F88RdSHGCHzkibB5lr6MPvwRAC4lYZJDV9Q90FXuwqr
i2/kMzAvilZRc4XrSBXbxiRVNJoNm2IgiNxAdQFrmPqGA8k3IAR7h6t83T81Sn80w2yfOVV3KIYt
mnZolJd1VkOesqS2RX+xuAPHd0E61lOGJlgDsnEv7r0jXwMEkXoXxj8zicSSm0OgAn3kIw4PRvpr
1d2H4FAJ/IafO0Va4uCLsdaEbzH42QiTEA8B+OB3sgZGQnkwt63lrF6GbtDUi6waC8mLFBnaCHv1
aLK69583mXkTUpBFvtfaOqDyFqmvfLwEtNMlrZzWzAS5dgm2MU+j+PP6eBQnwIcopigZx6/PKj/7
Z9n2I+TX21JAz8b+0MICTzkLLRvGW8nD60Ou578tkGNyk3ORDashQSks4wlBkeS9atdIKHwg3Hap
oMvkHINkMfanplKtcSnUiD30oCplPXwqCGFAWTkbWEZxZk9/wV6DfCu1qlnfkT8BCT2g5MO3W+WV
C2kfRG0BPHhZ60zjZuJ2JzljbnJAWbm3hmDhTYtw7o1ARpcV3xLSLpaau73usKdwL3L/rfgGDhYq
HQfFn7Dnffm7YL4s9oyRYvKo7oheCvi119HzsLg3LQEriYoA3t3wcCgKYIwzlfgxcA9OISqapwPA
4vPbNeYmiLxGpcJHeZoZpTLk6elnp1BQZLGvlnYWa9h2HLFd3eN6V9fxQvbC8jdQbmSHut7zNH52
/OlCQqiGca62+WpZzv5oXsJyZtuir5zmXFiEx2fHu0IpHXqtKvSXOmUYGmuXfhTM4uyw+YFxckhA
nawTRIE6nBnn1UAqd6TtRww6XUIIRo4Q/yBYkh+9iEt9VXk9zVGwS81iGLBNx0rXkgNaf5kHpacR
Zxvf0liBygQYv/Bu4p8wHLpQOsnGYxh82QgFhajbmWXKVQec8W/lmkvtwup5rivEi6Me7h+fZ2+O
l8q/4G87ZxH+BpjtjiVn1MvaCVaLLjpy0LgmqzCM/1FLxKFUu7a0uIc1+GAB3lES9timkM9JqSmO
YaMrwY6XEurtg5Lg5M5pXBKR4oGDshFu3CZO1bs4OOn0ttzpu2e8ObbVfhg5QUnWiK51fDdVI22n
q15NyoXuhXHFRLiFgaZsNx9fGOBHRBVZ+6R3VyodOPcc0tNmnFoFGg5FMbo0v9qOR0zk9v5qTCJi
X8ctXi4gsR+Y3fCC2ceWdg1VMdylRzrlaR2JnDOm02l3vJ9xnjXNDf/syFwI0AyqzlkusBt4X5Sv
BMsaBkHj4/tIDswQKv6sR0Y8dKSD74cXM8znFkiRMmkDcWl0AJ88lpiORkQPORT42tmGYHrWB5i0
c4QfKKmm4Q5642hPAXd+j4g5d1zRzI9e5a/ZOxE74+orXojZ+dd/13T/hYx672BdrPf8jNXK7xrB
lrDP2lmb4vkw5f5uxtGLM4zAOfqTPJ0kDSIU0wpeNqkZN2AUlY7ggZX5s0mw/lwogPcl54EUD/eC
7odC0YU7n9K/zTmbnpbN8thrdL4fU89+jqkPlCCwTZjhwRScD/nmwv9Qa45JMdpVuTzEAUMt4dn1
G//kVjOYbmP7zqx1d8xMuXThIdWD1oJxhMHCNtcD+dTnIuDAZpsWKgU1lGUqTugfeGo0V7flMgpx
ZhvEo+P3LDrkw84VDXjmwEgYJ6xcAPKb2Eob7i4huKzqlgFhL9yVby2juI1jLplTRvT8mjL9sFSY
nTAevl2CLYCBunmccdWQsVHJ92gBXp1jpmMemrSykmb2hglZ+GBeAS0sHIUD28jNV198/7RbDM8R
qcRQPz6phiCapaUXbk5DUY/IgoOuROCqZlKZ2egG9Ow2+WNSSionJvonXbfAfND0O+wAIEoFfoP8
Nw8kF8lbEemy1YlSCvBCGe4SWttrJHlb+slyZEwWGKnykFt+bxjJJUWKo64O1NAwZ8vqEx8OqxBu
FQhXtCaVHEMl8cqOf1j8SCUrGKI1ahoSUZsIGbmhmf8cqz6WandpZF09xnhMo79/+ZsIN7eqfTRU
rRk1PcZ7uELbKGebxVHBJYZ3OKY//8uS0DAg5mfQZx8kHtEfL7A09LbLFY3TmcD+TaJJUGOzsSyR
JUP4GGUV1PRVf6a7moxvy+gi6C3V7XTrfUfCY3TCTyGkqkinS3bzaEhQ9bPgRuLMz7h6eEGiJK8r
XrUWXeg6kGfWuF8sDDPLJG8DRxVEK+LtmiTnyXUU0+pRR3J8COA8LFQ4MlZktfItqVlFGXML6sRB
xKEuOAVw6CBUJBe3Ut1pKFlikMg/yDipuEI2PPWufpC2lZ6UsvJZZJfUYgvwTT9MV5FOa9HtcBmG
Q2qXEHN4feVwO69uIJbUXlrUvgv7PgXP/dcphLFiFe/XtesGqPs2Slue4WmGl90e9ycYkGYsDWpK
zOXty9QDGolvnjmbMwca3GhOSgrx/CkUGVqiuCJGXBsYgoRhVNJ8ZpI+plTKW8xuSvWG5t9XaLoT
DkWNhMXHRQ3206OXRBNvUkoHg31vuNvLkrlW6vSHymFBUjoWNYg+9645WR+NnTSmYY6Iyxg0+fwq
nTMr2Ls6axLVGRp0vDhtM2ZkLhgATnHlR6VTPGGixeRGtHTZTiff0/1lf5Go4qt00vEL2wyxAnd1
Ty1hAbuP5L2u5jsjl8i9zVLnwZ4YKc/mSVnJhOXZN0ddmvJNo6GIYT/ZgrMcL3TGVCapacWuHEnb
6y2Vem8IZWqNZq1tU3WC7k85/C5iX0Ttg30sWSETuSO7fH52AAjhgtvt/CnO6RLIR/U3NPE6EGkk
UcNB/zZt1yW6sxdVxnfVvSN+HfDxYQUSeZTozLbwVzr0nGGVhRX6j+mSV4I/KgwV/2PmDXR1y/1K
kZogbw9Me/TPY0dLPxXoQAuF2zHcGpMju+/YGxFZafdZdoNW/RcfjUe9Te3KvWh0hQjvcVG1Hfxo
lYNLFLI667YFIVHo0Ha9NqrwN7Y2fxRoMKyXCK4EWUIFubDJlgvNmYDCHjFjWBQLjIY4BEViZNqg
TKZMcOAS9XtxGpRIHAS0D/SlFH94NoHHC32z6Cf0Hl1ToortlZK+PN2PXMuHRkErPfKWnnj7U1Pz
zT0DvfiJvD8sDrF4b32tdBiyCObTY/lQ+b4qa1dO8FmhOb0VRZLrPpaJ0jANnvZuZUue5tfD317J
PteV0mkeYx9cd/MhQzPXCc0ZRG+E2MOIq8BFLWSX76++VLgLfbyf7NYgEmv4vNLhy+l1jsKoJKF0
tA7fnp44DPG+zOa+2Vxi/Y09dF5zI28rgwk/7lXnYhh1hzltkHrvKByZVmnwxM68sA69YTeqMoX5
p2Ius9LAti4v1zmBt4vioL6mtjR22lCbYSi1I5UDNsmrxZQfsw1KAL35014G1Kf4dM2hr1PeKl22
2/wolfgEUtWLMJX6N8H2hA==
`pragma protect end_protected
