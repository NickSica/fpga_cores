`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
V82h/mp8FbHcv3//3zVZ5VW10Mue/LSt5dvjsUkiSGtG5WaH8H9Fv7j37k+xy+3/pQvfXcpqBF/k
iaz4/vETUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n4WSOWV3uUjyMD/l4IGcKD1bHONRRplCKgax9lu4YRYlORLHEpckVBvOD9geZHtnlLIjTLNUcuHS
rc4oO2K5x66eEf5+m+hNzaPYWCrVKWQI7/tyX0imMAsD4JQXzU2CP3ATsQoldRyYOQZmggmbIMiB
stLQ3uoRuVc4t0kXI7U=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zgo3FUzRcS1G0FRTCr4C/JBs44dp3dv5CUvkYU2vM2fDyGtu9ekJcjDXnFGi3Qx2X0BV1gEyWxsJ
xqQkFlu/f/1mutspkUjOMtKZNCgPGDHkGfwBEPN/xT22fOBwQJUR+Oj5KSeDWe2U4t5UJ4XXcGMb
ZV9syPFreDWYOTWkkl85cAKcf/WXC6oz+tOUowqV4nSLA1PaSrK4ohf8oaOGNVX+4Ji/w6ViTIJJ
OqmPJQ151npm7Kbt4RW80tp1OmABkNI+o6h4rwtTS1IHzM6bJ1Krrp0V+2aEmmqoZkuKINjX5Pw3
P4Vi6iUmJI0uMpdsCPr3MEC8HH4v95WCnjh0Qg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A45QQ9IEoKpoNXpmniz3AuFZmGAAZIhtA2hP4/pi+Iwurx8nPI4ZkKpYXPnn4DfH42bSsec35aiS
Ve+A8f1Q00bmFgtclspinRe4YgFesk40ftn1mzy6g6sLCNXhUm/IIjCSNk+ie6jVQS7STfOdio+z
cvSm8QQePoJjzlJz/jkNhsD110PhDAevJWb+C5fforY6kT0k7ZmJmE7btahod6wU3o7t2HM6+XGU
DDNZ5E+RLS+IiJYVCOwsdqQFDuRaWwS0k8Mk4UuDiVWtU0+QLFZ/8UGJhy2ZDSYlL/8TrrsWcD/1
Vku2N+fkWCj38RSMWEEe5TmUHSSzP7uBI6QwVQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b+wEsHDGMmVXUM545W/2toIjDItLsHFsIOyFDid8Fv6KhzBePVZlc9t2c1LfdAa6UEpdqcx5kgIr
+oVEglJG3R/fb6dRp2mvlu6+x0AYh7FK0My5t84q7uKZ6EPBxHnDds9FLGQdMDUFv8E10WtGrG31
lkto5q+L5WLAzYgiD3//MgdbP+aqLc/75XWIRhw/PfRn4OqyBU7xSBeoK9TDxBwOscUv0cQ+dauJ
dUQ0W2ZCXwF6cP5c47k76Ikfu69J0/IO+FTLKMkjAB7Wzsyqbpl6RMVdJ/iYscNROh1xxo2k+52w
4l9VnVKN7wTWZdW75B3V/MsNTrKb2I6dBdveDg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyn/owx08GdB/M0CwlYM5XwpK1DLRGgNdNGvCa53fvz5ftb1LM2R7yhWTTXlm8iqXlg1S70wvPmw
WVO2ZNZ0csmDdQcX4HNMiokrI2gpR08Dk8n3nzdOhqyFyh79/eVJzQItyKMQmJZNCvFfww0mtX5K
FbNe2x6ria5jEBEBp3U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J8WwILioFJtk4e6vNsFHYZhWTjvAMbsqHcnvhYKYzsY6fpaoYuWnjTNNNxS6JYZj7bKOFgPjdnBA
rKaGPLghV6UU9fx6UcBVLjNOj95AU3CZPEjWGC/GqjGRPxOkhGtDka91PZuOBRTBqJT8F+5qIgQR
vO7WJHaKezpaUm2zbeC7+ShM5p4Wm9L4dzJ1OuUGZNm39p9FbORAZNzAWa35wpfJ6PPOgATFMi7Z
sN0Hg00oxMFCKSg1bxvN3p4iC3rVT+wV6yuzOecq97B7Fu+tfvP+shqnUhodTpF0WYfGWHeK9ocM
Mg7nt62XJybi4Tm5rgYGMIIM0i67934etK5Aig==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AF8EDKLpUnsf5U27caIfzjHsL1dKCT4FvrlOxjBwD3ZJ9vsXwbWO+EJTOJOFymKnoSSFnuslr7C8
ZCAbkJJLJrLXJwfvC9hiPRksxuYzuxWrtwsjJd+5KWtue3gL5kHClD8Tbo/V+Dnr3gvKzMRNdFRz
i+4p8dC6/32xR0/NITJMYT1uOYu0oBFDHGLR02Wn4PqghcTR3gQMVeL0RsDhJibeNnf4Q0NsKqCF
7OscDpis6r9ZAFao+mdpLGI93rreTlZvJBUPh2RcpqOjL/8IUv0iM922KOCZ6j1LtvD0igXehvHa
5hOx0DDcMjOoejqJiwIqLij0FB13lDBsu+fjWw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16992)
`pragma protect data_block
BMP9G5RAk03qFRu5UmzfhPRa2E8EtqJjN3D5ol0ioUjjwZl2c8nccWTnJ4vf5ZiLEl7z84bXFwuE
v53YI9pjuQTK6mt3ZyHLt7eCH7HS/6egyI+0gGNSg+KN1XVsjPjrGQ7gjPzcphQtQspuciLvbeXK
slYLK5huTlKtBzaI6KUgbmr6D4s7wbUxaaLe7yXBWL+296o0FPDZJtvn17qIj3hAkABbqQu/OhkC
qXZ+jXtAcncFP1ivmrgm9WEXFHBYJdWcBpP04qok+Gr1Hja9HKXGbuii4Su9pvg3qkg8VWS8CO+3
Bibn8dc18hb3u5RpVgujjazJbwyGjuro479YM7fB+hsP5+YwEvGVubWB61VF6pGWyDSq4Rswoi3Y
/+DZn9YRhR8ceuMTHfismZ6ns3V/PCCKvGIt21umUER/dFJJSfsxXiDm2NK52Ivlx05KO3lvT3iY
KX1WT4CubwVE6+TGV30fgge7/05hoZbZq57OgIHWSRJ8yA497AX4qAiezA8XQT+ZLXP9kxrhf8vO
fOKnrvrxZ6XVL4ucAczjVxxJzAEi8pY/ISxcs8DROsKO5OnhmG9BFupHL6LRIN4CAIIsN+31ToEX
EY95C28ZXN7YRm9eTkZDdym6W8y6Sm8rsqS9sciDUIIkWXI8b/S4/LAUsqu8SJ4mjbEleGjvD53O
h/vZPYS0IUzhey12B4PGlvu71dJ/sfJ/EBzp4rnX5EDHW9XBY4XzWAXEYny4eVyTvx2EvK2nX2ka
PxZhNuINUpYFodcebMlXUlRKdtaGSLQcMe1FnvwmFg2TgudMm4Alo7FFzMwftFG0sg494mW2e/qU
pI//S8wUf+TAmyNX82zFUrgVfcceupIqr168f3nV8O278Rc9GWj4lJjCyJ+9IrY5C2Z06WT2No9x
6wkOMEoaO51E6D3SSFtsOXTCQMDjHdsoCs1xx2feDGoQvVdCCngZPmU9RWf93DypZ91JBoIkwfsx
re+rtrLIS42bPOJSl1+YHhFXzJHIGptvld8zh0rxYmulwMmed9XzkSJWIA0svhSyr3FpcLODGgj6
2yXCs2kBWl2r82ouvoEPGTnnl62v39yYlD4kCpiwg9XjQ9reIuY3JoPuECGbzj2q2cm/QoPTADfK
qj/cd8TivgrwpjcwUSRrbGrMdyy7R16EpxMZAnJA9OO8Feca7ug+OARpJ8aSaxu9lg8NLmWoFRNO
5T4+dkAkWJ4ARl9TqpcyDT0XUFXU9g+IOfNHbyq7RarPveEAW2ITwu0oFYU/QNBjwXyLWOqoy7VM
GnKWmDm5Vqz0cKPjXk4+1lq61VFXcYg9602mJnOvsuGxi1HAp2MKmgpWFMypokvtiouGtdCZ4+AZ
+ErL88P0UEJ+W0Vdfzj4+9XAfUeG4li+bXjYie/Q2sB+OosNfjXtouw5BeSKap7gJMqt0gHc5c71
Zpz61wqn8Gpb4R+F7R2FW7jTWsXscdbv1dnm4PmTabsbjmFoOe+VBboiBGG2wSxuLa+DRvQ9Z/3s
euui67p5lu82jaQ3L2OaMnZmEVOVbFiSQj6ucmHwultNkBY1iwl2vEPLrs/6CILmD5GfEeoMxdR3
58Swzh+fd3Uz63QDI/ALkYGLG8j5BQqAz64og+Jpucc6eGVJWFVCZRxCsRxCllWyw+k6KrV0R6Gu
rtsKzOC30edQkWUDDcwKOC1J4ygcNn1NAtc7tPMLE+Z6/jg5rPYchxzziOBE7mAHuz+HeCll0NEJ
NEZIRVsuIWUDkOQXRkEr5qVXsnKiJc1rjcM9TrCSVMgUpkr5JLOAsZ/4WhoCY1U+jWryuBOSv2yc
15CEQeWJ0WMJXKAy98vX56M3hB2Ho8o2NxjuDqpha/JFQKuOtLXlDdYBD9RqfQ8UDSumDxMr2FRQ
CiKhK68FnEfz34/X3VVGNF0l5mRgyJDojxWGM+y1fhVdx/rFdmsvhnfUAHFoE5xlY3amv6werc9W
WjWtMu0wKA3tC/t7vFxlr+yn/ZOOg7DEsIIgWneVelTtv0iqlIx7g/TaAhJnPHKXeeHnXPreRNli
OVPJsD03JLfPOsB2Al51KRlaW4BVSijLa/mtERDoH/pAYp6/T9zXw+g13hr26IaqpsTc5fVPR5Mi
R/4hJRrQyn9AXG/NKDj2WW5iqTqbOVX18IuyqHeqIwGPXMr/LyJ6Ckhx2/Jzz7AwAuUxsD1nzCdK
fkvU1EFWzSq98xS6hgZzSrdem7Phd2C/ZDoOkYMpjYqronF2Vo86sVEAO1LDWdD9LD4oai6pfdpe
d5kMQjosve2nMniXTI+sMfAbMoku62ZgOQFC3E7EzCXDLLqeTfKKzg3Z2jr1ABpONLd3EOOqBnqS
rlKzwloOlPBveXPrRfCpwmNbSo4+MhlwrZrqWE1bT00Wx0f/tz1JOASfftaUtYb9jRaYxfvYCt0p
8J1qXPMXXJzHxqhoODSJ0RpHS/7IZMfnUgrDxWWZBtxK8pbdKdB1R/imfAHeN8ZWTbvin/CCFTaR
Kjmkzl5uWROjQj5T53+31FLbS7uIb8pjMnSsJyeGTMq8n3eZR4+JIgoB8Ss9aVYaPax4i4szt42c
9n27DoP3gDclX9Y/OX0IwlsvWtmRULPcUh3ef9I/b5MK5uXPAm0mJ3widzIo9rZ4ooVUEzPUT+/b
6DEmfr6d1cvFVaWJyi7puV4mWzC45uPU2nobtvL+JsD7SAlL1qbmciLxyb5we4flM195r5vT6Gqw
UmLAMjrE2fdKMq6C6Kb+oIoy612PLt7lsz+dIu1CbGMfGDtB+/ofbadYrNGH/DKo8ebvK+5e8pko
k/Zki3pkCQ/fo9FhF7/G/yBOA9DYSSrPCT9RS3RvIDPoa3g8jfpISwDqGIfgcDhS98qt2K7uxBmF
jBZ7jWcEfSiyMqKRlBvJmguTp4lT5C8LRZdEB5P4+Xu1W8y5ziYlGBoubCU9vHtLnhH/+g6e5ViB
k+Kh5m96uFeSbgFx2LGvw4vBVSX/506M0D1L3b9eJs15zIFR6p9AxTYZ1e5OwPkd76ahobkkUtfG
bth+9J69a6iCZ/W8INN5q4p6QhF9NEHfolPlWYM119ELHHk3eFVAob1sghcCTzRjTsyhKDXKj8wt
2ajTt6hiAL1qym5OhRd8cAWBvRbRezm4A68zSe8huNG2yYXRuSMqReagXMJcQvbi+1vuhBLgfwyM
DDulZz5dIHDjD2pEyeIbGILS7JaqOp3cl2egNOi/7Jw/gMyKWjo3QLBYO4Rth9xduO1dIGXZHw3n
qKg77/lKxWFoH9jzRpD9R5xPhKmVJt9z9PLQ7CWd1AljJUN+AtWq1jU9aa8IxSVOsZGLPIzoTzwT
/l/EZL1gcTU25iOVjzNffm/1Kp06zwtpulfpRD9UqjMolG04uS66tvEnbrxfK+nsKNd4eIsl6O6T
Uvsnw0tjLM9fbVbOJ4oR8yoy6aV2ssDRjGD985GQcGdAVa/7QZbcHg6trgAcBBAb/maK7MFYIEkC
V0eV2kcUONEn4WzvlukT/K1tw8NJjdaM2Hj8+dY80WnSms+05JwREEPpWgb4lH9iG+l2782RNgyA
eJspFFg0rkpWZoulD1ozR8zVzRtNET5l/mb9T4JhbE3tjTA/wfYHl1piBV7mAYw6saCiJgs8xkkh
ul5tVQLJ+bqmWQKGeV32Tbv6I00UdPMt+jXVsLuzY3H1ZOsOJ3sXE11Mf642HxpifbB6L3df8Wbs
4xuhCaGrI4aUtv8gZi/g/Lr3y6m6dqyeolZO13BUW4L1oPAjJNo9vbO0q5ZAZamSpa7j+4AbypbT
ED4fiTe+POYZLp/Ko1mTQZWaKHOxwA26Tv78/Bnf7lt0XPxtW5zyskuLaG5o7kcTHeBcEC8XPoka
QX+9jp9NBDTsWJvffyxgrCOO8bxC+rGlbrZRu1JAXEVGvhfLRZsNUzkgzGc5rmYCt3DLyAwX+EyA
z9QxB5plDTnOo34Y0Jjcbv882PKfM51aqRJiMg+35ONw7ehd+TGL2SzJcDxB+Relmi1Eby92Dh5L
07a3oF1hhNJ75GVOb87azjfDx5Z9B90dIBtySmZfOBDeCis+4v6htgD+RJZcXGAPWa7dtI8g+lO8
g0cduQehj+uKhbdCM7OOTHh6xbN/pH4OaCuTUEyuLRIFp6vJak3FnELUjSsl13QXcOEB4XVQtRx3
oVFfbAw9HiKmvZ+L3dr9dcNd4JAXChn7fDYYgvrovL4NJ91CzdCOPGzhAlcTra4NqQsXCsfYznxX
QYQ6ktNOlJyNFKQJ5IRn5imfK7H6T1fWAwKdcenaeIdI3njkE/oIklRQovdyaaco8zx9XdbFUaBa
tLKhLYesV5lE6My7Z4H2yeQF1nWX9nphKIhwyvjOw9vv4S8BHhPu+2sjaxRZDcFxzBqioNohWxq5
6j5Zb2LT+dsWsAERWR7WPFaPym60VCwDaJ5mxdaqG0RbB96ZvF9Yx6P9HPy6zy94/RvRZmcIKyyD
yAEeXHm/4CUCQUTX7mCQB+LTrYuqPY/eIRfjRxnpiDp+pQrH3w6wUu/MVr8GjO1XKkPvIDgsQaQ5
iQwOviaulQ8l/7dd2NEyz38l1D82Sp5sk4v+PLslrUjSF4gjvBaG/pR+hY3j7GNVPz8oUN5/5da7
p6pE4m7qaAie60DJuDDDCrCC1rpTsEoahGfWD3lAR07rdcjAeG9rv6HPSTPZW7USdZ7ZSmNf+y80
etu6BUicHxdBqXUwozfgzPpxILFL3zgaFhQMHg87VVPqHC5dCyLdxqnCYjn0UQr5wpvwZ6AZLzRC
Sw6Ui7YElBiB2cintDj1ykMKyNuTIPh2ATfriOc1zCrQd16IVZLdsh0orGaeIjjXQ85NsHgGIpGD
7jHJPqiT8Tehkx7bf2dJaP43QJ0ByB0+uBg3kOY48wJRi+eBmBdw3FAhcezDkvtEHpBadoTfdYFP
o7fEzzjFrptG8xHyF6x6sbXeDWQVLEOsHgM3Bh4oGJH6Z3tpYfOvcrL//07eFI4NFoxqb9iFHz7y
ODkbZePSXqQ5fqJxFV0hByxqHQIfDAKT1Xn/HFfUxvKQ9Kk5xQB/eNFv0LXPdRvtbLArV/cpBBIW
+5lpgWmw2yWoq/Q0XVmCy5A/URLzi+2CI/EMnm6yk83tes14wfrlE/IqVY1pQNdHrSgg/21xbVfm
S4h01iz5+ha2QLeoifl25b0b1UTROwIWpcc03hfs2oMnFbbXnK82ViKhEPpZ9WjHjvK6RawUHVvm
f8gBMkQpuXVoKQZC6GAoLDDYMHb7TkFZwJ68uaJev25wBLjMs9BuJ8lGk+2SoRCvNHsO7F/wcuLV
cFpje1nPxN9H34EG6KiafTnbcV4FQSBltHKSXy9pxwJEqmlw8wMISyQePQ+z+Q6etER5KIw0FBai
O+iLHP32OA6/itxE/7Fpyt3PHIKpR1XNSXSqq3pA/QGacbR2alS+tI6oC89LWt1e4WM7T3PLA1Lj
rVnL16gbx7pTVPicJvhST7iKJ9QRqifnIuVc1pUibSE/aeVKgH0nS0sq+L6jEwqzuyKO6zMZ0BIi
GceyRBP0AeBJpvRSF5tZEQBKdbMLj/lh8PwqRGkxAnTsrJlEKcJFtDvBfE2qA5IKgseTQbp04Nfg
DWPLjvOTEUg98Z7ne6w5uUV5itUBsAoO/Yg2NLsbydyJA0H+Q5hGZiUyMtxsweU+7eqkgXsogeBo
e9jOrn35Z56+krEZW2rjn9UjLBtCEFB3JSZmx6L4ajzWo4FNem1HbcY6nxhFGt4A23GTq+/GmibX
rzQfoKVMYW6Klnhr+AaAMdxlNlsbcc0RHDD7wn5MqVEgbIviNixSfVvDxPbnyVA7PKTRcG0JHyaA
iSwNk6qWXGK3m61QL89cSmLNvOHgIcZPUNCqjwOUz0FhBvzkUg1AG0pUQC9uwDtYWnFW2EIPp2zi
fKI4/vKyVEf1rupzxAcHVEtUS6N4gGVRELLKwj+v7H+i2RqOcN1IIGoZpQj8mDoeFQ0S/hJAAPs5
fofyBC6WKsV+QkJBlJWZox+KYgvE1VUsI6fuh4K5OngOwmVTiIrVPNSFYeH405AOJ64uZypY8hCZ
iFInfx6hLAMxVUoRMI3FSXfHbMU9nfJOaa7Ubzl7votXguyvw7yANu1ViqAfOJojPXcFooAojm/o
alvVQz8MXYw0tn2iMh2e3Khmey5AT7hDIihn0MxvfvAnLsuMYb7TToXwjHCv7LOSqC5SsP1UpOo+
pE9tcJDTvi/Sb1o5Vgk3SkPeDW0PYJuWZHmU1v7KLUmk3B2w1PMpCx/c6OqZdSHiSxG/MZ1V9PRB
or0t1vmYXe1pRw9um136kaczieKb77hbq/ehoYJcCi+3RX5s2KrDWEzWZxHYve9XRHnr2qq80jR4
IA9sIp/Re69DBU+lE7m35T+azHsrDKOM7IYUvtyJo9hMnoOaDbwwfH5NQ3ldHt5uOTPF/hP6FuEP
8g/18QTB1YwxhiS1MJG4bI+7JWw2C180JZ3Fb4wLU6jlKHhfFa2+m8RhDhsyzvyAY4w6LDDflL8z
byTdvL1lPC+LHnwpmWOdXxs/GrYXPjq/7JSE2peMCDmczusJ76NpHesq7VE7JrKgDk4Evchwkk7U
8j/4Ha6GSrHNQkRxHZQQ1mlDErbW0XKYwOxsrE5v6vuDWWcD73UsWPCGCRqQVMRIigqoL53alqNS
O01QiJ23jQ1KW5PTJ6ekouqQpAVBBYG09+gs74onxFO2o2CNxVNN3JRVpkcGrMj7Qjo3hzAlpzrF
HAx1gCwvAYyoPoiy3yENyTfJw2yo0rBBiLWzrF6lyvQ7YrdI8hPE6bZWqF//T9NIMrU1/NToidWc
7VeNi8KGwfAiz03lXwoXih6Zr2vz6dT6OqTZweLWXDb7jOScUF8oQvSSBYQOVVkyeNRVeDmmOdWF
7xc1UhgwRdfvWQhwquLzk6xX9NOUluw5dPsIZOP6jDugt+pIFE4YEFYVLeAbyK2iIhoFJn9DfhjH
2hLpHdtOvNC2aXmqbvCuxiT6eR6R/S/dvaVowBSJqQn9TBZKOh0IN5uhLeMZ4XbbYvB1G+yyPIsq
jjyOeTr01HcnEvd6SmhQp5SzGZzqJyFPUm02x2dIs6tByKEVlc1+4Ni/0uAspRAipIKr2kFVP1hs
DNvt4uLAi5SCcfW3mA+VFHPFx5ws9wcRLzMvKXPR5fY1jvqdFo3VW+3wOuEgW95Unq78FFXAr7b2
0xztHbSMDqNZpuZR2CgUkNr4t7ummzvXkleWPoxPGeIu/7DluLmC/JcUg2PII22wBwwj8radrXDP
TbL3tsdQ1lDuD/6fllyHolxL5PIqnaYewm6L746vHnvCL2S+XYEAgOIPVdGWTGxMk/3GfggUoX0T
BHKYbL4NVlY3C0kmT6MJNE4ibqURaqpnsYvBnl2QXyXoa6BvIRv1UoxWsS9PhMDCYUnqLk67D+nX
zAvBsOC90xNdjyCLeJWnpjC197W27LVw38ap02ePfXPvR2h6i+dGl2mlteA8Qq3IGV40iu/GwGEg
CBBQ4visyhajtrrA4jXddT2S12iWuypJf6xxDrM4IXMTGpMsoxPxwhV3HRUgqoYNP7U5htsR3txb
FpiKsQyU/ZR1Arr9nl4WsvUu12zlTIcmJxJlXBdG8dZfZhZ7223aLFLK3xX+9KraJdSSgbsolaL3
tRJbF8T400lHFkL9v+e65pekYfHxMSpWm5Xrb6zJi1xBISLNhSGUgVCIL6JTgKA7zmjCcYgRO55E
Mow2hsxJWPGN1SaRLCFrUZm8ffbx1Bsl5YGWD+geVpTXTWemX6UDXZK+8v1kl8xl40SYqq4ZOqZi
TBN8ePp8YgZOhUgipU/KvL4+Fvkbolo+v87l620IiyJ9NQj/HAjVy/Qlx6Eb+doQCQx2NuBuzej5
Dn00se+CASmI5s2oOvh8WBewv2uhNGYPObv23uwZbteUrOlyK16Yk8UP6a5FSCOOVqJq0guO1ImO
CEi/Ys/FviWY16h0dnl+c8A32Iay2G2YdGP/Npq0/wq3yOF26MIO1BiqtRo1qDHYqI3vNFUKkJq/
x1raHGH8kKZbc+kPBiYXsP6FHIgmYSRK3Jy++7d6ieKaz28clLPQLkUGE157N5hh9EpWQo8xZvuJ
BfJkGNXdSKAAXRmb/ZKMfUGVr4sRFfdswH9fQl5O9Bk84oiHHmmECXYulrSSR7V8GmF4gDxpUgkh
pOK+VriHrPyk1SOb2EmQPGRtTfb8j/3E7H72yz91ToAcKh8XjnaI2QoFFAhbgN4XBRC6gJ6x3ktZ
kDbh5ZMMvi/9g9BPrAj6/Z/ZGj19C4U04n8Kw1fWiN/Alvf5FkfHY25IrL953+N6TepDXWHdJzaI
C8Edcv47p2xQpcptZJMeJlb9a/yCEjJ6ijN4gXITM6+7wOJJc/C5fqgeXaP9eQG2AwBP4UKCV3eF
LwQOChDgqs8hRxFO+SLi5e72iUwyqOxmDFJZo1T8xxukp9pNHgjdLD2chXp5zy3YFZ5yNNA2kikY
GbMx/8aB9vKp217qsuOS7N05MTaQUdckCUtCAhEKO99X5/DK/rT8pbZvEUJ0pj0MiIsx4vm3WQBU
blUHkxSghssxDrBIgibkodDvKHJ8y5a73MExmKfItSb2emwGxW8qgysFB6liBbyvBpWqifOpjQz4
2k+Ble+ui7OjAYYd/zgv2R6wyZ776QdChIWVp6G9toDw72mes8crIFLMhG9MouVNpWdWiEYp1/27
nz8HVrb8BJLo1qwHG/kP/NwIcF2KchNbCgZ85Y01OeiXN8h1FudAnmOkdTFdsq84ITIQiS1ll1iH
oumgXQSxZZroYJP3zJUZJJqbmLFndZ3aTdymwY4dk7G3xtTX7ZsJd4PwmL8+URodBcUNOr/D8oL5
wpDMVab59I7EsBV0J+ejhs8zNLF9EctrvHFf6II5pIS2+Vhe6Wb7Ge98ba4VR6bS+Dr9D8DYYM97
ClUy1DikOhxqQiw4ZmZ/xzyo7wF2dZnKA+LKiSU9jHWKKPpBp83cWQ9i6lTaSQ8Olx0RAyrGVlyP
yq7GNxfDDC19Ry8Jn1VhMjPJFaqbCmL8bRGJrSzYCsfn4y2ng3RJPj//JpknlwjZcmxkUOjy/rOs
lrk7pukLfgWj3V+5P8YcgANIkZDokzlCA2kTw22Lvl9ayLctj5pNzoldXWbz9UZzXtmo40Wl9U+8
Bc3guDOU8gNQZjhr2q9YFZzOqcU9sXVzH4RwngbeXhGIEhhsOlC3rL47onZzUashSFy22DXaIMg1
w3E5Ei3lFE7XjWTUgXguMBxEQKrMKtRpYp1zefVIG41EC/oqGEN0spkHq+iAFCPPisBwe5+5Fr+G
44XwBFMAIJ3DWkH5E0oKp6+if5xq5/+CWL0TNeZ1adNFtYuYifLWfXg1n8RBNk18q25JaRZe9UZA
/rjds+dTDQpLzF3PXVmu3qmQ2/3ZVw/xuzdQVaS02lVnQCXmsgiAHkDfL2RSNVtkeRRV4/I7UoDu
zLPxazSxv7zQaTPAhWcsisBjwZwoCBA0yFhSltUZxc5GI6N8qqUUsWAM0VwT2A1+2ljz/TGhN5/p
254vlp6+GwqUqX1Erk/rgu1DFv7XYL2Mic6N5q9BMhrGp8KC8uuwQFNxUW0L18TnJMcKKFZTeZ2E
emsw+87Qlv3YS9pxUAEngW4VjdfPxQ57DNtZzlKGC9HtI7l+b+PtvSLaOOeEy1/Fd8uBL12j0rLw
biqsQMdLNHKTYhZGSc68hgakFC2KJbNpXo4USDr0I+nWxNgKyA4NjlspBczCkKTIS5S6o6fciMiC
yEbZXL2evne12/XkAQnN2/EWe+3xxWATWPlxSXgCQfzMxhLc5CTiWDfU6DXA4Kr5f7tfHmeI4tXi
Lmiw6gO4V39hXZkKVmC3BbefaouUkha+ULo546UcIddZmR6VPojcYk5w6hl2NY/oeLY57s5a3Bf7
QPVnJ//UuDBrCJo0LV3L/ro43JJETJVxiz30VgSk6rN0LOgymb37C3IEcTut9eMSw1t6cLERAa6x
fzhl/u2qiDVWGV3wh4TMYku9naSyzwv1pcKS3MQgRRPpGIn7wUHo5umQsg7VaCV8ryzOFbmsdpTM
neFeF0Lu1DbcW5yOPMTsRsJ9J8AiTLGU25VEQuQgJN+I46b++kyXIgJySXAofBDE8WL5NINENPXG
zA8DhF0o9qhTNeeaSkDzIYnl1HlP9pTlA0oWrfatjDmRJIWUsqNl2OLlnfLXpkwKDQPgioP1M5l+
o+Olbbe0K+P1j+Hjy/JFS30U5vwMnvQJPKui2a/2Hkt+zTpHnOFY21B+c4sZ0FcCCFKruYoEpPJc
/v+MDb0TTj6o9Gd/2S5qGdZZkwSNgOvWnGBeVu/96maKXUyPmN4yrtUoMTzE1K+iusX65X6cRmFd
r8oij8r1sbc840BFeliQljOMHqPsWtKZ7JdYreYhPrHsJykImKhxYVAumtA/n18AXGjBVJY6Lboi
PyE8QPPYpzmavSeM4/idn5G7HlYWJV6p+halx7UwTPHHVmi9yeTL1PthsPNzpO5RqbCbvGLJDzGw
oP2P8OVB9QNNGR6z5duAcaab7IQhYZVf8+FmDa8NtMJ94IYVDpYvSAs/O0DTfq0BuAukwbQUpMcE
PhejLqWPUWUsbnftpXxMzs+XC/HTpZwDq0tPWIqnkaIiXLhpJbqmfV5ZksIoRC/t87UJk7eeHyJj
mTslRKih6ZeC7lYVpXICe42Mwgw/WM/Y5YcFtFjDN9piAwuFZHor/530l6yak/EHwWLXQLo947tM
rIwIkVSKRJK4clvOFuUCPxS5XEkbjHE27Dvv0eUkIpPFCsVHKiXOEswUKyyo0x/mnrB6FyynrArW
8ybosPtahgIWvF9su758Jl8fPEFJe5cb9qSL74pTl/hLOW0f1ei/DXIN9fW6rB23uMg6k3JhsWgB
R6jHGVrz7XOQDoe4LH5Q/AvPCN1EgM61l8P06Re/GHOstwzw20svXME/ypJIo6XPerU1RHqqu93N
9upilOPIRab/8fs6JBOxJsZ5zBP5knDQVNtBzJ8VakCB5xXzP8ChM2enL4Qftn0c03XPYUiFs8mF
YilXnAM6lQ9hGHUtn2+uLy41FzVnbDEDwSHXrjHUvXDn667SOcml3jOWTIqUlT2eC3sIkhNwdVto
lzTDzEL/gsehyH+DBfrqOgl6f9leX9ETz9fDwH9W5Z+zCVKgP6GNLugaOoYgjT5ZZSOYar/m7PWd
IEwphhEhxKbXnfxQl4lpfpsu3nNRIHhFHsVfGHhyTkVSSIwOOyxdsIdgWqFpzIxoUZ0S6QPOtu7V
6pfmSlMy92f5MF0R2Ya0bk3z9Ft2cHeeiwcxjs8KprzSyhcDXv0B6bxM25LZzdsL2JhTnZ52hSQC
XvruRUhHMUTdhbE0DjkRFTwNcDEu/Onh+iwlhy4cQ7s7VfcrQS98csvTJ3hP/N22zj+X0aGyb7ln
dxynxM9POZXrA3HRMlsgWdIHW/lgXYZN/K9yMvKaB5FZdZGuj8t3rmPaX21r8zzolJagi2DFy+uK
TZc9U3zde601ITTm0znHSisblzzTaotyOa22bV/wMajojDFIDrrW2jSMIpMkloEUwyomliKk+IeY
tKNLuQfF47swrNsqz7L1kspHwMgOcZvit+IsahN8qPvc3M/XvT9s54VHKULbvFOJ/xrTv6jvlBGZ
oSvwqTIm7+iUWhcKAukQq+EsxK61ea3YW5PqGjWYtjjHR5bxVyRcU8d0AYNGOmJiSUGQ8PHKHGRz
5iLeXbMWqfAxSNZ2d0X5toSC+spmbDaeowGldk+63IKIlnbHng/rWyVVXGS5c+1HClCCXWYrjiR4
h7BZrYszNbj4C2QBSMbROhDQFhiqjhjIDM9NLXI7GMq+RwwSo4SgSHFBqrOdoYbc8SXEJPihSSod
/q7kYW4vkBaqn4VfICN/gsVIEWY7nLpHaGA7gaU0/ul5tGP6RFKMzxnYDWKHBkjZdD/8vjYYKMKW
pQMwPHCF+R/De5sceJZvV4INDinDMahvT/bmvwmItNPAwXNEhaSdGiqLRFp9es6E9OGcBQT8XvIe
/vqTZ5krh2xieK4qz3iVewC1SORdyIb7Y8f15DGgieJ9RQZ90hzN4XarVBHpYJ/G4hS0TOAR9I50
bpcqvWMmCTabFq5R6YG2h/rKGoAHd5/r2PAU7/oOszlc/l3NuU88q4kju3FKsthVQc3LvXDwTnIS
G+1AiKjFl9ROJ8lj8Q30GT6D36IkwSycdGye5RrKswoLStmLFei51u8/aOrf9JSk++z6H6owMFlC
CbaWv7n/GKGdS3ZWqE23um3WaQJhKRJu/fbDpaaTF740/Inr4rg6P+RrF8+OlGF26Vs/pk7PTCg2
+jYDOdEbFJS+ZriKAtuETMbG+WtVElE/ZHaFn7FYz8jVLQuIQBCav83Idksgrj8FuYxeOO1amujk
D2/frxC74Mlojup0N+r/ZHE2X/E7jH3EqvIEAbHURtvkN+8M6przBoavxiNT4oFAcDGSYoXbXSrq
Iu+rUPTASx9TcQYT+h5+y55uWhVkotoZqK/E4HisoKGxCo6yj0uC+wzmVcxnaa+bN7iAm7qspiFs
dfwRTGZaN0ikT4EoYl1mAVKQoGDPlVydhVO1TVst5oFclAOTMk6CZLDsqXXeU/qs79RdpmtBtgO0
Xic0zRcgOm8JS78tC3YeyQU+pH5zpYmiZUjKUWXnM0BlMCcKgDQurDvSyfQGzzQzFpRoV0oHU4GW
uLSZn1mP0YIBCPlgolPh3qiZD/90FMDo5m/MY+VRayKSQC3+dQ26wSbgW4+ZBGHoClFx0MCHJ06F
4PS/ZjThD+bs6/0QzUIOyzDgr8wEInqkCLH1zw9S0Ip/tVDJc8qdAnIt9ExvjfVbSS0fmj4RjWY/
h8RYfNwVwuoysW5PNYUhXkAdCpRtdv3mFbZYII/DQMYhDN/PcDQ9TXZ8S5CANTQsZjYCfe7xvqQg
Yu+ctSbVyG6Vx/KEG28Xn41Mlp+YuW+fBOPgnbtimarGEM/CMk34mYYuL79wJtmBqR2hLvmGIz8p
S3NBkjwJQE6NczNyYtPY0cs8PBBcCFqCmCzpPajpjL5+NgFlkaEDFyMn6Iz8RROuci82OdPkq3hp
v4S0Vo3Q8BEwv4/fVfp0nHyEqL0mrsqrO7YKmbWD0ov5zgl/E3Y0VDICxcQ4pGqMiQuetB2N4YNH
6vXwvgYdH6XKNsI+W7CFmictEBHaHeS2kh+WDjAk2hLUfFJsXVyQXAtFYGhyszvSjQTLdcIgdfpE
qXQz852aYkN7Bd0eiSs2bksNGdZIZkQKtnxm7sv4ONwXZx1gc7YwRvhNepWTihDnDyZNQsBWOyeG
eeXbRbb/b1pm9bpFfGzVYntMW5eZBb9F40CvuZqp13wE/dMeOKIZlOLN18TiWCzg/JXBNHlLkicJ
hBZ1m7nU1eU+/UuJROZFNplPbt/8L8T4rQfqsrW7FMEF9sDySTUNbY08eC9/8wqtWpjeVIcQ0cb1
RXnyipyGmr4OInoRisWRxflWcFW6mJNRYGt600XjJCP2hUtWCnFPaDFlSPIdxa4b/ujeGm8QsCqq
/TN1NxGjX3zh1yNXMcWdAznguOxnEoNYcm5ylzLVUVrXwDVTRnKLeKX1w9h0KRwBaDa7jTrFyFL7
9nCZd7yCGvvW8Gbx3gqn7aDktE2Cw9hNe6eb8WwoZ7cj+9CNR6PXGRINWnPbvpfM6/bhv+eZtjSH
Xijyr6lnlvFsTYfLdJtEV1oN0pss4lkUIjiovPxD1OQY8UzAK+Hi1w3ytfTU0RhOtIxOH2Isc43c
tFVGlsWTrqTLQulompUC2rlhLpOvdKJsAuRG/C5JU2GwigHHbPdT/dfEmJU9h+skTiYg4cPWTYm+
v6RJMeHOSSmbKktNrCedw3seAkT5oBvOklJYplfBKi9i/+gOhHlJzZm83C4j21vOMBa3liu+Ahok
szOLpYZF/3b217BAtU0zoqbh2aejTG0BAtDbp2J0kgEmHl57aGAbiaVeyvbG68uJfIj74qv7e+RJ
07qXV5wSZn6ZGiydTk+bzwcCKuOr4GlkhsNUWQ0SbZp4V7RVkhYFGIzhNvK/O+/EyAoZPSi0icP+
/clxg8n/psDngjgR99JahO4L4vFNpdzGePY1XgTEmeXfND2SQSkhRaRGDGHsicSq01gfqhGgcHRz
2EN4aTCgTrTIHzXEDj2+2THg2zAoxmBBRuX3ZXEAPDGqpHVqHFETq6VNsAzZbnuChr1I0YhHWaL4
exVzWGOFTfXezwoBruCGM3I/m1Dmm4JpAtrRHNvkkWGWMCVmm+duh1+vR0llOODVKd1wxpnnRUvz
c52AbzB80oaz4q1GIbYuqs43z/cReVr42oLNOSH8n3vSYn5S8xrhd8fXpTsk5/b5pUkfSvTqcTKN
tUkj3r19PV7Sj2X8c4yjxeb1XM+FgcEi5ACmcjjTHU+1/JRubyu/npsGqWiy21en4bWUpbOYk0TS
jpMi2a8bNwge+60uT8hWiMlrXtzNwjbqL04FrOZg5NUYizYaKrSCDS8BeyATKknVkc7c0DnzmwVh
1otyvTfOfAcD/a3xah9p9WdrmID90DvqDQCwc8M2dxJ73G+Tki/bARAe+w4YW6tJ5G2KwpwUJX3H
ALa0tRWL0oKteQ31BD+n2M/Jb6VsvCL4S+VFLkQiDQWX7ByjmBghvDu+MNbJFnm2BkCR4fSpGm77
RtFq/RiFT9HKpEQUb6Aw2l8uYIUCBvATcTX9OlCGSYda5syfYrUL6qwdPJ17B2JqrnqC5uZ1tTlv
Q8FROWerEvoW0OxZbEBJC2HXYEKdEo/SBiYHt6o191CGYatNjMfPFsEBFx4pM4GQHKqT0W9owBxC
gg+QlrCnGohpaY518i2ZHFTU3E9FeGI/Bdq/y8dPO0qI6Y1Ka2l32xEPRcsGbNZTUw2gfPvcucqn
JLCxY0zxLOaUOkj5NBTHRWyuZ7IbGotvFJFazDUR6R7H1AQCHe1bepZurgR9hy9nOo9hG350nLoR
2RGwFaiKjKKUZMdbAe0naL8JXpTb+CXBrjEyFvwNggsxWRwp8JlX1klDhFy+nxig9PfmDFB0Vlaq
SqUcyAI4gRxuXcvhYYL7Yk5ShhXXh7EsMgsTevIECn4v8BXU6tNmKcEgQ6QHUDRQGsnVEG8Z075f
V7cJw70ILE65FSy1QzuhHUbFukUnMzE3qu9XrxTj3fsEvvejRFFuBW4VZMvQb7p+MfeQx3OWJ3c4
9KXDbvOGNzjIHFSVJ/26ixRHlbVoqQNuZnIMkZQkjZ9dswMXpXi5hEPloJuCJLPdgRNXndWjraLP
VUu4Yvzzezb6b3m5xDHz0RV1rAnq91v5dhXWu8sucLt8ix2NIqY9HGd7vSJYYCcOvqiUBu+WnZEz
0Tt59wxjTCx6/xDc3qt3SYXnp7VUEjsJmuhQqmh+4eRgPlVK01wS9yr7AF+marpOc+iwt0TVDn4B
xtm9XzZNmHa47ewt/Nux+0a60gawRMekl9D+CDmfpT8HleenGzV4RLf/9yAp70DQ7bLV9lBTSnVF
Agu0Ze4xo74wovDO6wjnohGBAGghAXLN6kzdIaGsi5qa2+9aVNkGHSupQXt79ZstRNFHiAQbCQBI
NY6veJS5yAkanVNymreTzUZwhPjnEMNr+CCHyJ6GlAaso9OX9ZHAEEopd0WdCOwFjOMWwYbUnjcf
mRcqqxCpqU4mah8QcEJhNJC2x88PbekExywoBunPDUPJ8e65f768aM2E4XcdmBdK0n1LxT5ScRe8
OvPSTFHa9+w8iZ5PzPe300GfdCk1+/hyjh0JtxZVyttmVhBmFkJ3JvP59n218RiaRUAUK4D/S6fr
RdqYTum2IId7N/dgAjUtq8wKairtREUcQy0mDvW8WhgzSwV4jJCmc7tk81bJKrae5Ywtxcp/vlbh
RVbYiCc47nXihh/oab8/JnGDK4yQmQmNNwWyNPEc2bcilDdfwb/63Ib/OUnr5qjCGN5Ba1N3z9ns
i8R21WeD+FZvLT2p9RFdrDhUabssAAIwWlZLURXwja8EPc8Z+1bnNKyfQ/ixvn39umef8ZWbNa31
Ju29ywRskPdNqL+rJRUbHsPvQfAXmD4ssRQlWx3P3xJjMjn0p4ObPA2/ux6LUrEvLQpjAZ6bBr1A
OeiX+CjaJDox7nL2S01OS0HRNT3wbDZ7yZ6Ja+52u8W6q7tI2oThMQvcpLNkRuOCcbGhB7473Ddx
tXVxiKCHHdOb/BErKAu6j94DXcjqW4CuIo01Kwc2DyW4vbo8rAPkEsnDETlihGYXM7wWFzYF+C53
EgEFArVC5GB+pa+OjUlXHGEBDHi7XWRJ/B8LCkjS1zd2ejt0DrXtUcYQTt7g6zyHSgDQOraPa7V+
ac8FwBRywH4YVdVZ9xoWKg7ZbGQXmXqbgBJAbklMQqrfbeLI6XlTwOCk4wsL3Ro2yPx438wg6ATJ
zAD/xouhX7l9ohv5V5NdU6/YPErfWtclpwB7NagSolRdAL9ndbCn+6csxisnUi6HFoV+eopQUb7H
q3jRll5tn+jRkBX0DCcesu56OUK614Wian+yYmzQtx/jMvVyZs/Xhv4vSjxOt35Q/5CKFKbLwtXD
IKP9GeGMoXrzvUgis37lUXTF//qJKq+yo22oAnNthYnsbBVG2yW5UhebbKksGrPyXjb1AWA00RWr
9ghbSk/c/ZHeSwI6UHhfQSf5KBcQCAOyatbtpv/+vy26vmTxL7QhziIS8iwudSEc+eBfybEoz2Dh
at3XRtzVgAAhZeEbuciU1zqY+KeGDYqk8cYeMh5o0Fg+9JYFCLWoVPPme1lc1CDR2UPa6hfKaymR
I9zjqwAzQhNg0BbmgZ/OzZ6A8EGuxF2FEN7Ci0ECZsdCyyDFn73zOQNS+srJA9tDEPgYNtukYJo6
Y780gTq5LvyJZyUygDqTKFkB2VPdwO4skCVNOjrQomk9poSWwuVEehL3GyfCx8EizrNDmGbhCBuI
NLZJ4f1IeO3k2aUvXDrpYfDJQiW4w34ULzXfL9PMg4hLv8OSzWEBeA3bi0Hy2aXCdspR0Nh+HDjq
CUgA3So849WIX8Zj/6MMTEtPbs0quG/O94m6aJBunpRGmo+Lwj5p78vTvFHuS+C7NJlubjO0+jq9
H42yNxkFPjBXET+RcskbLUO0/zGuGGENqybwngJ71nGYx6jCgncxEBbHKNjQDKckW2kht2ZNsefb
V+2V4TKm0FQafutmnhe4tJvRk+aDUFmW5FE/hQkDxHmgxf11FLmfAOByEGD439YSWz8EcFkAKUVm
/rXKxTiIv+qMAN4r4mDapc7Sfq2nO5Gv8JA6qBQVbz2qOWOPnMLaBeKDhw96euNqdPE0DLI9yCFv
LHeTB/I/HRGt1z5CCurQq/+Rj2dEAe5Zf/nkEs1BeUK60gp0M8EVuiq5NTQHkIswJXbKObNmBYM0
tKuE/+/zE+4UDW+xZxnWvnPBKhjJw92LylNn4Tli+b9WiLDX634shlMxThIeyKFj1Kef5t6k+9G/
Suuh4YVRXoprpozYRKD9hah7GLXTNEP2kP9eBU65ZG2CIpDWMMQUIGnbNFGuPbB0SRiN6ZLPabQO
PpB2qNJ43JYlqkQcc5hHJgPIJnxHqb5QA1/eoL6/zzBmQY8axy3xLn3XjlWvD4LSui2SfLMNS7OH
R8tsSsI9C3vqzHMbVHQb4h76y087RIjlEeAfZQRCrJRnrndeUg3GiOPBawmFa8lgdh3WOuPqAEEs
HuRoyJgsiYU3DaCOLMZO+gay5pNG7q9LHZjBDoAV7aan2l07G+45KZBFjGOfbP1x2UI1//cV71DK
g/zC2my/tV8/AWMfvmyC4IMIho8gUAxRvwEW/3vMaJcIfXkOiLcQ9GflmPPXqPsQN61u1bSTxed2
11xTeYFEwGOeQ1AbMorxMHV/OCN53uYFvF3y2Zj+ozmrpNbF7nF3bHDd98xB8fzkhb2wNVVI48QN
v/xMd2CPZOvkf+IJOsCOaoPQ/SXfROw0ziBkIBkBEXK48ekNtT+nVbepl+AhIuxcd0FPs9qHVz/Q
Y7CGqTesV1lXAz2sqvIlWv9IDCZIQdThq9nBckCx2U3y4lJ4/PRXT7FHnfJQ884KwbhJTXkXCBcT
GwcxD+cSH+exp/Zs8Llh7ZLIXvJQxS4dCMaHRkggvdWhq8yOKnrwGbaIZABpIp6lf59HREsuKYZC
AqPBCVrgXsb446TynPkqS4EZ3hd8UWNrGAMS0cm9KNe5MuBu0/wPszE9GjdgTfTqMmifHFJkAiuf
q9Q06FiZw0aJrbbU4dioyRz3B8SMCtk/xIycZGlU5yRtk38DT7tnkccZsHHhyZoxwgcDHTY1/ArM
oRgcFnuJVmE2Eo8a4fg2YUjgBtruoGNNnx6kr4NoKJrcVDaIvsvNFYuCnhNv6uXhyqlwnthYdLAE
4wpkrjbXiU/vaFQF9PR6oU7IWFr4MYqHRsJ3i4OS0XpqDNx8sEin0QwCeWrrZxRW0AO5mEE4kMAL
SfT0ppK9jUaU1RjMpNGItsHfJW5pBIETywx/mWxYLwf9IIZiNzzaYo+5iOl1Fxsm2J0Aos2NtFB5
EHN9aBFds/LygMcN/geBopYjrDhgTtUqgLRk3J+qKoh+f7I26neIlCsAcSP37kRDMdaFWspS06GR
mCgdPLGmKAc90m9VABWwt0LQafp+3vswEmQYnAkzo736C46jfUPW6FyIkgAYsEId2hYy4zSyMxE7
9bCPFt6IUEpFaJvCNjWC5sOG0od1MYqXPgl/hTJk+haNgOPR13EsSu+bUtV7mRCsRcpihpCr1+7/
lhZdE1soI6wDizp33uqVzDVliFS+osCd+MehoIUtESzTo6/0QibvWI50FiJi/UPfUpZChxQVrLm6
5nkACG9wsBZIS54doLeA7nzzM5fcDiz0nlmZMB9TCWtRw74g/5VABRxIhWiREKhWHrN5OwFXnBCN
YIRrRw89wCS39jlz8kL2smwonwXpwvDY434A4NCLiwNlvvFzZXbORZIKxwF2A/7p2QXfjaxt70wA
b3kB6Yca3P22qHzsKqJQI9/fYNpgE8QotykDX80e6bJts2JrK5stqmjQ1apcMei1vwY5ZclIHK9o
ru8UaSC6HNJE0PLg/Gau4EeO408CCGpSksqhyXSk3QUTIEQLwSr5IiyZiOPg8K9uP1A/u8ByxeYu
KCJUsoYSqQk6ayy+Vx5HtU3w7N8YqbEXOGHICZkhXdGZXNhCevqVC/6J1WQngE09DTCHwgrzjggF
kDdpWcJFqMEAYfbK9dLcw8gv5FyDxUbMBT76lsOz8kf4fBrv/2O5BKZKwBR3bvjS1jZAMZrPAhU4
h96lq8tutFYH9drFiGRWH3iQX4Qnq3s4i75EYPbDv53gKmzpodFoamr8fXXsJOLvJf9PcRoRZayX
FDzAe4PXHCCauAyMktR6dNelMNgLOEIa8MieRnwLbRkQzDV5V4v/9oei/zoSPVUozV1aKNmy+jSX
kzhsly1PnzJxw3M7aINLaUcyaJBla6tK5jpR9IwzUvmqKWbSWqPiWC4t09cPF/cowYgi4rMz5co2
cDju8XeyAEYv/+BbeTIgIvBo2eEgRDS/TPR+RKGY4eBFZDJNeXy1dME294AwJDCA8DMmJvPI+1f5
6XD2gKPVPMTG2sphorEIelSgOO1ARnBGxZmWWoEh+VZ+SvcR/ppDn7m/bGHE4ip6wURlFy7mfxJy
EUklEKAGjdbVOjgzrBnf5nSCX4LtneY755kseiixRLkqOv9ci4UbZJO5nFbHPP8TB6i8cGVPfRuc
88pgubeAERtBphCV4YNRknypMg/dW0gTjrN/eqZHOZAruQreiG8IAEO27x1XNoK+NH4yIniOnd5J
qxio7A1kSbqEt3akWfocLC+q3J4ftKIgNwD87Zr5on8fZnp+QTZXfvRM14ZBxJhFWHlvN96DGIcE
Ubvv2XLLNWsfBPa9s6S/0/mOeGVsq2KM7w9oXBQr9KB8Psd9lT22Qo1CpSPqZg4lEBtCA4aj50nK
/P8C0qEQmuuDdILot8DPe6HEYNilLChAUayF4HzcglympHO3CB1T5OwzTq4BcqdsHzo+ELrZsWOD
YJDJr5OOD1dn6SixbZEfyDoVSKGZq0Go8ym4sDUqpwGSGLJOhKWzhbuC4NAxAr/ZpZSJfUnZJxhx
UsKaKciWyfv3CPmRNWa6jmjnho9/8QjixW++4tPRNVxXhMsonr4lz10SsTo91yA1gar4myqnZd0z
ZS8WzGG0LQ4fuXjg131Giit2ht6QDgk1ZSbKkU1d/hPsQC/VrsNq6JbFavlf0IYFFuFKJTQDbvRW
KlH7kM8hXX9oUopHkvxEEGhmPaaSRrRwjzlhqiQ9BQWiSv3efTUYqVnUb0KNF5/8s5341jyg2EIC
jYXvOCOx/KD0ESTH2slfoshi6f8tHAoz/yCIXsQ6CzxqUuXdtCVg788tPTzBVGn+Mlp+LmHc9Aqu
eUgKhn6Fm8O7cDBy+IEGKaOUPpTcsMwnRj+hR6pF+cJJOmRfXmjt66Nhsc1EpGWYSGXa52cHr/c+
hMR65zXSKouwBeBDRq2ndRCg+x0Vnf5j/C/Q8RbihfkZ5jEJAGHbJWKbnLYGGeoZTSdFVeIIkplN
6bCinjXU7RKOIBL/cgrhylCzcxXLPAuEzaj8OqFI6gBDTqqw5jEo12inxqm6kN7DpAEF4EiQQ8Ug
ABtPSQCX5IJNBJVDp3sllkEDuvkMBD9+7E28GCoc4nG2RudqzYv15ztVGkoSX8goNTwfMVTnQ1kl
Y0MP67nc+ME/Ywerd4BmBvXn514M48To3O2XMRwzUDtCRrwZZBa4Kre5QM8ils8QsvS9xWGbTboB
0JRKduhLBzt1sZykCFs4NrEPy0f4MdySN7zcnT8UfTctvnNLox7GugXYEnl4NAmI+aMtr5MRIfFp
rU4O6ZZKvDxekeybAoBHsk28pE7eVqW0nGi2BTOqslROGkfHWZIjK9pg8fhq2jtfCcd9Emj8pAFS
vIYyPuwEVNoTYNb10BhT2rANJqI6FK0aWx7QwTFKHauQeH/wc8SzyKHRWMsqr8mYcpc+HqfH1HO5
V5WZVvXCE/zoz0XZvojBWrhLxepdEqxSay6tZ2VTX7wIOp6SKTO+Xc2+B7gVCdw4OkGs66UpQ4DL
q26bGp7nLb4nwh9HW3r8fN38KojTLnKs9DEwv8RwGv+VzwEj6kuRH1kvZBkZcwP9ZRNxA+1rj4R+
4ZRaY8tMjxUHZRZXSHWkob8tT6jtNhXVKVMD34EPDjfrJvytMpXZobD/LUjlhmIypiLEiB6YMXZ7
WXaqCRUBjEXcq241wX+9wSE1Orm+zkGvTzWAbHgqi3uSFb7lSgZrCNRkRyZFIiSFRbBjiVldeLxi
V5wRB9/mCymCwSe2SlPDIljeunYx7/ODy9f5oAJU0Wsg2zJd1rACvsFNEF7S/UKXa/5K7YNG8RW0
p4PogjRk/3tlwRNWxAjNE0Rz6zCS8BQDExE1DUMW3nWzIqp0l4ejBAf6EnuOANSbUhoIEK8jfN+D
8EejEcgosuAGnog4J6JhI2GJUV78yU+6eKG1L/UW9+yzudiy7WHLUoGljgku2dSFf3L5QxyIinsM
QnPaUR8YxS4IkLt5esetQZAv3/t7ZH+6TMloGY3ASOHG4/FBB8/Qp7ElNw4VIqNqHNLm5y0z5KH0
zBD/9GnAtOGQr5A6/mCPt/CMRLcu0glU9zebVWyQQmQqdGOYBqOX6Y1a5yoZwyQN0jAfO8uYnHCL
gFPYGT9ZFGwlxGfRuUzYr5UIvgxiyi8jDIjo0kEOeHi0Du+TJ1iydXA8buKyBMCAXQzw/vYbeJ8Q
ztPSEOsPsUwk30y/EVCYbZ+a9rbMYwNVGg7IS0Si7pSNA9S9yPE2OM6tTGWXVLZ0UcI62V/T1RJh
YbTP5Okz6NfYngMhy589414kXjahd4RHOABo5m7ReXBvmiPwCY5fAVLp/NiFYoPx6wYeTbFl21GE
dnTreiPKxxEX9R5rDwv4bCMtVPFTXJs+jpdDbn9gqilXy8CFF0vXudzF+FR4b/45HlJiMldRRLlX
6HVggpoplYhMOsw7ltFB+8Neast1hesgVqzKoNDtCj6YZ8BSfvwLLZke7HnC7KsVa3fgpPT3kNCP
W9TeaAmP9BeqpPPFeitmOXK3/s8qbiIkTHFg6Sth/bQ8ubWyrKFenrEt1phAhjefVkK2w4QV8hQ4
3XYI6/6p6d83kHfu/W4hesSOZfyXi6w+OZ3HZIveGKGqU/dyabuB8pswVe473iS1IkI0uoywqT5s
UuK+Z+KcULHXeH3I5fQjshwbqQCpg4d+EcAwf0uAdjj6aenpqSWspiXNI5HpRgXG8nMglLrqBXsi
7OFEXGOwOB95P7o2wAbGHYmynK7hnp6iekY4g/9nM48Oy+EF+of+T+8vBYoM2rTsxGtdQDdkGqBf
dTzl+XjwTnh8mhbQ0D56l9HfomuKIDwcqH5RLcJv8BWvwhNayXYVq+9dsoYrguGtTHQy+QQg00Zs
19mO1x97vdGuV/6BXZlEtY5xjl7gArRxyqXz1G/swsFnSRSK1elpvAQZRn1HPjkIxtl80eu2EPBn
Ddl/eqLI
`pragma protect end_protected
