`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
iQbEix3JHZTwa1vhipHlmwS1/G9xw/soq5c1aH9r1Ikmd5PFC6vG8hcczrO5Gm238/UZKbDRHhQl
8vxxX1eWXA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NYO2r/VW0Uk9iILO9avt3Skw+TFdXKrXeDrkjkY6MrmMZXqmt1ljuTdXla3Px6GiDC5iNRfSB1LJ
jlz9x6ZyMo5VxrDlXmNLima4xlcLjwQ5Ldngl558uz/vr1FbORoJ+gk4f03PWwyf42EKOYFnCVfd
LJfFRdBml66XWTkIRRs=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hXM/negBdYIePK99VNL4dA9qZWSDCbIcZGIF+wzwJF2GeTdZiC6Sv8N9/cF1YoJ4PmeE+1cpGoYE
hr+rxDAb1wjgZvfDyEG1QWzKRSG5E+oNC6Bj2Xk8erPPxuHL0sXJnNFmZt3mRdMMjzJ/oBGkUF0h
iYE6DHIS9BMznThGr4tm6wOQ24nLfv2CkGw5FtsfpBEceglyVNwc5KmDZpqUutO1UmcXWgUVf6aG
3t7duiHDJKzCaRYGI47UkrEGgYTLtr4N4clyKbc4ZaAFsMfafXuq7UodHyHPGa7sQYA60+7yMSq7
lZ6oowJsQLQdpXSegbc7gK8ezWVXMGToMCUX4g==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
IZkumnZp/JsuGCxK7A5f04eL3wOhVC/HIkiq9ThWDUN6/jAV9gkhdECfPCdAYxhe0IfGI1mwNrRJ
CATeVriO+TbtGJF8trisSNtrtJxyu7w+ARrQ3i7xJ5OugSeDn5jrGtPVCeIVbs8Otz0RthJD/ia+
zMRiRhN8wPr8+wtwChbS7LbmoKzd361OLqaC8TX6Ab1GBUHFOMfYyAPJdl/jXbS9u43VHuRY6Yc6
WqrfDJE3842973TEArl3DaaLzZwM28WBp6JNk4Z1zR+7/fPjneoZl3Dvksdx4ThM0a5s9BNPAH9V
WF7gF4b9Me6TfP8DfbNOy0URIYx+xbfpe++9uQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eaRvVH2iXg+bRFhfU/Zdu0OhZxAtLuP0NVIWmdEUooi3G/jC4AtcmpPrp7p/DrHH2FZwIvu+AbK3
sY3ybtP3ICKGUwlnIt7XryFabcZX+wxEJ33rwyvMH3qSJUvv0NnXC8IHlKKyRjDylY/oANDzbz6D
+mWDv16FdHx/0RgRk2HTfCPx8qBZ+fT4hbE6exCfOH2KzbFjubsbEmNkNU+HUDcusYXP2EoAnNGO
lFufKr3GhljOMYxxaVeKpXEcKWjQB5Uu1M3JdONHHSUP3iVPekneDcajTRMfHD9FJggiLA6mAgel
cdhHqUxScYsWsL7cenQphjXngVDIxqnSMZgGGg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
heQDXwsWtguDyBBqy+N/Xr88McxL4tQSR2XBCb/lxs8IKaambMExKMCiF+uYl01VHmTIU2W66UkM
7t9z8H1Gdw289KkEy+LLNQNFvy4xiQp3che0cCrsbm5/JjwMeuGavzmF6wwMkz5sW4oMgRBAsxzn
RRGXDS1r2TiNXhNi68I=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WZqwWujfHGXV7wBEePMjGLVWUeV/ygCmf158CXpAhJC77z2vuuagSDsOpGgtqyakG2cswti5bhBy
iGqPgNkEY7Q4T3NMe5WssA5nf18Sw3LU1MCehsK5WrHeKiMOyz9QpdgScXEE86/e3qniqvFlM2/c
HpI+I2e/HN1QOgChXb7HzAEEqCCdY9VD1a+p15IoOmU/8Gs718QdaPMJOt3XdTu5pAmq/PWuICaZ
VFSPDj57xVELte/pDBIXo8hgI5sad9ci34UyXovDzhRyUKzLY0u+gqRalObdZFD1Ph6hGQiLfmwO
JTvUCIjoFwTzhh0dCXYGcwc8O9kaaOIiiwpgyg==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
B4GVIi6TGeAAKF2mV42cg9jGmUkeJ9TkEGN3HtEus1MF1Zmt7Nh1Y005XEEzr57ufgLlM872beae
bxX2U/dQHyW4OCP8KBTn49Kmkdu8j6t5b8W5HRsXXHYSGPOo9IxUSHBdhwxHpNWauRDmTFNl2lia
Ton0toY2wVDxIcyINRYIpxD8YGHOnHSHPMsgAGtuP7kRvUnSvNzqqhzVcNm3oeIMTawuhFgBXD+f
0S45sDt4HAERXJfO2RXmlDCCLpg7FQxibRHwoppbdhT48SpFRar2SU9FLaP1Rhu4f8UN/BXG8JDH
IE70hcE1uVmlqXL3h64Aaql7Kf0Mt19/bANOBQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3328)
`pragma protect data_block
8fgGNC4HfskTXIPOSZDcR0DhA1/xPSvMbOj8bNtDga7qhlRYO5M5dr3t8SjJxZGOJLc9YiMFCVdG
c8TKUF5fx5x3s+O7VteTbupS0RQ3vzB5laDxXb6+ECJh7oUlqmG52lrE15VCKKZrRgfNmk/HV7rk
uZJBmzcpDb68SVT20PbDG214f8pQUnQDhKduWvzGqXLOepaX9MoQSXHOs/FxZBwPj6hOjOS1CFcD
R7ZhdwDng5t8CyAmYKD7GK2UvY/hwn12NdY93GEJ15QB1gfHA4HCNJz0yMtfT+lkWm4iGjB78mq8
E6msAKKFHuc4WnhL29tEtr3mR9yejcSTV/t0EBjqD+ghjZiqiFx7SzVmbh6ImtK2m8OTlv6dlgUr
PkkPl6A7nDy754etBwLHDOxVCIHzGNiNOk8wsSpEco8cZKmlmS9mgwlbqmXyDCiRfjYVhAoL5150
Qdz8iheWNmTvR4mH9yUmcOqLQ7UAS94dENLkoVTeLgsXshbZWidd9rrpYigCJk38RhAsgPEOXaMM
mOV+eUZtEP1UufE0N4DX1u7hAzT8YQaODHrqNPHDu8mHpWGOvySd5/v/eLEaJWrW6Wz3NhQEqw2d
RxjiRGEHlNJWgn65gvQJHM95vROhobZ/AIBGrmjOW7DX8RLibThFfg5BXHKOW3wst+5ZcdslAzKh
5Q+KDf1TI7O/ZC5gCTe7MiZUZ5YMe784I+Fa/R3t8bATFKbEr4HTmqVPkjIafuip4maqCaSg4Gnp
adzuCMwHfl69couMDW2EtmM1aKD7HPLah1wbWsqSP1E7ZCmSF6gZ4ijR/PWTTp53pHCeCO4cuw0/
C+TDnbL9ZS6x4i3lbe+95Ixymrw7PDflq2F4js+mA/jBQ8ys9Z4bXFynLM3Fh6r4x148hl0G+15o
aF1P3o7rba5sraLYslTHyU6GkwASzb8mY06LicIbMRy8WYBe8AHCzcUkIuyNzFqwLPQjq6boKWCC
K+VOqKBDNMfzTaupQHyo0meJjuzlL3z2fi0QVvCGj+4dLgPT6XFtZtyv6Xka2GePh5iXrJoBYwhc
uQ70FP14PXQS//QrrTnIxPhZsFixBfRqrUDoEXas0XvquL7QLLafAND35NJTAzZKmm18DfvYyezD
JND/D4Zgn5yRUqAn/zhT+11Z3T7bpxMcqI5m3fjr+zj2CvykKTQokgjq0/75GPQOf8apkqhT/bso
Ny7I6Lqr3zOwHkgyvvW7ORxoU2njQjAg69BwCQnsgYW7Y6t4lsevGpaj2mfK9U4n12+yZkSl6Am7
rIBCS7liuiffQnvcbjU8pEvkyKZuRMLNRUjmm293TWyOFBFYJv+jF5DV+N4Vjo+FRMcIXxK1nroj
en4+08+iGyTtEHHPNySfPvzsaBcerAahFm0+uS6qu2pIdz6bwMKyWFS/uuI14Ex0QNi8+9GQgRJ+
p+vetJQY/SA8GTG9UDhdemXf+XQMMbAtyWWskekDEAsaX/RHTIne8DcOZVclkTrqX2k3kAo/0BAG
kFe+1Cs+0CHy4h8I+2Lgx3nLIJo5HBCvpuEtbZkMcnaKnoXSBtxxqWC3rXjpfS+J7DUmslPIrtk0
egubVaKZ0UC2JCWg8nxAWDJiCjr6PE9B3TErFVT2eJCttltjVupkrMIej78iL16xHEadMx93FrTl
y52qu9ElpkIo4xGcDAPHzszIiCfR9L01Miu/ru4Jg+pXELrqPAxw9oYtW5eCXClLwOf2SCYESsx+
v/99cGXNSS4DfHSPV3koXGf+HC026Vzp8jJ8hVJsN7hrR/9KoXGYLPJvGzQeujSk5JPqZiPaQna+
1oTCPHxv5dtumUAEp2q67YKx9QUx1Xlga2DgxFk4hDXpdgnJXcdXzEU3E7kFZNyij9/oL3Pa/yc/
54zE7hUW/2BkfJwA9+aZbL5o62FjOfgvt3PrpEbk9DQFbVPsIaK61W2lA6cPF2KVg3/k9QBSTmxL
F0JSM9lqXX/A5HlR5pIl8ho8cGhwNig9X12PCzjsEDMjv+Nnrg1X9/397A9am8MBYLSZSwQhTwAz
Kbk5AyonxFyvjxuSrXauYoXzBK/AlzT6Hv3u11pJqiGwC+EwgoQMXR35r0/ZrRQ5fVT6Iv9DZR+l
Y/3tBrcCYPsLHb1WBTn8J9gswitlrT8McUpdTsETVriz/oZXJu6OuLiIzfLYzVHmZys4ZQhvmJI9
udngUsis9KIr+Kud9c9lwW0SU4LhNJoS/y07Uus4/O8f1USacHhCXeFM3k+gymxg9FWZyU0G1dyO
xrwTe3xFju9xQ3CRiJ29jbUnJL0FYrBm2PysIAsQR9KvisSjqTXREdg0qNee63+bG+Jkenl0wKDI
8US0vue+foUsAu6nAsOI6/G5lRCTBuQytKw6MSvSP8Q5hXlIaC/TJdYWArzxrv6VXsAF/kq4Vx7Z
XGn9op2OI+hHeUhnb3fliunpvAh5mYQkMIsSXLw6y26mICGfGDBTwX4j2nKQZ9MP+ABPfiU4irXf
mt3jxPGYoGsHhC3bBtqC9+l4p6yVkdUk5JAkBfDmRUGKmwsVQSV5vtgDz9bhYWDuXVHinw3Y21lK
DmGLz7Hc1zMbVIh0Fp8YFXY+gobjEvmIVrZK9u7ZifYVq8XOhMUbwNtRiFatgSChTEHhQtpDcrfs
Mvl0Ea5fAUTpFBy8e7pDdOb8I9lcN1BFyDNvEFFJTk7HUNBN6mViYaHJrsdhy97usyeTpZHQWZgU
oy2gws4edC57sKes7HEmG/9f1Nv9FTIA8Zfv7bc8SAi4Ej28qOUxn6zcOTuARUDNtddtm3abUP1p
BpfhZmpHqfXGl5rD6sSrYjocBD94R4TINAwKmnJTNoxkDW2aUD/95M0Zit1N0ew7bPM2INDaNNAq
rIwe84phu2z+yYWX5Qp6/f0/rVltCs+WPM9V3b6inE4GOKF76KUxGmxQKFGMI8O33lFzpPipLPaN
XZwDjyjNGDZOOl9PXIZYn9kF48FGER1uzQc1nScZXDjQR1eFxkfoHqVORJhlYYDQe86iqfj0k2je
dzJjpwEFMTpwfEuqDDMYVWGbMxL7n6ErY2Evqyq2k90Lb+HnmUov3z8L4ctE/kDnscN6WX6fRkuZ
kAiPEyYr5CodEOM1qhw0S3ft1wvwXWEy2X4j72q3LPZw8quSN2Z6N0nAjRyab0FUi31tZHepyLa0
GdNruMt8Z/ruc+fAI2Q85YCRbb9I7yBjdKazSWiZtmPCbkLRG8HXaw7jppUePXxGuGElgm8cRr7P
TUFBH3fLgA1YyEg7aZPilGYahFXDxNQOiFjbdP89IinCYXdeGwG7bJfv9ko4DXFDNygCBl0NwTVt
fMzEi7vMc3qz0DEgs9VKIJJpB5IhEJJNyLirblTK0LdoM9me5s9W0oOa2bwu3s7/tmAYt31+09/h
g4H26N2evs9OAIkAKNZXy2mVzWRL3i8jHN2nyeccv7KsWJnU/WZ3XutMlzMDz8KEpNozAc8ylk5k
c9YzS4twJY5MeT+RduU6bvqDb4CACJkY8BED9ixPGNamuAGikF1pqpIdOjfWVqhcVHfJpFvthvFH
+z5hMGdr7QulUb3Z4LK9YjjP5iECfrG/bfiEpEu4sYC++S7qDSuPcuEmTVO7DtTxKOLGt5ew2G0l
8U80UAtGZhinXyIY2HQ6V4A6ejgBB7ZpQwCwqEmPe5aY92P2k52rMQ0wIJ/D9oiBRvGdGTUcrlSG
gH1Zw1N0SxBsENdcitMZf0/ZsfUtj03UcCIBnbGgy554unU9r6X2GzIadAYyXE6jmcRKirt/zS2n
EM9EOsX6/UGtZ4P+yk1/ILQ80bdXMPftpqMj5e6GDQBRGJLJx3nTv+yV3AsFijReuFYSoem0HAVo
JgF+gmm+q3XT84YniXv+rXvamxTnk2CTV5fBX5JtBR4vx4dnf6uV6KQPhkrAusNRc1VWbBabCO+o
NMO6jjfm43fALu3rDulv8LHtHDehwSCxnPMLZ27pAlfxL6GHC9nTSJX3tldR9fdwRBfKIfSIyj6n
xfq7VKaZWYXQNqS3n3Zf9zJIZqQ+L+m8EN8x5XbEvOeMWz6QMf6OG8YyfiVH+NEGybU0anxHr94w
vA4j3vxVaYEfUta0WeRBZCIu9QkTuK3bTEkd9aEeewjozzrC+hl1EX42jUAWyjaCIvtulUYqk3UY
ST9YoEBGAZz06jOUQqT2hI5w34kU2DJoWUBWcZLA9HNjb7BbS/43jmbUffUK5GYMURhd2RGZemGd
Y8EfN8bQJ3tFPtZmsBgW/vH8RP/os4OLdBE2qy+sjm3UihYBLdiLROcyvXfY3Lz3Z6SPFnCs8jGd
o5j57VmQkyFu/Jt9rra1Hg5VKiTSY++MLk3A73vfxblUQyXB6faWoGpZXgHQsWe0WEKJd58T++hP
47R5e/0K7fkOVGFk0dLcZen0ko97Bw==
`pragma protect end_protected
