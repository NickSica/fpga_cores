    .INIT_00(256'h0000002fb1809c0800000006b2009d080000000b21809e0800000014b0009f08),
    .INIT_01(256'h00000020a5500ce00000000b92d2063b0000000b82c00cd0000000001502063b),
    .INIT_02(256'h0000000ba252066100000001b002063b00000020a7f00cf000000020a612063b),
    .INIT_03(256'h00000014a00224920000000ba262085e00000014b003640000000014a0e19201),
    .INIT_04(256'h00000014a00206b800000014b002069f00000014a003649300000014b001d050),
    .INIT_05(256'h0000002f21b20663000000062b0364910000000b21b1d02000000014b0009006),
    .INIT_06(256'h00000014b002062000000014a003a49100000014b002065100000014a0001202),
    .INIT_07(256'h00000014b002062000000014a002fb1300000014b002062000000014a0020620),
    .INIT_08(256'h00000014a00364590000000ba270d04000000014b000900200000014a0020620),
    .INIT_09(256'h00000014a003245900000014b001fb0000000014a001da0000000014b0003b03),
    .INIT_0A(256'h0000002fb1a1da8000000006b20324590000000b21a1fb0000000014b001da20),
    .INIT_0B(256'h00000020a551fb000000000b92f1daa00000000b82e32459000000001401fb00),
    .INIT_0C(256'h0000000ba253245900000001b001fb0000000020a7f1dac000000020a6132459),
    .INIT_0D(256'h00000014a001da200000000ba263245900000014b001fb0000000014a0e1dae0),
    .INIT_0E(256'h00000014a001fb0100000014b001da8000000014a003245900000014b001fb01),
    .INIT_0F(256'h0000002f21d32459000000062b01fb010000000b21d1daa000000014b0032459),
    .INIT_10(256'h00000014b001da0000000014a003245900000014b001fb0100000014a001dac0),
    .INIT_11(256'h00000014b001fb0200000014a001da2000000014b003245900000014a001fb02),
    .INIT_12(256'h00000014a00324590000000ba271fb0200000014b001da8000000014a0032459),
    .INIT_13(256'h00000014a001dac000000014b003245900000014a001fb0200000014b001daa0),
    .INIT_14(256'h0000002fb1c1fb0300000006b201da000000000b21c3245900000014b001fb02),
    .INIT_15(256'h0000000d1ff3245900000001b001fb0300000001a001dae00000002500032459),
    .INIT_16(256'h0000000d9ff0b01300000014a002088a0000000d8ff2066100000014a0022491),
    .INIT_17(256'h0000002fb253246900000014b001d0010000000daff3246400000014a001d000),
    .INIT_18(256'h0000000d1ff3247b00000001a001d0030000000020032471000000250001d002),
    .INIT_19(256'h00000014a04208e500000014a04208ba00000014a04001b000000014a00000a0),
    .INIT_1A(256'h00000014a04207a200000014a042085800000014a04207a200000014a0422486),
    .INIT_1B(256'h000000062b0208e500000020a72208ba000000022a0001b000000014a04000a0),
    .INIT_1C(256'h00000000b90207a200000000a802085800000025000207a20000002f22622486),
    .INIT_1D(256'h00000014b00001b000000014a06000a000000014b00207a200000014a0620858),
    .INIT_1E(256'h00000014b00207a200000014a062248600000014b00208e500000014a06208ba),
    .INIT_1F(256'h00000000210207a2000000250002085800000014b00207a200000014a0620858),
    .INIT_20(256'h000000032aa001b000000001b00000a000000001a00207a20000000038020858),
    .INIT_21(256'h0000000d3ff00cf000000014a0000bc00000000d2ff208e500000003301208ba),
    .INIT_22(256'h0000000021000cd000000014b082063b0000000daff00ce000000014a002063b),
    .INIT_23(256'h000000033022085e000000032cc2063b00000001a0000cb0000000003802063b),
    .INIT_24(256'h00000014a002200a0000000d3ff2071600000014a00206610000000d2ff22491),
    .INIT_25(256'h0000000038020076000000002102006d00000014b08206610000000daff2069d),
    .INIT_26(256'h0000000d2ff2007f00000003304324a0000000032f01d00200000001a000b002),
    .INIT_27(256'h0000000daff2008800000014a00324a00000000d3ff1d00300000014a000b002),
    .INIT_28(256'h000000370012071600000025000206d50000002fb270100200000014b082085e),
    .INIT_29(256'h0000000b40e200760000000b30d2006d0000000b20c2066100000020b8b2200a),
    .INIT_2A(256'h0000001450e2007f00000003403324b0000000005401d0020000000ba0f0b002),
    .INIT_2B(256'h000000007a02008800000003607324b0000000006a01d0030000001450e0b002),
    .INIT_2C(256'h0000001470e010010000001470e2f01e0000001470e010000000001470e2085e),
    .INIT_2D(256'h000000008202066700000001e002068700000001d00206f1000000037032f032),
    .INIT_2E(256'h00000032b072088a0000001d6032066100000032adf225440000001d60220663),
    .INIT_2F(256'h00000001a002259100000001900206f100000032b442f0320000001d60401002),
    .INIT_30(256'h00000032acb206420000001ce400bc3300000036ac4206630000001cd302069b),
    .INIT_31(256'h00000013a000bc0b00000013900206b5000000108f02064c00000009f0820642),
    .INIT_32(256'h00000001d000bc0900000022ac02063b00000013e000bc0a00000011d012063b),
    .INIT_33(256'h00000032ad50bc070000001cd502063b0000000bf310bc080000000be302063b),
    .INIT_34(256'h00000011d010d00800000013a0009002000000129f020661000000108e02063b),
    .INIT_35(256'h00000003a03206d50000002f911010100000002f8102088a00000022ace324d9),
    .INIT_36(256'h00000004a002071600000014006206d500000014006010000000000b0132200a),
    .INIT_37(256'h0000000bd300bc09000000250000bb08000000370000ba070000002fa122200a),
    .INIT_38(256'h00000001a00000f0000000019000bf330000000b2370be0b0000000be310bd0a),
    .INIT_39(256'h000000108d00d00800000032aec324ea0000001cf201d00c00000001f000300f),
    .INIT_3A(256'h00000022ae50301f00000011f01000a000000013a002253f000000129e0324ea),
    .INIT_3B(256'h00000032af5206200000001cf50206200000000b23c2062000000001f002f014),
    .INIT_3C(256'h00000011f013e53f00000013a001d05d000000139000307f00000010820000b0),
    .INIT_3D(256'h00000032afd1d00c0000001cf300300f00000001f000b03300000022aee2f015),
    .INIT_3E(256'h00000011f01000e00000001380032504000000139000d00800000011802324fb),
    .INIT_3F(256'h00000003a030b1130000002f9112f0130000002f8100300300000022af61400e),
    .INIT_40(256'h00000004a00365130000001400620620000000140063653f0000000b0131c010),
    .INIT_41(256'h0000000bd300b113000000250002f01300000037000030030000002fa120b033),
    .INIT_42(256'h000000019002fc0c00000001800206200000000b2373653f0000000be311c010),
    .INIT_43(256'h00000032b1503f070000001cf202ff0f00000001f002fe0e00000001a002fd0d),
    .INIT_44(256'h00000011f0103e0300000013a0022523000000129e03253f000000108d01df01),
    .INIT_45(256'h0000001df0020b8b00000003ff02fe120000000bf392fd1100000022b0e2fc10),
    .INIT_46(256'h0000000b01318c0000000036b200b2060000001df300b10500000032b290b004),
    .INIT_47(256'h00000022b2120bb800000001f013e53f00000036b201ae200000001d0001ad10),
    .INIT_48(256'h00000032b290b0130000001df022f40f0000000b23c0340700000001f000b40f),
    .INIT_49(256'h00000011f013253100000013a001d001000000139003252c000000108201d000),
    .INIT_4A(256'h0000001cf503253b0000000b2381d00300000001f003253600000022b221d002),
    .INIT_4B(256'h00000013a0020900000000139002060500000010820207d000000032b32208eb),
    .INIT_4C(256'h0000001cf302060500000001f00207d700000022b2b208ee00000011f012253f),
    .INIT_4D(256'h00000013800207e100000013900208f1000000118012253f00000032b3a2090a),
    .INIT_4E(256'h0000002f911208f40000002f8102253f00000022b332091500000011f0120605),
    .INIT_4F(256'h000000140062085e00000014006209200000000b0132060500000003a03207ed),
    .INIT_50(256'h000000250002200a00000037000207160000002fa12206d500000004a0001000),
    .INIT_51(256'h000000018000900e0000000b237360970000000be310d0080000000bd3009011),
    .INIT_52(256'h0000001cf203610300000001f000d04000000001a0036107000000019000d080),
    .INIT_53(256'h00000013a00360fb000000129e00d010000000108d0360ff00000032b520d020),
    .INIT_54(256'h00000003ff0090160000000bf393255a00000022b4b0d00400000011f010900e),
    .INIT_55(256'h00000036b5d1d00e0000001df300300f00000032b662b04e0000001df002f033),
    .INIT_56(256'h00000001f010d02000000036b5d0900d0000001d000225440000000b0133256e),
    .INIT_57(256'h0000001df023256e0000000b23c1d04900000001f000900600000022b5e36544),
    .INIT_58(256'h00000013a002066100000013900206a5000000108203654400000032b661d053),
    .INIT_59(256'h0000000b2381130100000001f002071f00000022b5f0130000000011f010b202),
    .INIT_5A(256'h000000108202066700000032b70206870000001cf00365660000000b0371c320),
    .INIT_5B(256'h00000022b682066100000011f012069100000013a00225440000001390020663),
    .INIT_5C(256'h00000032b791d0020000001cf500b0020000000b2032004700000001f002003e),
    .INIT_5D(256'h00000011f011d00300000013a000b0020000001390020050000000108203257a),
    .INIT_5E(256'h00000032b81225890000001cf302085e00000001f002005900000022b723257a),
    .INIT_5F(256'h00000011f011d002000000138000b0020000001390020047000000118012003e),
    .INIT_60(256'h00000003a031d0030000002f9110b0020000002f8102005000000022b7a32586),
    .INIT_61(256'h00000004a0001060000000140062085e00000014006200590000000b01332586),
    .INIT_62(256'h0000000b0132d003000000250002f03200000037000010000000002fa12206c9),
    .INIT_63(256'h000000030f0207160000000b039206d500000032b94010000000001d00020703),
    .INIT_64(256'h00000032b9601f000000001d03101e0000000032b9601d000000001d0302200a),
    .INIT_65(256'h0000000950801d0000000020bb12ff1200000022b972fe1100000020baa2fd10),
    .INIT_66(256'h0000002f5042fd1e0000000960801d01000000095082fd130000002f5032fd01),
    .INIT_67(256'h0000002f530325bc000000096081d0ff000000095080b00f0000002f60520bb8),
    .INIT_68(256'h0000002f5370b001000000096082f00f00000009508030070000002f6310b00f),
    .INIT_69(256'h0000002f53c325b0000000096081d00100000009508325ac0000002f6381d000),
    .INIT_6A(256'h00000001607325b8000000015ef1d00300000025000325b40000002f6061d002),
    .INIT_6B(256'h0000002d10b221720000002d60a2093f0000002d509207d000000001100208eb),
    .INIT_6C(256'h00000001100221720000000160b2093f000000015c3207d700000025000208ee),
    .INIT_6D(256'h00000025000221720000002d10b2093f0000002d60a207e10000002d509208f1),
    .INIT_6E(256'h0000000b911221720000000b8102093f00000020b8b207ed00000037001208f4),
    .INIT_6F(256'h0000002fa36090160000002f935325c50000002f8340d0040000000ba120900e),
    .INIT_70(256'h0000000b4311d00e0000000b3300300f0000000bd372b04e000000012002f033),
    .INIT_71(256'h0000003abcf0b1050000001ba000b0040000001a94020b8b00000018830325e7),
    .INIT_72(256'h0000002fa360bf120000002f9350be110000002f8340bd10000000112010b206),
    .INIT_73(256'h0000000b8341ef2000000022bc41ee1000000032bfb1cd000000001c2d003f03),
    .INIT_74(256'h0000000120013f000000002f20f13e000000000ba3611d010000000b935325d8),
    .INIT_75(256'h00000032c972259a0000001d4012ff12000000094082fe11000000013002fd10),
    .INIT_76(256'h0000003abe21c0100000001ba00191010000001b9000b102000000188400b001),
    .INIT_77(256'h0000002f9352f0130000002f8342f001000000133001100100000011201325e7),
    .INIT_78(256'h0000000b9352fd100000000b83401f0000000022bd501e000000002fa3601d00),
    .INIT_79(256'h0000002f80c207a20000002f20d2259a0000002f30e2ff120000000ba362fe11),
    .INIT_7A(256'h0000000b70f2d0030000000b60e010000000000b50d207b20000000b40c20037),
    .INIT_7B(256'h000000147002200a000000146082071600000014608206d50000000b30e01000),
    .INIT_7C(256'h0000000b013250000000002f70e365f0000000147000d080000000143080900d),
    .INIT_7D(256'h000000140062500000000014006365f4000000140060d040000000140060900d),
    .INIT_7E(256'h0000000b4392de0700000025000205f4000000370002df070000002f00f205f4),
    .INIT_7F(256'h0000000b43c2dc0700000032c3b205f40000001d4002dd07000000034f0205f4),
    .INITP_00(256'hbf8abf9cbf8e341997098ca79eb78aa48bbfaa06aa12141e84b08d081cac12be),
    .INITP_01(256'h9a01183807351b241024a78da582931113a31d060f249d331ba79a368f3d219c),
    .INITP_02(256'h80a5be053808148d1e84b2b91ca585221d3801bf1b24351b22103801b91b241d),
    .INITP_03(256'ha221bb04bb032d8ca181bb0405a33a98081e331a849f849812179e0611263222),
    .INITP_04(256'hb81ba2119a8fa934b92eaab50630140f933db4312aaab7143b158c999200bda6),
    .INITP_05(256'ha5b322851b1bbb842e1a963d2b20a8ba03813f8f863927b6862d14352abf143e),
    .INITP_06(256'h8aa32aa13a18973c11ba9088222490853ca3b71789110b22ad3d930c2a210a1b),
    .INITP_07(256'h1ab91f859f14b52930abb21b87a3af1db58f1dbb9394a48804a2b725a12e181c),
    .INITP_08(256'had2c3285272196040382293f05ac8e8b0a3ea0a3aa1d9d0792ba2636a0990524),
    .INITP_09(256'h85842918a51aa28117a0b280beb629102db2879e019e332102a0ba970d8f0fbf),
    .INITP_0A(256'h850ba709a08684af020cbb1904b70d11a58015b33e3bae3d021e0d09a430ba39),
    .INITP_0B(256'h1293bda0382db2049137b408a9021cb31202ad3085b42a2799368b8d32b49b36),
    .INITP_0C(256'hb997052a33931da09732093bba16b4881c3e3c12b8b333b2b88594a50fb08d9c),
    .INITP_0D(256'ha9300e21a01227bfa6389a0880b5b6adb3801c8e23bebba6b91781b82d811729),
    .INITP_0E(256'hba8f242f3d1397110cb6b82d8903b5be8d27940b212c952b3b1e05bb9a251591),
    .INITP_0F(256'h1aa63dbf12b5b83794831d80ab98bf1d260f832a052ca9951f9e3b2caa113c25),
