`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5264)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5IQJj49NipZ8M+awYasSToxFXS4UuUEeV5rGiYBnae8zaBiLxijauuTi
wh/qiJw+J7W5DaDng1HCv3jl1xLrVztCZOUlIPg2a158b7bkH/gBtESeBxTmHYrEF2lbXqnY2dmD
fGaATCnjbLubIqc6LVxs4vWqp4I8V/KWIaSEaoMHdaAyWRqaBFOy5yZHp2viskKoc0FBRefPwKZE
TkKB9TkoIxRLLdbpICpPFmrNKRnLgsHOatqA4OmW+ljqgbFTATh6Q98Qvf33mAXAqohKF/toIxTL
/CrYo31tl4P60sn8Viy/911Kq5gzOuSmFePWA4h7azeoTIzJRznglSbx/sAbWqdtVFvY9s5zjjJQ
HJCHaptFJvKWLugyP5euxk54pjGzG9krpRdBc8mhJtSJhK/x8w2hcc5M1VdNWEPP3aF1L+hrJHOE
ALChnJP0A7Vz5ShlYEwFASIk26Z7yjG+TsBhyc9zCFZJc6AUmxU6LqFmzQMHSzev95NcF0EFoA4p
prFRaKpk98lVRjG59HYAzDCgrhc+UYYr2pD5mruTaeBYo+wUM2OyhdUDh4BWNoAVHBKx2pknIKp2
Ev7wYFZv3a9H8fQ2JqBPGfuXetKA6qrT/Jzwvh/t2akGlKRMQ18vMO5JHRlD0+Fx2fgbZg5VxHsc
NypBNTsHXu2gDBbhQhQDSGjqIwAH6F70wrZ83xTQTvx00/FAH2+CMo/hU8og9lfxZ2X1d7BpqeWs
N2OIXdw5XRw8CHNy3u1YiIQie6RUqlAXcjihLHIUoDPS+sPHxdpgGqhs/27RxLkZIbXJkx4o7rVJ
UhyWm/23MJrnj/6RwRIik3UzMhb3r5Z+9cR+fDIGUeqIzcnWKS8EwyUC0HmTt8HIVlyxHryyedv8
Af27CIEp8uCsJm8t/osD5h/VJW0PjanFxzEI7zaQ1JcI+0CILan3c2QZCyGBkSdEqFBaZS2hQEOp
2Y6BLjncT8CFhQ5/4oqAunryZrSciNbQT2XjkOGmf3PJe0xkAuWCmAAuFwTifilvOdNGxDtBTaN0
SEPwsMqtimnzmV/hlWagGwR2fTOTP2AbF8+WypgTkEAX80EEoZhVtqo9RGESnvBXvqIdp6gTDJQT
yawqB/yUMWEvRJ+EaKzeeuU5wsJW0uF/eRhgykyiHQuXs56ZPXDEFwiUqtnPENpAVjWvu8NA9o/r
7jLSHZaPaEF1b6fZFgIgGrEYfRSdgtr5VQ7wERWUPcG38he2q3a7avQ0SE2DWjOFIAM1EbbTaP/H
DVXm4xhxT/5WFruKQM7ZhnAKEsmDYJ9ws/vS5tzcl8SojWK2q0ttl/98Y2hlhHdiqYDve8b1d2K3
HEXvyLo2lWxO+cgv4uhc+l0UetFTscZU11xbDQ+Ms33VZEDoYpaY2HHwwMRz+b2Vxer6IDf2Eas0
H2IRIZZMV24XITBzjoTJmg7ISkr+2QWz1RrRfPQQnyeiDuUyLYe6UjPotYk2jZOypsUIz0bwNgaQ
4vfzDpYd9fFB3YQ+4/5cgxuSaOwayQw4rz/DqQb1EgbfvcZkmRcazBSX63piABvA/Vnx1X1q4TBP
rqsC1RBwFUpsdorNuIDB6QZ+EUjApID6+uG0QZ1JTFEtD8qUDtoHSpLUEUdSIWwai79qX4Y8WPIu
PSs9nIWpWFkvois+XXXkcimNrLs0ByP2jzDO0HJ43pRzfHOPdtsVZxmhs4phz0JI2yNqa0+W3Hso
jMP4CqoGOuSC+HchdoZG4Di7R0peoLaqU3Z/yBom/jNrFFWsI25M88BiOc5O7Nn4+ioNzARudQRR
mora1OLWXwgvKnkYIG1XuqIOJRjCGA4bRuin7gpzzqhSngCC/wvA7Lz1215UGB2tRNvwvr6D4HlH
UrNJEzYfXhc+8UirhvFwBft3plwsu31yuDOxEG315B5ymumQCII45bTg3kFk7z1wRHOAtuUz8SH+
fI/uRlAty0AmAe381c85HATe95OPa6+akGFQULw7NNuV/upqlsypNBByQ7gdAkJlR0CyDztxTflO
sjDCHLDrl1ql3uNVzHBN4+DYgk2JI0Ul9Gr1UMo1Wemw1ZirOcMqPjBbyQoHvpN/PZ7La8zPR+Ff
6WyMQpzINfX9kA3GvdQTpS1YRGy5uz+5h6GaD1VbyF+0kI2hVhTtwRKvSpgyNI5MBxcNM9wU2QLN
PS3po01mOl7/zUFxew/DIDbtLzOuUeKLNJ1iHW0gKUin6DYylQCkn2uHcdN3uf87HUnzvHQI06tX
kTaZpckklz/7mAL3HDEXJy1YeiySUWuA/hs9UuVGXVoizSWXbun+YGGA6WGa5gLhiDVo9LoWe5sa
eQIEUe1sgdURBQBi1qzPdes013LGp++ZyrN+bqLwr+J/1SQegaurFNQvR32fUFJkZKYEECshR1pI
iWYL+IOaYTnWh3DWZ6xnTctmHAK+EFr0kTcXS0lk/6f6lhOsw+uP8dIfr5MDuMLULvc6egCdFvB9
qIdSUMs5bPD4OrGc29M455epRxlf7h7LXxfakCF7lwgRAhuNievXYKUx5kQiQQ2EIVVvLMsX/FLP
BF2KqX/m8p3MdeMgHyarYcizx+aerUh7gIR3Epkr5W6pg2BmlRlb27wv58iWhqUDMvbIb56TQ3C5
r37FgGqwuwcBP4+ocJ6Qx5A/Li/yHr9DYbgwm+cfSFCbcdb9clWZpTQyLNFTSRBuduI7sZplLklt
lKZvW+vfb4+tiVSuZ3HN6jlOIUy3MaqcNyvQp+iuPD9DM5JnTbaR/mae+69eFMe+ovta7nOM+vp3
XhV6cJ2lPF+YCGSL78d1w/ZoezdRl5buOIvO49EkmxLUl1umFHhEboYUthGuNNLj4Mg65wSt53kJ
DjEFTdXcjNqGD9JseOORonw3T72dONpPuJjCm/rwP1wN6iX26dyRtj/HJWRS2hibn9XdbZLHLdaU
BmMA8JmEeKN2BVDOQZFugkfSXE+VpDgFPpN2a6rj++L037OtUaQfMo/HP7m86qrjGzfyadUxb482
MnyJTw4/0GMn8XDTldJ276k6V+2O7m/3iayVaNU1NAJNfKMCCHnGUryp3Y1q5BNBaFzuNoOOYbkb
43Bq5wpgut/DZByeNYjTl58oUxHCiThBAMMuUlPpcC8SIUKLAbYTyDAj+WMwMbSpIx/THcDuSt6i
qBMXosorkVufSbMhzncwKQArelb2CbI1qQ7kIgzxxX6AD+rBe4ljY1OAXJK+O7TtDGqnq8BmSYyq
iRwjmhX8oLjwFDHATmjtYvF/gG/cYCKdLwyvdaf+TecWyJ6KkRv2WGflE4K45opCxYMiWPSDQj/6
xUrk4uG/TY5/7TP/mveznl7psEouVQpL2OTT+N1JcWvmc0TPqTbuIY/FQLuvMr1qAgF4ni6O1RXt
S57hgrRw6jV/bFC5t6QaqeSIGCb2JAYbNGP27bh+DFo0E+X8zzM74H1qTdmQuD4keOLS8IZeiKa/
6G57e7xOFsRueGCpoqpm1BESK03OtiI+OB27dCFzJVRZjstMEJUyWspPtJWAR6sP9eAeSzBr/izS
cpIS2zSAbWQQ/AoLtRizx45bkDxPE3a5nfQzc6IgO8iDzINxUJOh3FRq0331Fzj6FzKmswEgom8L
mgjVl5Ar4bAcgv40Y2nZ7R1m8S0uZYNlRsbWZ6Qi2kAy7Nsf/4LOJvYBsfF1INFcxnfN8W5D059X
u6eQUG5Nw88tvrGSEy4wByA/kgO1ky7iUp/+pV2hJwuAnPQjQrGg6WmXMHgPOh4Y9578kzOwrTfD
asG66sf8KXWXd5Wy/fGbcXDM2R1Brf7HB8KNnJ/i+VhiJsZgt8sQsaB+CQ6oZX92pCNADfiMqviG
uf3QxY8rO6Y+Jj8u8Lrj2TOW8UjTUZgunl5RSFyZ5uPLnzF2PvD425m9bGu0U3Y3hKlPb+qgCydn
3B7oSmgeDybWMqsDVd2o9PNdSXrR15pp9WQMJ+R5uPvUoUX+Rwt0l/56+e/rbr8DAKryz4+71JMl
5Z9iKD1TQGTvo8umj1n0k+Ghn7yE+W+v5TA1xYQirTqUAS7GoAz4spv2mdMIOgc/g+chlsspcli6
3ivPFQEDbpR/w/JQ7xA/i+16njwzzr+xblcUX5Q5CIFZz9EXQh8VF9LLNHyCpZ6AQz5Nd0tuQLow
2i16lfsW8v6Vy8x1A3CDC65zRRhonPv0/FClz3PM6Je8VCCZEGXng8MzyfK9eNPEDzxl+C14ECXG
wGHXe4HbUNvy7/cKoiGf+VH4jmRB02kUKSqPUjIykoNpy3EQO0SDsH9bTVTxmrYjVzP7YHY2/KAJ
/L11k5+/9A/p5J4GJsHWOUQW9ci7mdwmzBxvlskMUx1LMgs5uAo6LNK/cqRCuwtbrnt9JVzmAvyX
34D84jIJtIi7AVT4hFCiNkdN4JANtz8K4byWY0zJ3jFE5Um9JpH5lmFGLIJ1vRyR+U/ZLtGUOh4U
iL3OpQj/XGD8dYyWSHiw2JpaOt7XgrVLTWZlfsTQnvgM413O5diASNL0emH2nvXdUIjJ4dxCqwQH
fD7lNmviiieg4KPlVWcrUTuHPiKPT+sNUl8UHaYobgel4hco7Y8WGZfRpx02ps57TPk9ylY5mHeP
IqKrAUdSC3aesew5ST1wUlgFDsZM83Tik0XJVIOZZ5gG3Vu024hovgbcT5dTdWPGzLW73B1SLI5b
es3mckSZ3l12LT63fx07ISzYlHPhMEE2a69VUmU9uQRTCSIEd9OC8Al0kzaCCtOh+BvA0bhwLgR+
LAD83/uyIlTm+AjmkeIBMnZDDjfL+9E99/kcVNlk9CWoIZ0So3Oiu+w3afw9DoVB5ZjdkW0LXhQ9
YjE12iFKX6gl+PYpZVDLl90k8LiZYrSgUT7T8MxCtTjmBcKVbmSc5qrQ1cf0B5G8WLHnmzR2myWN
YRg73tAJKZtqqmm3GLnpQXBg3d/AGVtXyCTflmx/D+/o9yscmQ2SSI+CBHzVmcyMKGhE4mkVvzhD
lXapLKUeDm6PD/f6d5HTd4rySSukiodWfCxobJeLwMFc98jmgYdlf6fdSBtBvsiBcoYd/Qop0dk0
RK7ycKxpgbqyU/gl9Hdr7e6iVlJY7IODYcB7A/IP1w7iUgbPDCCbwXhSBIQHKY/sMdba+Pt5kZ4D
hnbwGK54SRQv1cSZ975AAZliFeka+alw+48M3nGqPdOlCPWvhPAePt1KEgLEaUVClgaTlFOjMuVk
LXvw2FpZKW0jcIrrTwrJg9NgLS6KgZEN1E5zYyJ4VDbsi7ruBMLAb0JgRiG/3Mdfm+tGu0Vz/KGZ
WniQg74coz1xgvUr6KP1jOcOywHXsysT/Y3lJM7GN0To6pp5dECS55iCTGQR9tRuJHJLdasRNCWo
AxTB5wQBCsgBfjCIQtxdaj1RjxUk1/MIByeYZRq1SRF69pziZ7D8xsLis210jTm1W6v3Ch7G/ohY
l5/zCKOIsXDFiUjyxsC90zaU6QZ3GV3hOl77UKaP1vm9Fayn4SnGSbYNy14j12RhcqSnNN8Rs0jA
aaTc4eM9IwJkeyw2Bfu2OHsaUDd+MbJDoutR0jDI3hyepzLRp5cDH5oMLEq14VqPe5a6y6osvb3v
/w5NMYucKd0eBbC0cAmtVGN9jFKzbvFqIXBl8PtblLGMxrrGg9S1u+UhIOBhtAKUkY6dduWYGD9a
Tsz2gg9tNxn94I1XVMFBdEdtRirBh9u9dSbysw7Y0V0++rheuNIqxX3p/JrkXetyZ/ewpVUe/VTR
+zjBS2ihgy7bT735hXWA0osc3H8ZTxUPlTLfC1aQQ3QDslF+7u6rtL6chiW+AfmsUX4exNTnXyOZ
4ip7fkwElOx78C08lLX0MXkkYUQNxTxNGAMgP1lo6pPKX38YGEESt24XGvx0ekP5rJfQH/hSenjp
EstJPCWpAW/yks2lXHM4J6yIgMtI+xI9CwG70D7bft1majnHNATSGobPBYWslack7+/cQrsON4OW
4HmXzlhlemuhuMyz/ioiPaEoT5BatOgYvxD4UFEXWufVK0hGtTlNn5Z/6vxbvMlKd1Zv1pK1yWAv
DFE323zWdsEYN2bLLrvQ2O+S2eRwii7XVZGX2htd/5I/yov7SKPgQaYEZbHtFIiQ8e4b59kMoG5u
3rPQozYYTKGAEuMe4tio3XSNarlJlPrpHQ3PWNG5Wv+UG1iT5e6xSmWjwbxiFtQsL+Zm2CIhWUjn
eg/ddHBY1f7aKLCVv9mdDeHLFRQDd0xSlFP7fzOFkC3O7MQoPQSgEJdxD8re0XYkh3Uwk7rPjvqq
ww3d+/mHUiypK2VwSvxEVJB2EMAEDLSCcKEDs3mYL/MavA6NxSpIFFxmwIfrS3nRwqqxZSEJypml
CYzpv6c/P9mTpgdFvCwboGP4O5QJX+xYqSG7cOs40oL7Te4Yugp4qnPk/EppGMZyI4OJhhlyahAN
Fwjh/0od0/AYjTTKbtQ4vOdNg+lEX8FwNuA33zfTQLTVTKLgnJ8ny8syD9Wyae/Izzp8UaaT0BgQ
WHSznA/6MaewEuB/c3sjbmI4y5Li9sbPvBPuG5jVJIvAlyzQFlQyj35WCePpa7F1TmmqZD2xlYzs
o0ZD6R7mWoDXE0Gbe4s8CzbWXugQLfti9VLHWJyIN+zGHAODn8XtBnOQVGmMulboM/pJbW/LNGXV
PFgNtTfO1eUkYIHNjIc5vKiE5pmaJyEhLVaQa5FPiuJCzlhyhBFDUuuv2/E7ip/rKtd12z5ea4Dv
k1SUIaQxgi0YOzY6PswPm/gUVadE1g9XCx00SKv1XDaHZeFL73qqozVAg8zrBG/fwsa/Nbwi3ywD
Hh58vmU+O6gXRHA/cHwhiI7oL9uRUyNu5sPPhkKbzLOAlqH1gkpQ4LUqAzfpTV9k4Q5ybwFINbRy
wjm9L8cxbdJubyM0ifxue1jmfVFnrbMypFvczVVQ9JaputPdNYsgkuZStht0rxuRBmgrSE6OTepp
TcypPV2xRp40/u0Nze9mfME8VVA=
`pragma protect end_protected
