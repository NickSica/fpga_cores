`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
iQbEix3JHZTwa1vhipHlmwS1/G9xw/soq5c1aH9r1Ikmd5PFC6vG8hcczrO5Gm238/UZKbDRHhQl
8vxxX1eWXA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NYO2r/VW0Uk9iILO9avt3Skw+TFdXKrXeDrkjkY6MrmMZXqmt1ljuTdXla3Px6GiDC5iNRfSB1LJ
jlz9x6ZyMo5VxrDlXmNLima4xlcLjwQ5Ldngl558uz/vr1FbORoJ+gk4f03PWwyf42EKOYFnCVfd
LJfFRdBml66XWTkIRRs=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hXM/negBdYIePK99VNL4dA9qZWSDCbIcZGIF+wzwJF2GeTdZiC6Sv8N9/cF1YoJ4PmeE+1cpGoYE
hr+rxDAb1wjgZvfDyEG1QWzKRSG5E+oNC6Bj2Xk8erPPxuHL0sXJnNFmZt3mRdMMjzJ/oBGkUF0h
iYE6DHIS9BMznThGr4tm6wOQ24nLfv2CkGw5FtsfpBEceglyVNwc5KmDZpqUutO1UmcXWgUVf6aG
3t7duiHDJKzCaRYGI47UkrEGgYTLtr4N4clyKbc4ZaAFsMfafXuq7UodHyHPGa7sQYA60+7yMSq7
lZ6oowJsQLQdpXSegbc7gK8ezWVXMGToMCUX4g==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
IZkumnZp/JsuGCxK7A5f04eL3wOhVC/HIkiq9ThWDUN6/jAV9gkhdECfPCdAYxhe0IfGI1mwNrRJ
CATeVriO+TbtGJF8trisSNtrtJxyu7w+ARrQ3i7xJ5OugSeDn5jrGtPVCeIVbs8Otz0RthJD/ia+
zMRiRhN8wPr8+wtwChbS7LbmoKzd361OLqaC8TX6Ab1GBUHFOMfYyAPJdl/jXbS9u43VHuRY6Yc6
WqrfDJE3842973TEArl3DaaLzZwM28WBp6JNk4Z1zR+7/fPjneoZl3Dvksdx4ThM0a5s9BNPAH9V
WF7gF4b9Me6TfP8DfbNOy0URIYx+xbfpe++9uQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eaRvVH2iXg+bRFhfU/Zdu0OhZxAtLuP0NVIWmdEUooi3G/jC4AtcmpPrp7p/DrHH2FZwIvu+AbK3
sY3ybtP3ICKGUwlnIt7XryFabcZX+wxEJ33rwyvMH3qSJUvv0NnXC8IHlKKyRjDylY/oANDzbz6D
+mWDv16FdHx/0RgRk2HTfCPx8qBZ+fT4hbE6exCfOH2KzbFjubsbEmNkNU+HUDcusYXP2EoAnNGO
lFufKr3GhljOMYxxaVeKpXEcKWjQB5Uu1M3JdONHHSUP3iVPekneDcajTRMfHD9FJggiLA6mAgel
cdhHqUxScYsWsL7cenQphjXngVDIxqnSMZgGGg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
heQDXwsWtguDyBBqy+N/Xr88McxL4tQSR2XBCb/lxs8IKaambMExKMCiF+uYl01VHmTIU2W66UkM
7t9z8H1Gdw289KkEy+LLNQNFvy4xiQp3che0cCrsbm5/JjwMeuGavzmF6wwMkz5sW4oMgRBAsxzn
RRGXDS1r2TiNXhNi68I=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WZqwWujfHGXV7wBEePMjGLVWUeV/ygCmf158CXpAhJC77z2vuuagSDsOpGgtqyakG2cswti5bhBy
iGqPgNkEY7Q4T3NMe5WssA5nf18Sw3LU1MCehsK5WrHeKiMOyz9QpdgScXEE86/e3qniqvFlM2/c
HpI+I2e/HN1QOgChXb7HzAEEqCCdY9VD1a+p15IoOmU/8Gs718QdaPMJOt3XdTu5pAmq/PWuICaZ
VFSPDj57xVELte/pDBIXo8hgI5sad9ci34UyXovDzhRyUKzLY0u+gqRalObdZFD1Ph6hGQiLfmwO
JTvUCIjoFwTzhh0dCXYGcwc8O9kaaOIiiwpgyg==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
B4GVIi6TGeAAKF2mV42cg9jGmUkeJ9TkEGN3HtEus1MF1Zmt7Nh1Y005XEEzr57ufgLlM872beae
bxX2U/dQHyW4OCP8KBTn49Kmkdu8j6t5b8W5HRsXXHYSGPOo9IxUSHBdhwxHpNWauRDmTFNl2lia
Ton0toY2wVDxIcyINRYIpxD8YGHOnHSHPMsgAGtuP7kRvUnSvNzqqhzVcNm3oeIMTawuhFgBXD+f
0S45sDt4HAERXJfO2RXmlDCCLpg7FQxibRHwoppbdhT48SpFRar2SU9FLaP1Rhu4f8UN/BXG8JDH
IE70hcE1uVmlqXL3h64Aaql7Kf0Mt19/bANOBQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 44400)
`pragma protect data_block
8fgGNC4HfskTXIPOSZDcR4TgLnemdzeM6AviUAaUSSdE0upH2s5nrjqEJUNPx8Yka2y2wNknc8bK
wDdnWgjKEc+4qC7pdVXffrpP1tMF1tjkvoWB8xKZwLoP5bfj5JRs3mvLz65wVHZUSzhQFV9n84Qj
eUvg5RjUZoeMSBccYPgVjoyv/WFDe8xI526+YhnOOClVtq9IZJl7Hwo4gWfZeR+EvEaZUJsZp4Uv
wIJcjtVy7qrKydnQ2bCzhaihaVkIAsN4j+5R9BpbFUVjQUS2ve4rYobxf0R2zJPGsKI93+CpoKmY
TgeYnPrJw544S/DL7BAbHU0+k73kWnyhU7IFfVQiv7ZZRNBz8lZ6CrV+PESMpNfO16Ivry+hmywv
WXcnigz6DdvkdQPNmqsXKuLedNfnG3hht9U2Mlb/0WdHa6+iC07MnfnxlSuSIiNu/WKlh0o8Adx0
mSri5aqaTTbRQV9YacCaiQKOWTs/wIMMSzyM4IYpositw982I5oBvozBSVX1yDe5pKFzxmSMH/RN
erx1ium+K+Im60OUsBQfDN8pvQ0nWnF3UNQPVL82ccW+kU8o3OL4YgWym+JYeif4u3v8ds4+FBkU
fQnTGbR7OhgEpVUNEN21GMkMWPxhpS/MKGMrYpmP52Lq8agCZeWcL3cJIIp17ZXOkXOEjQqaSVsS
iQcygbcrR0VQGIQ70yEZXGJ1mfDTzm4jrW4DoOi2JmXN23LYCElX+X9Jc413Awcz6mSx84QcUg4J
n72aoj5p80qkH2pHtZqY2yY+FoKPu2arzyvXj1ktxSirsaJlILEcc/h6tMfjB5ALx1/BmBalC1Zx
DNrnu82Xm7z1GwwNi30WFD8rbF4A636zVjdWyCWd+SmSFkQMMoKf5/C7zZtVotSr88u/1xsJGXKu
pe4W8oIqFy5V1+Ns2g2/6FaDdoY1RWyM1l9xj3ra6u9ZXm2gS9oYmnd0OHW+mmFsG9JqBzRukf18
VNefZmIkS00Ilc2irGDyrI4zxpPHB3POl3w4I/r4BuBBU1Lvsh7tKPV4o3uKnNXIzD/Zs68SuJwW
2tR++n66PiKGce61dKoVDxqPNt/RoMSBw4KPeTv5jY9sWv1NQMaAnmTBFIUwu60jFB3UZepxzCVx
fRs0uEnmXtxdHH5tnddOLBasJHrbIOzVHjnJzsEuAmKATCRXXGBt0FNeo6YIGw2a0ewDVoQUMF3D
cJdxSgazjVN3Bl1IGKcJwlK1JkTcyUSfY32Om44KkvnE5MPlpUxbCqbZ2xukF/+9a75pcOKj5BzF
n1GJfXEyKB7ZMhOASHD4BIcsqpkI6Re28x9iIUBqV8MR1AJz5SXrENpHIgbk47T+cSZ5lfH8f8sA
hjrapgk4ayuGTfL4dgMm9isrEd3kBK3eRK7cVXkg578MfS8rr4btVZAwAde94v7B8QsKmS0K2gcV
EgtFgbHe8cN2NN+fKf7fEDXUGwPijk3qcdrd0nLAJdH+eoq3i1xhnxjLN0hWcbizHKk8j1Je7UWR
bPLGlqczA2UqSBLnFm9qTSK2VcPBYC/XZhNGlVy/iN0WwbCn8uOXFF0L8HeizlJyjqq+qheTHqby
jXDoEjAD4lAiEvx0rd1rhEHXU0EdtT9QVsFjUzNqfPia2pGQau6+d92zwJf53XzKeD3+b8Oj8Wx7
Cq3+rzza970VJ/RYdMUxdimu4fDD1DoHbYrb18OLmVIP7beLWkpaeF5BqZi/LXebj7Cd4TJCjyFI
cwm172qN/XNTsEBICmfNBIqw3VbgZobnoaIa0x7BTudPuXf0FNnVBB0ie+Mu2XpRlp12d0wgsutO
nxe9kHbGeEHoslcj2XM3k+Epx5/l2RCrLflq/+DthKJk1/SVy8OgyPKq1XLmdKPFskbUPpytOnNX
LImxhhI3bkwLkDLEwktvNsVZLbTHgFyv+7IX74iTGpNSp+NZpblcAUqvZ+SOq/duTus0Nn2UiGiN
4HWXrueDFaEtPR+WNiYQBawV1RsHIxqqqSRUL1qrWjV7T3OIkGFC0fZlOP2S5JhCYInoso+wWbJt
GuaWh5NPRJ/KP51sFzPTp3m2O9zR7sCYoP7+zL1b1Eb80RMOtlquWt+skwWF2yI8fWV/yQX2P4RX
s3UQadhK9inVezZ2aSSgIK2o+JS3p9gObrx/7gveo//2BJCursIlOvwnerlb2kAxt8/NVKsflOOh
n62lKr7gQttSex+M7T6SoOkd3IB/7xmI9+OLsdTtzwQ1Vh/aNC1fhSC8gD/FT82qt2LlXRi/0P6c
YNR1y4mRSTJ3a6hl+6MgWjqf774GvrRNC8WrIt6K+uAcr2jv+SURRjU1BVT99c3gc8sTZMwzUjko
Q9cAMQZByRlkzKUX3IP8hUECqmZlk37A8Mh4YKxCMClEa45qk0oAM30p9Sc13kp4/2EIuttk1Xn6
LBJmSowJJBgEomvtKYZfNQxsxnRlzEYB9l1mLKfzJaUGrz4f/msCRgy71vY8gHRI++jUAoWuUX7K
yGnoYtDF9kYycsTNOAhcZbjNrnrjQ+R88RPTU5WEY+lFEekooCZyHsgQWN5+hWyXelh7amfNp6ip
SBDsCJPiE2N8XLkJtkvui+WdKp+HS4M5/r4Tk7gaYVj1Kq/1OutyI3XYYgLN6eai9gKxkXI1sCRa
P7aMYce6boooD1ZZicTjRbuXBrQhz2qhB/gZa4scO+PWqZBqrVreP6x+j1qa2+s0JM5yzH7jNasS
7nE8W4jh0+mg7qUp+B2el8A5fbyyA1nc9ZUjZ5vUQ4rZh1y2mLoJQGxhF5k/IXHunV0Oc4Ts1Dxs
betYSrzSazZFE+hz81Nn1JpXkYmUoaN+NDZmNMjwJudEVmaPJOqhKx4HoUMWLJen6fhl5/aSv/qn
gFEjtpIEHFJc8VHDijRjsGfFs8GioAkSDfPqxiKuwPwbfdh/iaHGQ8J3NOy9bbWzamFKmILg1pyI
IUBGG2MZL62R7bKcTB/tAEcCeEVhs/krN4/h+8I1rlGAqrzg/Sp4pLIZpVdPtvqNDGLfXqaAdZRd
ZELskgYaRP24vtOQryNDNRWAVAnhcW+kU5ny2VpmD39Tng6aseJim/uTONL/9vE4GumT1lc2RmUu
EXkNo4zazlqFKCSyyKHB2DsUyrzffqH3nmZ8yaRt+NMjfsHfECV1oJVvyqBWOkagJHfoY5hl2Gts
L6CDaTjygvmnx4bPpfYKxJIK4GNAA64WV/OxrV4N518tfn6a4PJzXfwosX9+GY76T9maLIRMWvaU
VBJ1uCnLnAYF3UGicKJOSw8jq6x4lCSiYbSOS0dB1q1x0fUpnGhzG6WxgqoNNptFm/HyWa3fGnpR
AYeaETbn6Lnu9DZdAurjZdrd5Kq5QSf1IGdX4u8di+Cy5JhtS5T+71qhIm3GwxhR+jGUdoBUYS8U
3ocEEdymt+YjqxYkXWW2guADbFwRob1dD9cihiLG4EKvnUILl2UuYDlQqlZ972XAWICPiJ87TE1I
21bTYAY63j0328AM9IHRkuehjXvWkpXb27a5Yp3YXd9cDV34vIfj9eo5nevVXqtJOCYFlQYtBmAB
cSm9T3ErVr++mYOk5KB1yPjKQazcazYUIx++95q5zsOYlKdfEtq9/9olKyUe1zRALNMEJGGx6lGQ
ckhNa6xLr1QoReLuufH+cQR6wpjyBzHBlwuWyVOF4cpZsJlAfZVHh4D8BeIjx6C+9iKxMrl/4brx
58LGszHzCGA6iq+bVt7AZI0bYHRffLmKBrzk8V6lcUxX7obu6F2nY6vGxnDozN6NizEkpNU3IsA2
kSPnDBa5BVAYkl5WSbZeouiLeDD9dGzgBPtac3XTpda0mPm229bCQq4pmcDm3/Ij2QfRKNeeQ7GE
LKgFkZrkXHEt4fuUSWYplre7GcnykRHczKxqWETMry/12JizDQfj40eFyaeAx7XX3m0MMJ1olVeo
ian46iPB73xui1yACiDX8E+o0uqKHLkzl6gST1ve4S3vvObvGG5O5fV0AQR6Jo5m/K3vv/v55BGz
09sJDLWaQFtSHmhOOwsgrZ8MC1XAFGKvg55oUs1Xof5VsUpdYecCA2luA2BAp+UcGATAhaf8d/NB
POAFw1hymkH07noXYEs/O5nOQ4G9Tea0yJoLeaehZbzhk0rg5Tt8qsqEe86Lc46/Z5qzxOw0nCdp
e/KJqdD+4yBddVsyI0DFHoEOoCG40EG2aM36wZXSbyLaCxp9TDpSmSOZlf4idA0Ym3ocCaKpdR87
7rOiCCWJee6DdZt36Y3bsScqnlDoau3kLybPq0XrAJDPzaKZTY03CPpukGpywhc/n8DM1DDP1rNH
SEBSdWiDIuviRxa5fNnMX5EMemmxrUJLpQApXN7iNSCylVALkhurH+haZGraf3cKwTsonPpYTMUC
skIFIRzhK8o+lkXCZm7n5VYJWEt1Wd92C+u/urug408mdqZhWESvRdmqOUbiRwoMTJJ4u1QQM1Wq
P2BgffF6aFsQD3YYG3Z+ShnFKtXlkQeIjJdSQF98Yn0pPE6WxY4Zdyj+ATAOVU241dkEnhCk5UC5
w0BwtTIRF30rMtLPlpBXYEYw+TvQznm0Os94HJA9omxY+Hzzmd2m/hap6X7+86u78IM/EaSk3Eg0
2LOTBYLtLijqdD1RqsQ5sqiZnWaiWgKxErKw8rI7FXZSlEB/sLZHQijvYhJVzn+t9iTWaEMKvMEW
kw6Sv3S0chXICCQ7991OBVsEPIXrREBNyaNS4+6vNlU43j14QXR7DRu+gx87B1RrMY4/QXJRRveL
EsrWhihqC+fN7V5PuA+OVsM7jC8Irtir4wAc9rtBkLymxaJXYbQXp3Hqkwm6d5GVPeQBZUpFWCZk
du0xzWhE5ZITFn6XP6rBcF9j1jHKJwe986CHyYzJzTg9C4Om8UpBY5EF7TUSitQZRUmN7a1ySBy9
Iw1ARsyWl1gaCtAT+oY2dSLvxC+JJwyEs/QGTwI++uAjIl14NPgxZ1tVZsuCkDoPpB44WvAKExmW
FMYZzGpIYGty+6H1fzpUwRCI+pd1Ezte0aZM9Y7EOi4jfM4yUH/Cy2njgFNCYy2oxJMhEp+6d9Xh
6ysXAatrPXSQypRLIn4V9rpISbHnt87+B48bSLTITrUm3s6wjodK07qkw2MxODlRtpNwT85F1KEK
OL5VDUkA0Tn8L0aoZbQBq0JwvOx9w0HhTzng6cPHVFxPm1y/cztElfgSyapyu5WZeuDNOUOU+4bm
SKOI9beOmcHgcMGgEHg6hWZGgQBRFP6fxsIm8CVfiC5AVni9vz0r2rYkIsiETjKCtj3PvcG0xDkG
4tpMsicfdh+G4jx8XDEXtS0qt+ua37HBRe3MsiVhPtCJMGbsNlEp0fUFEVkYNVMUNJhRY+j1wmn3
g3cGi0GBjmAFZEoSaSbSwZ+X+aIZG7bGivs6/sd3PkD9P936Tj0A/7W8PEpXqqMafmlXY9A/+w47
53kMbF3jXafUlRwhtWw4qUhrMSjAlsYPuo/SCy7HOT1h20ut4/bW3DOuz4WvPYr+1mOrbi1X9k0v
7Sab13zMy6WUDSpUJe5Nr2SLX7+J18YOBXrbtGCB4V3KAtJwv3bdEYfp0TuTst/fPMQw1s5rb213
8xBgk7/ArwpP/f0n1cStxkYXLSDZHhSlJpy4fOe2aU8XZRFLoH8Qpnl5IUn19a0PgK4GIhGFoV4J
j7LhI/9UW53eRozQ1IhbaBSaPq+6fwDUrxJWCmI6VAbXYoP132+/3IiMZ2Er+CwIkD4dJTjVtYxL
QOC0SdSa/ELwuHY1dqJlBZD5t+oBGvwynFychPWxZ/aCwcnJtu4fKm7FTdZKW0IZl0zQIjr9L4eS
k4SrkTw5pQ0QnwKnXjiQILymmiukMT6mCCX0JoXvVM31x6Con/FhaC1uPMUIATL82dZWNro/Mxh7
ZQDKd9/rLGinLBWcqKtJb69uOPeQq/khEz1oYrIZWtoA7yp8GhCCiomxtKrFx0qlBVVwgB+7vuvD
TdSH3fgj0fVDgZwkOsY7mbXJO3yq6H6oD95enrSAI/4Sm5cDtdGYp5oSv9SDHNFqUm0TWQIeAK3a
Ge9GOFy/cZ9e9wYo5Mt2GvqPBVIopxe7I9GiPeUu+LdcwQrZXCF8BFnze225q1DuEZNUmXPN0Haa
9T+FtxOpQ3aKZcwgOKoCKdIg0RuXRpNC2WIpIBzFehoteiMgY9ZcBrZXtWPdlYyBnReEp94m7hqG
6fVMEicVVza8sJ3Mf8D6hsBWGdqZy6Gh65AUb3zvTCU7jp5IuFMStOULIQ1YsCYcXM5mOIifvFCh
n9WeVNax2d6CbaNu7F073+2PumjY63V6pzBc2+X1GuRWrjbWTDb8tkkG+g8AQpiyK8l85VbTcCWR
tm8v8uUz0k5l2f0XbYESiEAtsVDsSI9dtY0BF1bb/BxA04eBapLtm9aI/MhDvKI7mNzuhffCGEio
mB2w8kUxXfw5oY2oBVUH1YH2TbLxx5xU73I6lkgkPTWEoirC8yV5p+fleW9SydRUqUv3m+TxETHO
Dh2oVCCn+gs3ksZG1KM7BfhymTUy9OnQiMgoJqsBq0pEHP6Cf5iLAUZn2watA14Fl7fh1UTAdt9j
IvJvBPnHSHEfUuNaOR5KPJmcwOQ+8E7o4/g9iBZV1x/7h+MWGkn0yp3eQlqerZqmUetlh83OBWmm
RMSAhcGeq6hYJSmrcOCVYDVP2I1pFlsM6ONXh60qhdh+ZsgyBqRp91QcPd3psNvb/fzapkQ+reAJ
qoTfFLuMKtOaXuJ336QSATDu39l1zYw6hR1rZq6/eR9nQr9m5hlxEwM73gwitd4z7I56p1oGKL/T
PJoI0owugvU1l4j3mWIJ83BSAki/fJO7GBwDe3W/rPY3MVQ6tM75enlAdUER1zSj0WTK//R271Xq
8i0YOmlZTBtxY1MgCwXq2s0klPXSiGPoOTdQlHS4MRedJiitawvhQvsyqZDNN44cX8gcfJ+D3FtN
5SjMa2uNjDfWyA6RdsogeKv9Gl0qJF0CHPQ7SK/Nr5NprCCYITPpssNRTHCU779Mh4hJnPb49MK8
vrd76uIL+oRFx7wlnS8/DdaHI9u/fDGXslnKYohn1L7mHlrIc/3Pn14W4d24l1UESjUW5xHWGrUu
gMXB5UYuFYqyb3VUputxwwJ8CoXtwfmMocfmmYYIPvDQEpursHlPfXZLF6IqBivJ1x+6jjJB5ZRS
n9PLU6AyUoRGptFNca2h+sKpQjsj7aj+5GIv2QoNMSaP3qXGpcX2QGiohPMWtdVEfr7n0hIqDrYZ
yW0mi3GBRW5VxzDJGs17TJU8DgcciyhlRg8CQfdWjzkeKeRpHlmB6SwTJ1q4Gv8ALkHi+nzlRXqh
IjTKo8CtFQ41sd7wBTLmV1rLTRpCd3KH6BGOEYVE183PoacCL6dxPg/FDOPto3DVVOrBs29iS8Wg
luEweQJM/Z6NIxMCciWo8QYoLLN269v9iDvy4NKthEB6Dt2F5/jtI1eGEQ3FdEaOvNQW09vm8dt8
4L0KCw5aj3hnNagPmhnB4xU4xAHiB/fquWHKrDKPb2iJFM/cYL2bvAS11jZZ6zRWyhqKTiHlzJOe
tktlgaob3LypfVMf5YCBGTfCCG0z9UxH43J89ZYOjhUgr9t4wPSgaYtAvK+1NhniQJtuV1mT/XNk
fMx3gJKO1JyWsuv4e7I9c9NSgLlPXuogIkQsUyDK2SNuacSE44tJxot6C7dLAgYTFI8wNqG8WQot
Shc5II+/UqXR7oUEe9FINOCctfTeMPXyEnlnnjTYFpXZcv1OldoSFQNINg5J28KXvSHCMbrP/FnS
jrrkTOW0pYfwW1Tn8rqpPm9OvyIAkLEsPGuRxLjbhXr7sOzaJbKAS0jCFfYXsDq5moI9G8Effy0v
i2H05dbL8HcpiSd3vNGqfd+cpukRPhV1ijxdgVxfkYHVdVZcY3DIVJfD3F3q3x69lViHgjZH4gcC
ET5u8Q1BB8WHjVzFsRuWcLB7CSSnw5mt6mJSgqjJqBqsQdLOVhF3iYLS9/1IemHBl9ZEc3nrgKT5
48TYo2bP7Wf2o0imF49dpAj5Hd0jxg2mmhoG57vnvnVCHAOI5j2O1gMOm3PFGsdXENqThf4SBaQK
D61b5p9w6DYH8ueO3CBwoZfSW7hMLHlBx6Qw18gkvfScDcBtdUKlD+KhZ5OVwLK5hdyG+GPt7KUI
iho2TbWQnELrt+MEWEe/VjHm4/mMavCLZEGDMoKQIyNeSgd+mhGjE5qS/uWxlaOPMQODoxEEpvPe
QyfEcoYaqfvejSiZLIE28Mw/Fh3M1cG7aii55wrP3MVtBxB4n+oEypdfSXBVWJM7f3hmsCOVqBE6
qgQsye8q2h10eMbb0nNmh5TobW0Ooegv7TFofbLuqdIT9/S66RWqSQK/m2pqCXHiLv3xz2uoIF4j
ecpcWFzyo28yDyvdACvup5Ik4zsaQS4tQ1WojIYk5qXneYjGhFN6qUCyYXUg8e6jwkL+3XdrZGnf
SF3J7DYi/YAvq1mfDWWn2ih01KfIU6UjDyQKgqVbdzh5GiSSh12QAL4apz9LsIWANte57A02qmv4
o7Otrqr5YtHCAP3zz/wA8k5L+QPluzTuDwMXQfQKCN0Ys5lFdrHmFrkvvJWWw0SuQ0dtDgm3H7xg
cx9qphcBIZ6inswLeXMiuS2bBPAYj6cmBHaTBfFHarMfRMviBfhESfe62C2x0inXhJ/aMyDSk4It
pyPca2UXGkKysnDlXGR9Sny/VrmDcvcVGByLn+T7wYg0geqO6V9MAxqR0F6V9lCfg14P8NND8MdO
aSFHFvK33wuCogzQESCPpGmoPqh3rOLs5h5KTrUAM4mfdBz/9htK+b53LHfDrWjQBtlW1uyRK9B2
brZX0CuycwW7wqkuhsR5qQWSG2Shj27QEzf1JXXRbslN2r3v1HczfU7wKukIheLF98StWx4gncIO
MNMHM1A6PCvkv9zfac54rk8gM097b3N/cVZeRijNt4oN3QfbYJRacObkln0QC1jmIZoVOOd35R6V
eR1GBJSnYZOimaAetmJmJ3sbEEU3NIXR2TVI7KlRINnvl2wXJmJ7leQVYi0iFsMRpIXZp1faKNvW
r4R7Pr3QpXCrHnkPdDIFuilGrUJqFbOshMrFbmx5wz26P4iJ6P+8rAUIOHABLvEkJhSVfnXfokOC
mkEksAnYt7n4ch8cqBwBTIMEiud2Gvot4xi5JLZCI8i3N9/joHgNumoj7GmmBLOvImqFABwZc5PB
J/5jKMXsWlVZdW5/zONyyNQ4lfDpY/Lv4RMOXQo3g3JGQPCkw9bRkpoFalV5RI8AUUUh/Rf4P0lz
t7uB3PabG19etMbKw8s64qgaxD7ZQ2AILnTRsQgehPKsT0rLKlB2BsqcpR35e7B86eXsOmlzPL0r
kDDex1ir6Mlx846S5wEc9IBWJpAOAnzFEmZZKIRXc8Fe+h4Z+XPtHvG0Ugd9M7GmuL+b3aEu9JQn
55DLWepzZ1ERxuHMbeNmKbQbvhy5X+PS/JD9hUVGjjAoGvwWtiuyqz/ShZvj/4ZQnyhcPwj9NAGJ
rX8lLcUfNvEl417z0JFYEbbbKptSpMJbHP9oO7+01ml0HYH4CSvcS89zCoM+2mBZtw/gFZmDbaE0
iB/YlqthAVjnO7WCKk5Jmjp0dcZ2ES1hvnzYUDBuqBqxUdyPPEhZ7nPeiq6ghzy59DmBbCnEYmyM
CJoeW+RX5IGDh9SQ2OOKuBCXrf4Aw+Csw6ekHA+pMTE5+M1UCv08j2rFQU3iBvqi1/enbeUIJhBe
U/8B/llw+RBnD2r+2m01BNASlVCYFIIozJ2MssIeSijs8DDu+tFY8wnltMsL5Sf7Ggq7cJXWfiX7
zTiVPffyQVtPO3gk+ZvvkOG8TGyzMb7wfkRR43UfyeqVxnjzDVa9irKm09VedFKCGRZFSY2bxo/X
5Az+AGwVWEYp2JMvN1Mdu5x+fc9p99U4BvTRZrkGlB0UT3xGhsFX5Ul6y70sYiL4ZayDjVfBizu2
veUrT1Dv1vohChu8WPPiqnCe/Z72ECrpHwSbTNtC3f/aS501I9oY8bCSjDz9k6hQWEfW5ZgQKoSp
8zqY8M66sVrWFHm+DAiQ0aumDViv+b8cJOd93gcO5m3eg1OoKDayBt9lxg98iszFRrV87kZBL/TZ
X7OtIB/GUfC/Sbrczzi38vWrAYrf8XNWZt3bgsKt6A0Zx0VX1IUOX4rGbiLpQFXAy8qT+wJVN1GV
goHe7gQxYrqAJfnUCvGk2Yyag3W+aprof1r4UZz+tReTVHd1GK/0EyzxSAu4PupkfcLBYL3RLRok
INOHWsIvTgf5Cxy8IScWcEVqcWYwxvPkfvgbbRBO43liD95teRbz+EGj3jkEjlE3vgtqdlr0HaYL
2qzLVDQZo7/1EAXTVzaUiguHIUQ2JjKvsvHRa3dScnHkKCgF8yiOBJNXMUj5805FpYShAIaQ1qdE
kY7jFHk06bbCgErxK9iN4E6lGTo9bzrIr5mlpuvxoLfCRuU3TFxW7ODLUGkMQGCIsQHNVmJ6Gry9
hhlZfaQ6z+QANGznDQX5rnXYbSxQA/3NWe7CT7IlWtXbhArjkdDxuGVNmPYO9mrYI3f+iiVenvk7
tXRrVezaYJ2/IrCRr9cuHwM666yCA9VFNN9XInl5rBCz68JKcNJE/6fWddb31//YHGy+T05dHwKO
U6UseBlu8NgG5od57HCZ4vFow26S1SQACRvcT6n45I0VeuFr/njK84E35YkrPHt5QSLuN9ixjNwh
eDqB0LP96NA8UsMYnUTSrwKy5VfbdNuv+xCSU1g42LQkpCIIzeJ/NVE8gPLV3UpUfv+JwCslcz6B
LOQ0gg85O/e19ARbaaEg1b6XHBr5BQkq7YYCZR/PpKoaqjre4pFGZygJnosMfkIyuoP5m7yP3rmY
uglgbbH0J/vRCdGt4SJyIlVYa4pZW2anmhuCRWIRaJApbJb0nfyFd5p1WYoaRXIw2jsCJgpoG4I2
+3ejEOPuvNQJin+PyW3DPGpWneqM/U46jZ5Zxy3BtkG2MR+ucU6TggaVmtDirZG2iVQvUxU2SM1K
+8BARg5+X9sklsodVChBB5esCcGjXvbZA8T3myhw23XT7J1joFwALbR3tYdRdF9isD3czVELP3zF
EhcQbPy9/Hpyu9YiyYCPHDttKtQv041RI+9QVBGW4DrhY7ghQy3iliHO6981PGe4tV2lOtw2vPlN
ASALA8HLihKaMc5b9kYT+Cc9LfWCCb0jB/JKM7kF2fL0negpn2KFLC8U0uyq1Yw26d7Lfb193GJm
P50XlM7fYYGnAEREXH7BzhsyKtZAqd1qZQXKgbw6045CD6HgeuuX0FjF0TX0P8MyYZrvSWrrTQ6u
xUYF4woil+J7/N4iIuNuAtnZsU+g12DslEZS+pwogmpG69csGM911jo4p4W8Uo7X4B/2UG78y+Za
sLxez0DIPFkJzMnhs0vlA073VSJVj5WSD9VyGB2mEmMwMkR8xSZZzqOb9+zFFTtzZp+kfLZbw9A4
lXVcI9pFSrz00O4cQDz/Z2lV6TW+JZqP3gt77d/xyuTAFTi564mJA1eWnoSnKHr+0wXfHlMFov8f
NLMMZdWUNlnOy9ypf2msHtofA00SbMq8K3JXP9wrFcOiLFtQsYmuZ+ofgSbBxFcPFp8qOjp0T5ni
CC6xmNiP+nFgbl8wZuznlZ4nIMMyBkYULgLGBxLFdv4t4IF06ZhgLX5hRo3J82L2uqyiVE9nzdru
c0+Ok8CmYtYRg9+hdaOp9EwqMl7wHBxAIxIPkWKjtouPklJCJgOv4W5zV/qG+8mbwsPrEOGbb+aH
QIMPjkW6yNHvi7fwk0yFK3AgxtBhWxROneBtymNduTwqY6ywfJj+Kv0DGMgLxRsEPelSNtnmC40J
a76kcNAFg83VOTM3hex1u3Ulqg0a2+KKON4oV/+D5/pn0yQUoZYzXUsqQaY8Hm95aYXQWyaYmLgf
oWf0DySlbneSBHJkCsO91ZMZMYedr++Onq/0atZWB1xkO7ULL6YErxLP/+hXh3E7ryVPPHK/Ns79
kpAYHiwMw4zsdBEM2ue9YxQT+8iFroePQb6WU36Wrcu0eKX8IgkQbG6mzNjeIIgiuNHVnVaDR6O3
JKDjYJag1tKfrjhzXFAvK3GGMqm0f1Tx8dgpk4TR22P6znTBdKbexc6tCilsEIbisJcDa1esjCjQ
Mvx6HWEby++pvI5tKo02xhKofnkHwy/Nd2HArkL+Wq+843hXVdhmtDCIJtSLSyChYuyDKCa7jiR/
LwbYKKGP/08TNJQQrWuu9bN5Gv0pq5OeMpTOZpwvOaRh+YBT723PcNmn5PUojMSLqXBxwaxWE+go
UbkMn8qNlfVKzn3LT45m7GZBAXBCavk5Z9F/r/2y5JfLI1rJvO8+kUiZxFf1tOxTTfiFwxCb41pA
77HxoSaBLeUpX5TC/OD4utePdWJWtZxnuPp39bLFgUigEWcix2GN+9bw7XAE7ewlJCdvO/1o2wfs
EaLL4aOsf9fHzhQSWiGRSQfjv+oBF+SL/C2znxYvaBycSoCfUk7h6/ReBB+3RwZM2zaB+RCY3m2S
yxnyI3aHlOAcdbhVeSvDGV/lOuOZ3r84MjvQ86Zwh08FWZwhpCr1haYCWSSvD430WUasvH5HGsAO
O04FE7BfK8mxF+PIp1PhqpkTUMfVB6oieMumcEFBttMolutQGhthQmHpNwvuP1Kutm7sYFPZyhrU
R76LJa43PMU9IORAQHfSRs2TC7Oi5H+FYoS+s0cx1iwEUr2JFQ+xO8vesZYkq4ygZqXrhGKFUsKj
MNLRGNR1Z30yjVHMRQiTA7oioyqYghhmJYcXv3BHKucuNgv/qtbBYVy0SfpPw2QSfJbWDOLZ+wnM
qrFAR/eF9dMwhni9J/2uJW2k//qEYLIXDSs7U6E52d+XJd2XH+xekGkEx00EedvwSM2a46VPaJ60
tN/hpZJv0rORyAG4gR5OfnkzeeM8P0YaD07fnS65ep9II8icLAj62QxuOcgwwp3/MHpLKByYpaRT
Ah9ZmEo4wy03TSe2p0n6+EQPBWJ8KdYGnqFI99IJWuT14RwTRie/xMYyc1LhJNOLW8Uut92l0zc5
Nc71nqTdTuipW/W6aS08uN7FrXmGvp/w5625Z+VN1JzzNJL3GynYRYWGxatt8BodripQqAX1hkUb
U8ZCRNqEv1NN90sthfHo3KBjRCGtTJMr1+gPNwICA8qDu4ataqE0FTFQ0xe6g/UG3Qlp2xUhPFwJ
+5zf9zskIue+SHlW+FXycKo8dfZOVGkLkm/qzioT9prBIenaUdOKFC0ggTwYnW150U1PM1bX+4nC
UHJ3gdYrifoCv5MC8nSU6NdHJzluV1HdyYdOmLAXIHdnf7LseRpNOw1u5nikYHR1CaVUm1SijG9I
lZLJLRhfSqJ5i336lfwxAizSooIdzVYMynPOxdZA1aWdWmeExOUB/03xi1LO0asz9IisIQHsFlAH
Blfm82YNz9TJHt1PBuM5ghujNfIrT3cd8wiPF3qh4bb4f8XXkpqLtzxsHRw4Gl2rr4yle2hDf2vE
CPT1oGLC0YTDpuBLRFEAOgd78WEI/EeyAg9aTsUqge5sfzuKOquni31HwntSVa9EqdLMuUX8oQ/Y
a+JXZxGo7wcaqaW1//4+9cON5KUAEnANJPKSuXhxQhx7ubNMwpcLMP95tUJouM0jDc/SL4dpH6Bk
AIdD/2SWp+bAkgrfin2gTj2mCA7yf8w+VJO4UBVMlQjF/o9D+BIcak5GqN3XYy/vNXn9FP8g4KTC
Dba0lkD9GGDQwO0bd/hWDo3jOCX4PVaZjfitO4kVI5ZJv6kT4z3bH1ncTuF+j6NE4SQISozQ6lHQ
XLCTTg0QiPKASM91ObgwaxaNeWXjA83Ls4OxHFiPDbPQ+SNBj0lJRPDiUqP7EetFlwEMMteoMNiA
tSy+8jCz0VMRTY+tIs1+rJ6kJVsJXQrWuQjO5q0q9ET2kd3XBivwGEfHW6fCMUnH4SpvqF5KRnNz
5deo8SK7+67C5ftf+kDR6t8YA0MABkgoRx+yQb2X+tQgWZO+Hvq6dasp0W/BoTD0GFmPRBzcyI95
7OEnjznbN5MY5nhQZ77QrZkDfUdahtRuQQKk4/5sBa94QtYFykCHk12/EoMkHhnd1F9Og44yWIFO
eU9dqrmT2jJaPuRWHiIhO9JLexu2wXnE5RiaB+N57Q8Gy0s8YzwJOcEI+9Cp8xZwkrByZppySzRU
vQiVFKwyaGNjlGxNEwbvPs33w7qV2E8Zowzrc4HQGdPbOUW5TNSzaIrcY6VWhr0hkPuso7MyfgHF
4Jiz5Bets34Hj7sdPqUEVSdDM2H4ribsCEBdG6BqUlW7lRhKXR2SHfRBVZNMi0JFe3/h5uANLQYX
jnY2rK3I7tDnbZmXFgV88Hobi2LDMksOtmJQhvZPDCuhHReYrntFj1TkybWBPZHt6CvfteFyRtb0
qmKABH1BWagQaMATCpdpatiS0pi2xcE4tBeIlqg9mbSS7CfgQ+hB4nOJX2QXxLvMji63KD3WS0xM
J+S9oX+GmL+BWrRNiDZPMOE082jqp5XfvghkDzMg3vsIJ64+jUlwLSpKnQMjLMg5AZ13ND8CQ4qd
SFWt87Kn0Lx06vO/Dp5t/6r2CcEnogrrarhltft9y4aOF4GmU19uivNWLB2Eo8WmCzbkntUHPg/Y
r1aurGWW7oV+QuG2uaDCRufVxJJeHzjNklSn7bHE7C3g5/1XplNNU2Z6r+qMO9sMiTyc7kiCoDve
lwxCSWwzrU55LriqSjQKRDP1QvHANCjJuVB5Wz/S91d/PUrUaB8EzbYrCkhJCBa3mB/fedPpy1b9
0YhxcPKCHxZQQze+jyXA5gScg0NLVyQbndT6xVWg+rlE8QvfsVSMFtOkpk703jgXmOF4aYQo6IW9
mpMJruI9kkZnVyyPCOUp+U2qFLzNb9NidGXWOJoUhV4i6SEFYdlMqxlxO6Y2tqtfvulSjKzdpkeO
Fn78RWTvjpa6Va0UBkoDm5OaFMph7gXkSjpt0idjtZFPlun2dxu2UQSbuk7AFZSgnlSL/eMfXKbu
dSDfN6LS6Qz2SSJ4V1Ti5UWn9HfP+uwBY/P3mYJDthz2bg3DegnAZxi/kTSqSWbZ+T0fEsDIyMXI
Ub57TXXzHGaJx7WFjugvr1kVed9LyJ8Xz0uEA85guD/OyK3ab/Qpy2nsvYFF9IUgsSNfywyp3DeX
vbOW9auPu2XkWB8jUYjTAiUFDo0HOAYWTm0tBwa4MRY3johtDH9OkgVKdO8u47n3akezT1cy2m0Q
skA3Oq92C+eJ1FQLIE+SXBnhYC3whfXbQZ26GeAlpE5kUVIMKGh6TlBlk9hVg0TBwne7H/kC3yKu
1r2gb0oCdfbqQB5Bsd4i66JDgY38/lXYcrg0m+bvR1MhfWkikCMODdSwzbGImIt9jXNzUChRbOev
pIEWUrPkFo+lHYe5FHZmxPPtuhzp5MuAEZAwuREXvYB9Hk4jUgBBfo5hT87iSMXxbPZOg0P4fedz
ErrWRXvI8qpt27U0C4rp+Vc2ndcxPpgyVS6mdxCetOP67YvYEyC8zt/ZVjylvxG+08z4d1+ptT1E
Ftcr3HzgrcLBE6vy8AJzphKnfhE70GFVhIuGstR2kLNQH5mV5Qd2tIE18Q+CJ01la+Ek1xhCyf3a
XuR20zzGTvR6LIy92oFwmhXpu32zHZE/XKbDLzfi3lyiUyhRnOhU87G+tVUi637WWWpICwSD7Dyu
W5YeSH/YF+s8iYTYn1gO2mngjh6K3Pjpf8TqQuflj7Fl0VYUBu21WNG7k/K+Af2OabRKxtEE+q/b
f4qU3UpDnrk/wT9NCvvgODcp16a0jnYBhEENSJpm1HMfFUO0RPw9MizX9m42GcKSuOBykA+nA8pR
RfAp9BQ3hceqI+9xSr9QWZZsNvA8NIOZv9mgmKSNRl63D/WTx+vwzY2PPAVJbwcxRiK/2TSs6geQ
8LRG/Qhpx2bgqej4p9CQjlIqzQKbDVEOUoWmn9Cng4L8W8STj7J1Wqz6flLAlEIqppOBZgZnNgtY
rkr6EAcNOgHLa1rQBQD8xGaEidvh8ad4/xrJboRC8OlJRp3X/UqnD+QMALJnE0tP/3InluSEPvnm
vmM0JXpIKCkBC7/uStmxaKNEhmF5FPfOBBj81FQxqTpTtjnbVszwIguS2bJikUWs3kbx4N2I0Yi1
kdD/BaEHLzKPaCr+c+mbacTBjiW0dnvvqXuEb+bPfL9drlZBZXLQm+or+5UHbVKj9QP0132EaZBN
ktOdOTg/WW9rI7NCL1E4Z1eYqy+oX98a68oH/PZfokTqA5AKkPKCb/EP6bdSQVh+DFakYKdz0SGd
KoWicsJ2GS+H13YNOO6khNGM/YLSp6WVxGeho2rS3gyU8uhbL2LiZ0XmbFcSGYnyZSzaiqUkuU7R
yZ3cFFCZ3Dc6xvlh+rqGoyzJ/RmBqF8dzMb5EjYPsIlapJcfmHRVDGtSUapDTcoTRLz/cJW9SPz9
GS69cXya2kQPIf3ohpXdbgupxj+13dHZ9/crgJqAUkVYNOQkUr7c+Yjj45KxT0MhmDnkmoP9CTJD
nWy+tsR8szHl1ZdtjJ30spaHTwdEJnsd0lcO6MciTEM3GON/Wy+ncUQu5dyG9LX/38YzR5Eo2PA/
binVkHaveoxGwOwUe3Yw72gVU+1nmmdwouJEq4RMxbuCax7Ud0PEcW9tSxlYs2m4salPZB1ktvfm
6PbtrRSYH9qfcQUb4W+sQHeLfbrPV55BLnyzYhucOU6cPz2ztrlfA0T4HIHZtGzPcwUgS9BcT5vA
AopD+ed/MFboGMG3uPKWgXgGk3XxrspJspJMtjHoVkHqV050f+NtOr13bB97tPxy+8D5Rc5ZUp/9
0KYIrNgXbUDdOmt9gSwGVfBv6ZcuTHqaO3Mv5QRcmGegbxsKJy7P6lt/AUb83pCuLUTTq0lRhJ+H
8zbgMJD+LuP5F+DMfGwQ8CtYU//Bgc+0nQjhdvoe1l9i0zMyS+CUQwVTWi2CBAXR7uWD/dBahCp0
InWwa2ZPTrb5Rcq/bWDbUkJr2QRfMjOjgGN2jZaI2shrxfEZs5/oiGh79krLjOYHuiToSoPGEh5u
CdNGUpk3/1Zj24gvsXQnRwYDYdry4EooZbMz/NlJN0tROuyiBApyBTn/uonjhXvXSQIOIIm9l7j/
Jj/Q1Xz5v1qUQbNr63lOo938DH0ElBDL8fTI7P05yflVO6W7/wsp0JZUEeX+qOrUaYx5On6mX2y6
WRqzKwSao7nOmHUNAf/HKK3pPOFBj0RLVMY3Zfg7BgqwjjI4iu5SE7NbYd+DuzUOJf68SIS8QbNZ
oNznInQI0xa/xRlA2d5OQovGxGlXVlYC89zqd9DUB5ASoNO6NA0MTmxbMEsiayVODmlT66jcqowl
CjGrGSr0n27UAOKXwcs3JDOvNVWN1m55jHQAjuMdRu8MEnWWzv6xlLkK57FKNVWrXUA8dR7xEqVj
hB1C4LxEL/lHzvbroBJ6a0x8/52dJcxwPzxXHXvSKeUbb7Q2Xl6IFnzKUic5pnXyc2GDu41lcSuz
NOXCnqTSXfYs5vZizafRjwa50TJBLBbhZ45MG+LCN56jURLF0SEsNg6dcQxKF1LEA1mHkkL/12IM
dmZqNQKg9+fSeIQo6+o4KmGVc8XY/f0IKHJJDbWACpFSAQcsOK/TKmg8KUlQR9d0swJwhY85CQfe
YxHoIKpUWN4lW1C2GnEu4GwWlB5Il5RpeCyXNFSyI+m3fust9tEy+Bze6je3c06bj2jOnuae/0il
RTAFjDXONxS/GXjWIrJVJg+5pQwf4Ri62SZn/TkZI30Wpts0KXSX/q1yVm+8xb1TI5OOIIVKmypY
G2DNFIKhmAJvG7YbeSrqHm9WHwU6xslgCJf9fhMPel5wkVZYF02hksdQZsvdJ8mP9IrTMHD0sQ8v
JGtE6DzP5xMZzKGY3IfGLyxWa4892PwLKLPbCgOI2bwSeSZwcmZVLE/dhH0Qe8zKEnaVq4bbkdFn
nHceL70I1QLKbyiaZ4MJq+kb4mimk3HcLDni/aMmBT72VQDDmn6SftNCFsmlLnW0lVN5X5QkmLq5
6W9S4Wb4nLeQuwv5v2qGSsxD+ocu2dgm4S9OJGZPS/zulUBVq35vFC9aP/Yp2T7YEfOqb81Nlmux
yKa0fIp6dTgzYwohMoXx76YJWHrWIPL98SkFrpUXoikxpoYe49UnmQPcJ/sZDf75Fa7x8z22iMgb
Gk/qMqAZLUo73C/tR1r9YIlmgOKzmLL2DedVLiBQP0wS/eV/0/yyfJi8GJormatzF3Z7GUBp4D7w
XQasgAtE7Y4ocebMgZk8w9IU8EEAsiuqo7KvufbTG5vBoF5Avinw1rocPeo6swoEhbbPigEkI9rD
xtthqbOV365BTDYPvk+lI0RJwmiOs67RKlF8JrBF15oi0RJybBSsnuGLwvdGOWMoBV1hZd81NFW9
zaEw4vajz+AsnFSHa742MDV7o7uvJfn2jHGiHm3QH2L3S+j6m/DYhvtYKZXXXcdnk9C40+VlvmDd
RZtkqo6zh/A5F0Cu6gDXF0gT5wSjOS1+D22iN0c0iXv2QEFBm0xHk8luBBq/iVM0ja2Kmr2FBGfH
hXjaupTrehczITqH9+gEtJnHhrx19Q6eAXNQZF7WRJRxr2DGzmHrAbvK46haabC+mhZJdvsX5lC8
WHhx9Jp7tUSs/tt5DNXHTXwE0e+0O1+wY9EiEXnDo+4SjKVZJUqoV9qoEDbpb5bIWD/JwaCDC1YN
IBmksbEgcuX37lgzZjoadWZ+AnfwXoXuhOt142OxTcjE4VvHhmCizaI8sGo4NAs6Q5q5Gg7l1cfQ
1YRsQvWVvqVTt/Rhh/4DTF8fVNVA/obLTNpYlqHdJFhwJZxIY+LpXxVDTAUFkCxUNVd/sAz7pvUF
G+FhclBjt+T4CvvK1dW/MU266W5NodCjzT6rHRbsQBxDjfClKAGJeQWupXcRSv3wMAhNMuXKuhRc
H8RYfAHSxpKb23BYVQs+jbvOx5te8Ke458ly1eu+oXhDyEwj9nHh1iOdO+b2LBdil0MAGJHBDdz0
p6Vv29FjK2ev7cpOv9oWqITrlJ96qT9MLSa3dBfHWpqbKFFKW9hFCt3Tm6GjoetqKftRDi9rJBf3
Xw6O8Pt7GYixAhXSf3IN4lx1HZ1kZNLN+eBTBDjTC8KmXIkhJW8+fzCLMuU6CWKwbHZZ3oemd9zl
LYoFBiyBrvwUfJRsHU1YPq4ip1/ZnjkXlYWzMI6pAzEWZn/tPQza7VgCF/VAzH0YlcuklxOMrif+
wyTVsZHHmDXLG3PrHNRhHtCA92a9q2WZBVrFFspv/zmTZT6mf9UjIBICCG/ADAUZNTsNzEtQiZ07
B0dnLYXcA6MvPc3Ztph+jNr6dcojoern5+yIQAzyLyLgwO1dmDz/1RE37jkhkOV8GVEY3HrI2SyZ
7yecxwtNjqXRAq7fdm0cCQDyiKJZKZtfXrQhWt5uJhNCeHEcathLbOSXlO1qrYxwgiuFICo8OfD8
tSd2iO7PqQ5nAGQvVZcfVvNTJhqB1S9112aespuVsdOEUYu1P4BTja04cKDyd550DFahsQikDyLE
YaLw8wP0dPWKlE/pFFgjF/RA2lZBFiWIrnAyLoCHUKIcwJRzY+qg7pCiHOLgyfvSRE76GHjI3jJ1
KtUlnvrBtxT1Lw8hPCdWZdpRG3ucDEEBU3iqKUJLerSHPD20CsmVtlTTRPKb/17qlN+ZNmLZoVdw
tzYTFz4cg8XX1YdiIdfsP+KTX6PLsQoKd/zGbqOo0TNCnFTQ9k8iWJe7by3cRAPedIo6/oqswWJ5
Bda+NqAZ33sCDva4dPdlHBuuCkEh7MWaSfq0xQ4yhxJOqZfVUatwB+LCBQ2k7Cq73MzUx3n4qlIm
44c0QjYM1FCyXMQuCv9FBKfn9wO88WrQe1QAuZ3nlHINRKZUnymMQ7LKOkP8UdjV47DXOB5m6pBw
uxrfc4NfS1Z0VDHfQWNAINoWxMVW9H56X/05wVUUx1z57w7TCTsp6PFrW6VuD6QIe+m9sTlyADg5
lkXwl4Ckv4K33eywMX7Bf7jYjbNV6IsIrB27HVGepVYdZMqkRiA7OlCTpDl89q3p7cqrJ9lrYWtA
2g0iq/fqlE7KyL0ncizgTw51vJ2HIKH5XNZtzduoNB9ww65mPcboM4gwaeqPBjceXze4Uyp5sTv6
4tTIMOtDlwbrjRvt3OnTJdy7F7l0d7UV4MyeJ3kPYs7nbFuSNmncLgYWKJU8AGw1IP/uH2WGODnX
I1VYwGSULN8RnXSQbYjSKMUobYQslyDkfpht7mqJXn4tk1gw/XiPXU7EY2tKnTdNDX39yEbfHvLD
JycQ9rcUBQR1ZTlTG2cUKiz9X7OZXgVsy5xnnYfh23FubBM1mZ1hQciYVCrEhMCBbWWzTYBSmpaJ
qkgDwkiBpvs6rxVBXsOAK2wFykfF04kuwtHHG39q0f6jIdI997i18uHRcxmoMB3UYzC04GAP59al
HKyrbufDRFKsBQlORZea1+nLIt8Jg8cucxFSixmkAoJEHA3DRPMbsW+tPBiK4mlIq5hu4pX0aAs5
gNrnum1fFDRhmViS/cqZJ5/45Gp8bGvYZu8+imzgKT59hGN1Ii+uxum4eYmJq+blEpSO2ql+QJaP
yZqyKD9ia3BafObr5QJLWUqAkTCgHVDRyQEslQk8OrgzU02idENAs/EvJ8Rt85IkWNf28ThxrCMw
E2YPmwGCHw+tt99RrfOlU8KpJqc0v1Vryd8ay5EnbyRDwT66stBQzBGDUfC9AkJm3J9Br8HSLGAU
eC6CR3ltmt2GE3MMe/WX8AVpWZOSOml+XGUHM5UDZHOBwYl4s6mQEqpDexmdKZuOH04+LiZdPnHT
vDaEfb3zlMw1RACmogzXWeHIjsmBrWn1l2eBEoxjVhBCeMDuBepbzN6a71xnfeGpl9pWn0QxzNxF
OKhLKfZuZfJMyx6FHczOPCo8RUq+KDuJsJHvRd2MmPd6UMfP+0Gr+POO9SvHP+oFjQvDegED8VEa
fJwWp7RTSY9BOAAU++O+w/C7q1TlSwXOxo2se5/sARetVQudE1bmdCc3HSET4PthLo7N06Rn8yos
2EH6oA3ZkQTsRdy0Xvt7GOnT3UkJlaoJSVDpEDJ2fE0qx92481FIpKKIdD/fIF92N41+CIjuaxfw
5khuZdQvhn2S6hCD7QnCkYvvs0LlzjaNrt0DcV00UlQtLLkwKE0bVY9LddgBQNycECVUMv7XosQL
e0MT0Yq6VqmcP4pn//+kY5BOSYddFcppyF4fuOb0QoYIIB7DXv/R8XmHJBSgbnpXd/k3CF3O30Os
NhaEvqsW23SPXOf/TbofCle+sI8dMglUq4GKPAaAGVoyGyfTdiYnPWhsADRpMBFAIZXSPkgOZStS
Pp6sz88rmIJrd+6xLAhRenjWz26b6Kre4D0Vpfrxvf5afu/zmNE13z01y/iVQl+qnNibEDvrVsnF
2X88TRq+zDsr9qAEbRuJkTZHrGjREgfe83HrFQXr1YvXmTOE9lOCdcEayiuPM4AtZgzwhmlPuBvo
/kpjyGTo7OuBpCPoL5z7T4NyIymh1tXj497q0bhAf96ybWQH1YXGX0SqZ/ZKZQwfH9zatRsggOkf
mmmBQ6R9HjPjWs+moZfNBIPOHYe6b9fhaHFiFXG96UWFxP0A4SvE2aTivFUCrUl2NF50tNUi6pHl
+JjS+bRWzoYvWz4/OkMrPhhUfaHBk5GMcfHsAmWGAAdCBV84l9XAU4AdZyHERn8HlT1phNiW0rGl
HPMkYL9cyElVQxXTRVhs/jTbwXocRfWXYN6jCPgEVJbqbV6T2HmQzy9PmIbX8BjRTqkHNK9ho8l+
dVXAqpNhGWz+Ln7eZfIgpi9NNwWq7O5Lo6ktPrBMhx0rctIGRtl8/OsD5/Nw6oZNJ9zMXCvGrDHC
y6JG7z6FwXtB0++Hs0vDoti9NvKgyB8DyQG3lvgf+UasRtP/dLFkSaj2HsZWTomstyZ4Kk0u41D5
yXMvPBCRaktjaNewaea5NQhYlIz1ESpYhsjjVjIbEXjfZyi+hFb2aCbXSn6J6iDW2Qk+e8suobiX
tMobtz9vEbSiUHbNYuWv7vP+prozl4Bu4/HZmKDVIrQbHpDpgm/cFhiNNxen1bxOLDc3OPVEI6Yn
c/JJIHnMbqHO22U/Vy1EYXw4DnOtPqhT1TGFkiUIROVZjPjOLvayrRKOcFscqGPMpoXKo3B2gUsW
17aSnwND5ZTBKTKJnjhYVbyahcLAf+mr0SvyUKv1WaseYkfhEfc95rdE720YrgqzKW5BRBkbpQWn
eLsqcfGEQ8njnac015RSp2slEmMUZTUh628iGFHssEkeV19R1iH1aKdooGtIsS/o1vht4NA/oIc2
lAyidop9GsxGBZhV6G0pIz3YNoCEFn6NNeTl1Q+32lmrrzlmc6t3fuYGd+dQ/e8TBKpJe7GjQGKV
L1GkPnWyU9tv/eU+J9G5+GMcpdgBURy0j3q2uLloiyzhEz+bYaKTUP4FhRyn7UG6L2Ho6he+1PYM
ojcuKpfbthkwpMBobpWfGGCb60VG3hi5yUwpVmHkoRYhGySX4gsE0dgU3sLRnQgefKjBJMI1TL9X
vvWIwz0fxc5AWqvoDHsOsnIeoDlH96rp/Zhtdyp3SGiA3zr58Y5GUcY6HTkB7FFQwTCJzwY2o78z
/vLICHRQG7IGlLcLjkiyC5LZd0y2LVy37IUB83EY4LR97zRaYORtP0WU5+vP+cqW5bG9z0OvI9xN
U/aQcELJbUyTv0xaW4q2zW02VFJPQXiJBPWy6wqRRHmX13zDqEGVZKCd/aPGnYTFt45W3nIvQP1I
EGM2hpxdfAMja4eUtM6GPP84hbBChOoIwgeNOPTDGPiV4JyHrZbk+VxTKhVe0pNin4rnkElNZVe/
iutLV6E5JGKyhaNSnwGYX+lleccRoTsBWTC3Z7DHv5LE/wtoyLsWBOqhfait24DrJ9knzrlXy6AE
9GiiKX6yld4sIAR4Yv1U1BSC6Vz4pf50va7g3OIVRggNSgHSOiBBUtToLIB3WG3aZxeyjXviczzl
QxLgpsHM6YIgelh2x2BDorw/yHYmz82mZhridcUdisuxYtEDBQXG8zXXTPmajc0tG1YL14Gd8UEP
jgBXcPaCDtf5d6i39P4vpKVwy21wjJimpMeEBl/+nmW/UtQC7gP5MZdvqMUx21Uv2ik8vvDkix3n
NNNx2cAOMdPW32Yg5n0jd5xDlGgGTa7fLbtdCTes48B0wfZ7ot2E1nExkCfK7ZWVfvYEhAKquWuz
aTGDzQfe5Vx2pFsEx92mqiw2OfekrjtbVZ509MECcdNF7eeYQsMKSRFYAPz2Ww/3hRpFAAGq39RK
Q3Scm/6pfRHUHqGZzVozfrPmW+SSzL1C7uUPKAIs4SmguATpFwIGBqmKHusxYxnm1/bh4lpTB3rE
Y2+H5A4+Cr0kadNqxbXdOCFNyf2kBbGDW/8Heo5g6D/GRWCOtNXcNvhHJgrgzgeVE0gywEja3a9j
hQ4xAHeMNFzeNFhwxnvaKJbJ35gAFlqvdgdJYYUGctAnSsAli80KbtMrowbS/QSs2JYdat/d3wt4
dclUz7ZTer8UBrPQkuNzwCJjw0+qig5VB5KLIc92zSwL9ROCbQs2W0+d8yNuN5oTpCSStTg83+QD
GpKIjn0TXezDfWuZ1Akie47R2yMDVqStQPsKKG9uv4QPOJRSii/hJhpN6UEa1WFxzNLfEYhcFezj
UG5aLItarfjiiRIHZipFiq47Yqv4p5aazdbgS96sSeMphApsa0cgJxeStDDqw3oMi6hM94fGa9iS
yJd7V8O6pcjrt45YCfeNlddodrXlPqAnsukxtJHxf9G0W7BXPOrEqPdT3LGNjrL34ZgTrJEoML7Z
95KGdTbE70NZ6pViAiROTgeqJv7B16lF4CEAZ/wTZfBHycsgM+PDQ3/sfGKNGUtTroOjU6t1mmKc
SmvZrOgO9rezgQuF9D7a8M20eJPnmIHPZRfICM8dS1+f0umFVvvg0BeV5z+BbtXPRV4LKp8guPMd
ovMsB5p5QQQjbo4Kc9Eu67fEFwgbEJ/5hfs1XrcKisAARXLJZLESoQS3ipSXNCjpLgUOFs/uLLnk
O+rnJuql2zTxc+Bxoata/P4faUHO02T8IIrv7bIvDrUEM4hk6oA/CeYUbjm1LEvo+Fo65b5MCj3Q
czV66vGYwk4h2ac+olE555oWt/DLyZYAnABZMvx6AwcG0I2FynD7mTWTFLE984fOOV3nFpWOgO5D
uSVNG4dVMkvWC22MUI/IjLYxbVWfqMNmXC//WIm++M6/EILvFetmzTiYOFJBSW6GeSiSRXFodasE
mbP/024nnGBsk5xGCwQ5FeopkDn6nVTVyzTrMftEvzpzJlbWWhDuT6UT5HaiCVgbh99TzZXwzziT
03zqx5Qml0LuHzZ8ZSGwXWWt/6+AcjbCQoSDfxKG7dqju+SiNnbN5t5NgQSVbwgCvuDfBG5KAYDr
32jyjtQFPZpi5sOruK4Nvw9ZbjJZvoDLGV0LBKq6O1nDayb2x33cTG8qlyNiD4OFLgYkp7/MKepJ
L53h6JPF4T+JJrP/5zKBBUfNSnj2imK3VCWXy1oZue62pdCypmU+S/JcVkgVAfXEW1MoC8uvA8Cx
F83sy5aDCLQaXR194Zc4ShAGHqEewS0rcW0ywOMnRubOsSI3y/GltJ0XCHxDJLyF/pow4JHJ5YKL
DwZD4bXaz2WIq6z6C3J1PfbH1N5j8I1UUpqM9VUZMDWuqz2pgO/plAI3MzdJTxxGZAqebQPeK+3k
MAiaXPU69i9A2uP1ccECa162tckGiLfnAJ8QKxruJhKl9Nrh9doMvAaWiZaYuWOA20F7ifPDTWx1
UdsqIuqssymKoOv8uggMJAiJ074wqyXxQQHkciiJvijlok9CxzsoAUzCbbVKdMQUg/0t2ESBfDSp
gI4aaOoZ3bXeZp57oSU3z0e4yfwXllM9rDL6qAss2r8r1hEaAEvxiUQ0h13Nm9lSu0pyOyetPhkp
Or3h1HvsAr7MENRkgqZTWzkQ8T9u12fJEshWgdVsfVAQVUIhUZ+1RrtjqI9+DLtGhgJjj3tLAiWq
BD9e4igCKamg8+3MTOLBhsTtt+uIoZxIQJYJO3Vuf4R0Cp4jribxyY30S/C1/I7LtJnnkR8i+d6J
1RYH+QeCtkkInfSCaw3hUYleeaRpZkiR9M+YFC9X8YQY190ioE39M7UfbGqTh0WP+WtIB6IvHxNi
gZEAbptqZ+8sWP3UA43F2vM4NfZLzyZdsHbKaik7La7xJAJFEUmzgL4JCavYWaDKwod1zI8d1A27
koOeWPJKc3VQEZsBO6M7vRNxuwvhAZ1fkojXb/Fx2Ag0ageo0h77SFSoE8qSuhL0dd8EEDFsxzxe
f2GZJypAm39ZVLCGXQ34jD7f/nPxkWMb7fUqTytNPNyoWlBPshMiBy2TonZKS0ALdzObvblkzjQ+
VEJlHpPoztaQ98f9Ny3I96fosjB3PyD/uPxxlPVGhi7vU2/rH0UOvrUGzPMp2WAuRUiSl7g88nXb
7WhqH91dV4Pu0zQMJ0knWtqjlAUwTjWQHZiqcgWEhstFdJO2yPe3ALHEjjlETbaG1L5Isdk1vuag
I5h3hNzBo4gOVr56IvN1OP3We8Vo5ET7JW08mr2JMtLGnE+HNt+HtNOddvnar+vN3mZceGqilkg4
0DmEQtPf7t4iAGmgK3BwhuxKC7umBcElV4apgIPHipbSXLtXs53U9KD8wH/7zLuJZ8WQKUJ9ZC7i
SYq0GVU9nLsxg1yKyQjcYcbjnQHYo/hHndXDXUkRmdmXQPS7ubW1nWm2vCfwrS62voN0dmP5QOLH
r/MMEEUv5XnZNqcXrwyQT9pq/JI2yLxwBWHB/jKYStHJQbt+rqkQe2RicJriR1wmUZhmtoKX0/1L
RNdf3gBfXEk1jPf/kDMaIFJ/HLKHXnc1YAIlXpZhVZwHVB0s0F6oPc7WsHrsV83O7JeANof9N5je
JGkHT7Rc9Q6kGlySDSvLFt4nyYilaqD5dR5bKMvmBhSpw6ybEtLPT2SA8gI58Zj1xEhwNpuVc+eP
DeR6O7PqRHvimH4rNl2MAxsdhFbbAGHTjl6obNDACs7W5lpBUA404gbMjbIQgLuDxkD6q0Nx12Uo
XJeOcc6slNly6sW4GkpEN1BTNovRI20iviFmu65EOUtfEfHGDbLEzLFj/xGON567PFwyFG6pUyGd
KXwu0AwaR3y488Zori5YXRqtTGjdwwxMw1bJrlH2LvovFfFI/iaT3UWTrh00tjJn5J8yXv5g8+XN
yvzTOTHigqAPeUo0qvfdca1lVnXmPjMz7/Ys+hbZF2OHRx8S3KeZrwpWs9EO5uuAekWt1teWRFWC
b1zsVE3gApZDFBPEDTiPedwrbuia62SzQEz7oXW/XYhko4u0KqQRFy/wuVBTK6fXqfUzHilik+Cq
+52mpK3o+aeyfvFWLPIaER1WR4fpYNiV3k/sewE6iOOSocJ3eJg+Bzy1FZFxN5nN4nbGsoCiWdE7
fC/4aVm4+rg0puWVNpejadSIzXrRcFIii6uyaJFKPqK76S/cI561YQjfCDu6wbnv0jTP2nUU3NYn
oO5HkuLQSeV0yMeNduXo/WVDXz6f3P10kH9yhue0U9mwq7oO1KR60c4LhNFrwX0ViqNMJzjftJck
OnltZWwDIAwXVH+s/qpWhP0Nj5uR3MJXxXsVo9wvrdgFZVC7bV2dkS3yrlFvDKybcema5W9+Gn5M
PzI2gnGjuOXsDwWKe7jZ1ljNXGKc8HFprIiPv0tpHZlKmTfZEZNt3+AaQmt+89VmaNZ/aDNdecXH
iG1mV9c8LfplonggKRXX9TlgoQfjCZfoRcRcqBJA7RrKfw3q/H6Z8DvR7zOcydF2mQK4MORvPAE5
JpGL/k3+XGWtm0Z2Q1xTtg0swpVlFPvl01uFEOA2zlPcJdpbTgggQre53t4AqD0PYjbXrBlVCXPt
Ygx0cp0Eh8BwUzSygDj8mZHz8u/HdT2KZQSmeAIgDkjvvYXHNmrl7ysVURRCg7Elg6CgIaMBwp4F
9AVveNJxupIugkrNrM2mpp//TIlFPJ9FYI+w5sbLSBV4AvVw1uCsCjpwnGQFZxpmkGFHCT4WkfKK
ljmeBD0SghSaGhJpzxbnevYqteVj+MviD04VZA9IbkMONJY+J0TFlS2zXlO0XsXj9SBrTmKMWmkd
H+KB4MD71aU7G0ebvmQg5R0Q4pyLz+A02ARL+8ehoFZYE4cACK2ebRgsP2L8Td/zeQRDqYcDf5mp
UYfNUn1EdjICevsZMCdDvMpzfRKhoLRarkQdw/cqgSHbibXGD+FWwHS06elhmWAzAlpFGzGAl65F
0QuCaOZeGUETfHcJuH/m1i1GTeJu8DC/v5twJHGjs+oO5UAmh4Hb3tGB6GXI+WySn5LxsxduUqwp
eH8I/tFGg6YnS6ljAJaWwfAKGcRx92QWYyjLHNF95xBNvkFXZmKFj0B21IYfnP1/1CWk2bUl4f/k
kfwVjAIEodZaMAOPPnwN0F5+AHYqoCyP27q22ePgDABPXSRUqsxS9/0UDchYmWjw7G5q0kHl01d/
VJYvNKym91bDvZmC+OQUv5zcDluWBHtAfcYVjPAkwidQrEg9pYhoAveDXi5H2S3KZ/UmlIWPurS2
0uOvj/jN6OqyAxn9hagT0D05KGkHloUuz4MH19nv9Bm2eO2s1+1jPOzp+f6uA6LVZkVqAzywR4XF
ha4gft9u2Smj+f/cB+oHVhxtSdZCRc5FVyOZ546DgkFM9TMzkms80hCM22DLmZQKOT/ezwZhKt94
joDDdGUBd6G1Xnod04hsSbIhVYmJBid1vEu0mxTSHXNXBJRl5s/loidQzHkR9wEIgtA4qqw9uoDb
u1HJio1yW9xkysgyOY9OHVhAPDem6j+nJgBOxm7glisbbsEbk7oNo+udHU4BZOgYX3pcDslEDZIm
tjAvXKbDn7DckMioPzV0hkCVTFfc/Z1VG3P+frwVsF5/7M8cSpLYNKG0VrQNZnQL88rvaTahkOCp
0JQ/3+MDh1sy38uEeKLMulCXysBw9jXj5yahzDSarK7G4ccdAt8dpV3eU2CL38k/K64GnfRit/x/
rrvEG8QUD7lchXbG35/JBG6oDCFvN4KfaSsyiYeoSm/5R10jMnloG3J0j+WCWeVP3+7HvVkg2yH7
CUhIRKOetmdrEnFE5SjhEhzw/pP8GZNl7EE6va4G/m5P5BrS9aVY1VJVAGQmJlt/hHrl2LlHjBQV
eBItzlcIoji7oJ6xppGMXATVX/dJB17w4o5JDBA5LnLiQ1A4SD0xH4CBaq1PgdQNDsZm24bldQbC
HLgoTLAAc+Mv/K+N5usct6Q0h88DWZyzt6hE3dS2PAnXMRFiRsMSiZ6mfl8k7aiwKtFm+6l3VfVW
6CG001hTQdnH61SsBJ/vfg3jlT4PVbK98co2Ullvk6PUdA34efWpGdAiQv1R1he7zI/vL8FAvku/
i1EE3FZJnBcNjY7N+wvUFKVAcQLMZhqIbjpqBFs6rwM+nIv5w6ZSEEh0wN0cDOIDZ024G+uczppl
AHfbvgOnNO7y1FsP9wUs76WsjcaaM9c9OaPPLITx27tHxXjtZtaXJ/f9nxJAl2IuYqv6zVhKLqLY
Gir/joFIo2JXcntX1OBE59RHVa7oTHZVoCBYqYFgdYyUB6s1ibbk9CbYGrRlARM+B6D5u/ONt8q/
nDl2yaCnZDHabsKSODw+kgF3RXoMSGeQnh0+e805vzRX2WohhPJoj94+pjPuPkMmk/5RLLZjPRje
hURgvxeI0Bttd177b4dHBDXpO+m3Wnmc2O7GWMtOKFVPzXSjedA8L6zQpplkFs3LXcSOYCWRrdSD
XMhVmqyM2+pH6v+2wR3c9lVFpkx0pHFW2VNbTKMzitu/4TU9zJqR8yMHquuurpiNTXanJURCPbYw
MgsAwl+V/Z3MciO7WVhTEB9ur9DycI3LE7QG/JAWF3wRq4+9zXwGZpbXlXparfML2VIJx2CxGu8k
meV97nZqgXakVYUs9BLAg+BHHJ5BPqYaXSr3m1SI2xWe0mgZBGY8aqpYoS1NhP3ERjOZ95wQZKYT
BUqXKLlKU3/yuqCFYjhfd7d5Cueql9+WTG/J9deH28BbQOIj9BVB6/A4WaqnThVq2uaWr0oWPtKM
3Z5DPLCm6+UhdO4qq3WIRfTvq3cayPPkvS7zYUm3iIutb9AYGxUgHtfRBqmlN3fkHox/wPWNtM64
ggmtDna0iL78g/H1+WyQuO6WiJd+0v7SCK19W6WEqxZvnv4TRVtTFNuiCYa8koYU+52jE1TS9zf7
UzozUNzmc4dGCK3GhJ0lhqocnTd3Aw/4vn7YNT1deI/KR1dkif5prds2PwBxig99lfDC/uUuqW5y
ObLHg8jH1X0IhHKDPMDxPvsTK5apYW+HV9iZHAlv0HNLM4DIx383qu2XrU1izRucmCNB08fKqdVV
8M8qFwS253ZAFYx/fqqgEfoH3PyvH0Psq3hEEyKY+bBzFhvFAkS05NWD2O1P7CWp0liM7JOVUC98
ysBnepkVOi0uNPwcc8SoC4Oehus9GK12bfpceEg9PSnBHwn+SeD65oLCX9TPq1f5sdGn0fbRhtLD
K4pK0MuW7Bcd6xLaTj1KbBbXYgU8XrIouhFYDmG2jnsDi6I8VQ6d9PKdGGcv3Q/oNqg/8HQHrkwJ
4E2FDW2Q8m/VuwwoIbsPlV99S+hRMc7m1vZeUO21p3oGTkLdZsgnOhRdA+wM3+SbqHyDhS0GyoMO
QkXuaHN40Scz4zehBLEYrgI9tM0f1KpwEGPs+ex8X3lAvUcb5mugsz25fW5CkiZJVnB45AqLmlud
ih3RiO+NIcQwfdEbEiXsMXkSFQttAz+HR9CAtF2L4HYI+kQ7crYDCxPlt/yI6xodJ3j/N4UNJMDV
QfIJIjM+LdXm4IP7aGTJwRc77nsUy1om7R5ZWC9p3RIFDzX0e2ry/10NjWyOU4NBj09N7vjupK/Q
4s73/u6x2ONvbrwKQU6rwIqTl1KWR+VXRnMKnzjFxIzZKI/nbpR6LRgeudPGKXw5uYud5PGBZnZP
KfJzLi4WA978RHZypIrljUWXINuoWHVQn2ybPj1QzdDQe1sUnw1L92D/Xm7AupBiJatWx4dgY/HY
Da54EV9VMRhq9XcJouLLFNxXgGD8EaiONx76MHsT6AzGzwX+/MSCTCSicMbaW8vw/mjoQzMpJK6W
HB0DfAlAizn2ULUj0LgviJDYS9i+ICbNDFSFRUKQvLHrMYyI0BMuDwvt2onCqmEd3jARkzaXDqTS
CiCxUUY4GcZ2gBngzGxXN+c8XxsJxm64ovNEhipHZSuCzJzNr/7UF/naSAQ2BfkVnZpBbwTdSYzs
QBiWxvzPxi4UPvU7wHjS1nQQnYnmlSKqNGbNnerEe8Ink9DzmD3VxvJ2F/INfyDskFYYFcPXhVQo
kD1PWyAf/S9zOB9NK5iZz8+Em5USiIztxCOv8M9TgqRykoEkDPvQX5p04ycMBIn5Vc0WYkXQGsIS
JveAiWt6iCVFSfFTxmELsACIZvUhzbSZLbHLVJcTZrk6CzCpJn4/dwNTCO1o9/iSWPnntIxrdMHn
fq7I+uYp56tx/scIro2AZQtU/yj+G5xH776dnWpumulrqdq7a1sGybcY9AD7TFCN/Ofkd3GomE7v
AvLs9AjEL7n2cFXf/995wd0TG916oPbesSrVo6TlNVIfHxXyHti1a41DpQ5ikv9PemLTtnIf0wHK
922vrYO6VWIxezzcmAusvXTXOmg2D92qV3McQbaWrzbmAPeObGsfAO5Ei1JaJ6yFMciVw89pSOLQ
XeRBGQpuKKWZjslNNuZzNRubvcXpbGzZVNejA+EgH3XeaJDqjIqsDwJ740qTWBmCqIB45ql72gYC
H07Mx5yVT4YzwrnCHX+VJU7Wr7yjOvSSn5tqY04eOH55+zJnR8+2W1zF6Hb0ySuJRyUC/I3T1Kkj
5c0Z2YZ3H414tg8tDCS4u7+QBqLoFhVSHZlFU+EwYncAqC2ap73fV/sVYj8kcosOxZBvI/z2Is7H
R1B+Nk1SwUGIx3NJZuqpGhQ7imF9unDCYm4V9LSReRvnWReJpSFvqBtJqxi6wg/JVmNstYbs7snj
eha+DghhGyzk2fgU1D0sE7RruNXDKS4AITz3Ae4EAQHc/ytX1R+QN5FpjpOdxjHWAwZAdumaDUOi
NcirIdJg49tCa1hZM8AHuds74pKSgzcvWJQDjDiUzQc5jnT6PSIEnKsVnGkBHzgoHAW1gQMg2uw8
0mW2JuVeTI1dKe/pCqtIQU+yHKzbmj9u+czzqXvMlLiI8R2TMQasydOhR+KKX76hs9b0PevblLtk
TzDk/m1+CBl8bdjBC54ppp+GGEQe5YKKFVvkLWNcmA6ok6i5SYq5afr1ILaoT2gJvIBDEwK/iOeV
ldiXZF75gfqeN0/FBTUljUT4YJvO2RnMEyyoKwrJpP7YYoyPeBNpaq74B6+ntg6CqHEUqpiDJDH2
v55BSxF7gEFNdwgJDTEwKlIAqpQHQ0VV5sk7XvFFQkMDy40Ljs+329WPxNnirtKhK8DliY1usXh9
TKFGV25A0ZF6DPX7b7h00pvaLh8//0rhELwoxmYb6T3RlFmqwPhUwNpysjH+lz3rrFFEBsKLe/ko
QhgUkxo/lzptLpTn812BBxlvpL0EwhtoaLqbQZAUji7NAmWYQNT04ehKpPFINqwXZq9sQ9Q1fftn
aijgDk6+SQtXhIRWeRPb8G4ehqkrPKdKpFOYeaFbFaFNZ2uUZH7asR/k269yRrFj03KcA/OL97kw
dYI2W0GbtQ0dWXCjnLDGwYtiP/LKkEJ+1/7KB0ZAphWRKO+IjHTTgL0NvEVM9ycDNDgAOukqjX/j
pEyviTNTDEwJ9Zt+Qy4NJdCFhWB8DZx0//4QBfhhD3ymOdNaAWRQC6I59WGjEV3HOL7gJeJg6FSG
/B9H2WpslnGI17CmziZTG9S5LJA6fYNj4CYkWK3iISd2yHEYGILbzxOUkn5JknVx1lNF6R0hQOb0
xaW+2brEsUUL5g3b3wsNtSg6WZqyd6SGitjgsOhBHktudrp8h77DiVsqHaczcD4uRKaoynjV/A++
hOAQyyahgmqrsgHGLTZD5YnA31z0/Oyh1bWCH7OLdzrw0E71Whe1hdzlWv5gsr4XfXzMpHovzTrE
ZDDajusPuxAHQdV1NrvAqve2lWWbfHibQMmlb+bOG146YqKjWXUYXrq2PCcp6CR/ceSwjOJ2yM6h
BbjDophNIvYLqkxSPxUJUNJHpXkOSxkI/kxoN9cIzWMw1h534Tjr3fwwXZthKi/CEjcMZZzvAq3l
o6mRyJiQiR+561hL+fybbgGWEtLk7G8431X+niN1AiUeP7MshOZLzKSUlZHFWrFTIQisF8txhUfB
e661+Y42TB6+AvbdS/ffVO9XC/mCIWqF2EZWfAF4w+9oiToJoITFoVJLn/9/u1cCEwAwd3uFp1oE
3sthknRXvNhsDpepuYFH6JCnNK8mMX22Ptr09hZdAiAwKjVmyeRwlHo1Mrcvhh9xtg0iyBKI3Fbb
onOlxtPMeFB2oS76oIiQpVHOi1yiu4oTZCLNz9NKrTfa9THkekYtNkOn/+ph16SUJYURsmHsu3dH
18LPDj0JuHpNLhapw2f1vJTtS0jRjBjanGrTdZArfB7muZlDH/ml5BliblB748y69ZgoivmckuSk
7UUPPKl9Srv8a0USW/n6OwXJ7BoV5TBV9Sj5aDNJY1RPHkeL3R2FPKNcHXSvEuvzUTjE3dJroV+v
V9QjjT5DW0pF4iCVyBsGfHQM3FG+f/JlV0vKbl78YSxJRvU/abftPPLzvnje7H5f1VLu3LxVY0BK
ujPEKUPBcArheW9A0IvhHgBSAnJ0ZtrRYHCxBiNGSqTEuHK9xV+7hgNCQIiZ1kiJCvq4qzY5ZGAr
EB5vp2eJmDx7XM/qL9Ll+LNVmpHC83YSs80q5nsCB/KRRgSNukleo+f1JvGRQfWtdlWc0VBq54/a
km1d/jxVtLAxfFG+0ibLLunHLjWjcqaQ7HCaW9EVlwj63Fksvdx9m0bQp93xLL1cf5HhBXkTwJ6b
JnDkse26ueml0/R0iOcrMyzARzcWB4nA669CDPCuzkS7xU3s8Cu2Xd3P8RYFKaIvGCHHDUwsnqP3
6Dye1Lkq8T1bTrm5hA6PdOF6YN6v+RKTbShOJsSOx24NjaT0Scfg7Xds9dL8vViWkZQLWZ9Dkn+n
QpwAJ2a7qof85d0S7bDA9tz9m6j0mDb4bIlUlTXaukSUIdnrLh1NZoGu5KlSVACSIdI9vPiSKzF9
kFNrEpu436sgy9EKM2Yp/6BR/cLhr862pDVwqxJDoOBfD6PQd3AfQ4ovwXoAdIAVFldYOs4abtQD
ZD0vuyBPLPAHz0hqNcTJbLJnGpGvW/kOqsSTdS/R0k5gihOXEkpTV8Dpett4lrkhjie7ztkVRl08
sm0qgjMa5TjabLEA4WTK+Xf1zWEGpfj6CLMJwhcSO6vp90cZwD/Frn51xbw5yDIgEkMvPvofu8QB
BGiy8Gj5FEXq06Uxpay25TxHgPAMiUv3jB4/lcCd8U3/bpzNIawi30HirXb3DBqCgOgfEX/EttwU
hMFNuBirKLS86I8qE5l8pFTN/pYS5NOdV101lOwB6K0M0fvxiLvDmvJcCh9u/wzjNhoTOnfalRs4
sNO9l6D6coSq3vOAalBYrPFS3z9sBe6uI9LTl4R4xhGtSd3qbnJs6MsuaJIhBpSVE0qLe2DJ++O8
LCJVZLR+pj7UK6kjYHA+do6go1xrwVDM5jHQ+6lZly1W6ZPRQejNwZKvhvRxfzLNfYKNrYOJBuX8
VmfmeRnLHgyTgq2P2gH1xsd5oxo9KnzbxCE+UHkmqUcqYVUdUQSPYktddZy3pZf5045VCRp/HAMw
0qFFiHgbePmmaAw742La2WEFLcM0a/hW1ctR8PCQ9sfrcsiqz0/KdJB6JvLVEPOXmwDhNjay7wwM
2M4YO2EDDCsKI01SNBk1q2r3JfZF2MqKHmbEQC2VCubdt3F7H9rfDMv+BZPU4gyNvn8NKrBxqfPr
RZKdGKF/psgmoVCrbCleXsLVYLnpHvzPm6Shb0EKi4Fb3DnAtPYDNmfkLf9dbzEo1+E42ugsJp2b
agHstHfpNuMwpnr27qmqvPvMnpLEX6dTTMiLQqQXFXwXIsWXPJQrksgjSZAJxPLCSP7Vg8yDaKV1
tXus4VQ8jZrkwGzq7Y6Q1IfCqCYBubhMw7esMxpF3asgshmmowJSovY5LZZgWCG2t89tYYRAZq5M
amjePIhqO/eJe+B2y5PB4MqE3nrfOjRxk37m0SRvy1jqFE5qRZ9g/6dhmJvcTgo2ZPS3gSb9BHFt
+cIfLftbWSy8WEQHwcJs2CxmEP7bO7RvsB0fIROxen109Kpo0KPO8yC4NELL9n3oNhdz1Ty9QL4t
ewqpFE79xjBSVDs38bIJhRgOcBUzvhDniwsNa6DSxUTIpHS169KkBWPO/hjxDOxT01wLsq9RMZrC
mNvSsRNW5exnT4Vk1bPbmgrXE3eAIfKx5QDqvYUcu1gcf6mjqpKohUemhy2Z3G2307JOE6QbBoLV
x7E3H7GKrOHx9g3ATIAU+MCNHm7SJmdrmQwBp/20oVPEFEaP1bcakmQK6I54w4aa5iGSU2uBdU5s
bNMBmL5TN7DZhPhb46ZKs02TgR23LCNLa7xzqB0YeBktDtHFF7n2tegOZUVXpYOjS88n2Z2UKGQY
EHifBalwZJCzDasgz1K0VO2OqHZZhkOcJi2rt1RpE+htFSQGjtQTDgBBWoils/1sCayMLgZyI1Fk
nuuHoCpH6THp5gV84B9p06l0OiRHKBy4Xklxt4LflJQvNOts3/KaTlQ09UIRn/+aPMOwRYo65e/F
toWHin1xfqmDJXskE632orDHjERvkgK9WjJlzMlpgHKHK+5a75OS4+I35u1g+1ZslPKqRdsNLUcY
J53nbgsjLdC0Ryhin8G0z5inT2UdAAblcGeniUvnqxh5ayNzzktsjJrUd/kCppWYcNWt6f2d3TR8
y2WUk3eC0g/+fvaJpMYWdv293SWHSQslxb49flo6MRPwnAuLPFpRY5lZJfSfv0guTq9tw7FUU8qg
POs7WlDeri6ULNDM8a6VsfYMoHVNlps/XuzQxIKRfvKViQHFqCuSZtkqzWvWo+fALnBOEDbFUiGz
lNFUKNAMmuJ2rJGO+sWKUfv5ZHeSTmUi2oRsif0JhDE2xr+XWukL0rWzaeH3TPYTSsf3fm6UdcG1
Ih7oC2kdhDoGG7LhIKIaTcxIzuFTBqaIa5/9qEaEWGd4Lpgul6+Uy1/wU8Cviw5pzzLYlh2Jf/cG
9R+zZtRUTB2yr/G3wFlhUSy86iQRKdfNTia1cuGsXqal91orJblPWyv4BKTgtVN3c1ELwuVcXu+C
nJdgqzM9kEPvIcLjwZgm8qibj3clxo42SHjlVIojewcx369E5D3/lpDe+gj8/LpeJsK/JquNhHWL
tgbiyhWeiKMp+q1O5b44aEyc0T1moKVZA4O699LP5eLThTgWhaOP9cx0pg+q+cOBCoGaVpolxkz/
mYLwRrRuNcB4GoSqWgzlDLhnVWzkYZ1zdoVqydF6C2aBtctlg52t18tEu6q7GJXvVZpjw+6SvJC0
i8CHEijEB7jLwcYpIwxkhx/um46Q/bEW1zUmHmPWYSg+MX4nkmgUV/M+lj3AGeDyQK6YZ8UPzrK2
sg2AcQyKJlFQ20CN18eZzytfx+7sFcRJmy/l8H04UE784xWVytd91XdQDkPqeP4kbQTG506EYiOh
wHYgQc+hfDeWrdF58FMhyQ34uflzwfBOpkpodk02majotVIYzorNDhjkfWludS+/Cku1gb376Om7
RXdfZ3A5PIQNR78Q00y19jyV4zq8xp9hhNVzuhKyRmDRHXy2hhfRgD/n58nmB5SNKvJ+lIiSY3xA
LTDLFwFUI+fuR7ylsjyoAXviFGBYiaRuFH602hs9ZitfRPkvjqP1k6ey66GbwiVVltWkajEp+XhL
eQvX0yo2LEOj5crsVC5VBOQEtSwetwDcmd35FquDVP7JwjpTOcK53F+GZWGZepi2sWj8CDRKP9zN
AAf+Wmq1Ytj6ahZezEJujpemLRIIfLREvRCqiT6YFe65uY58oCMuDSyhmuoTyndfDjY89IQg6iv9
Wy/qf4iBNNWMDPb0A00YAvGAzuX5Y/WjAmhgouq4otSdd79tRJeE9EOI6w21ihEq86b4arAG6BuB
q5PlrMEnmz/mLFxddSguKdxasIMwuSReB2BwrRPFGSxlPE7w3E1uzaIOevIQwwsIX6FZaxQKcO3T
80Ezv9M8qhoSzKyAPiY1J0RmADj71vUY0cfP+Qu/r2nB0vwlDFetFJDGczyhDoyfA+qngZvMqP5w
bS5n903ZVgf3xJbrIYh9tFVLd48PmGswWj8JvD+O2GJ4mNELarVdL6AF5zlb2iLCQ+JanmBZyaK8
ZuCtdg1JfqRVbCigZ19CU3urTJZ8DAYA3su2MkzkNIlbmTIB8HCtIDwlTUM3n8U4bUwnBR+0LJ1K
QcSnpq/2I0HSVsB29ATNtOpZy26TOqKhxgri2ygYYP54gCUPuRjBsfAXGeOBqOHkRzPvRbR8G4ws
AedBOpC/+gbAf0KJk+z/5PuioagGePRY/KidvZPr1dCCZaUF8ObPaMzC9+de9uvNWjti+kOfje6E
ylgvq8pR7T5Ha78HdzMTopqnlLoTq5G2Pqf+ifTOkJIpzTxlohOdsxcyfsPUVt0PWjgs1/W7oP7D
CECVikp7k8L7eG0LiBhMwvm4AseEHwNJQwrR+zrQWSJr6yNdDFvIy6ooXbaPpN20otIBcUBOxXNF
6oEtqj3rI+1/5SDCt1aeiwDssfgK6Dn67e3SJf1LIsD65o4jvkES9ZU8kKDyteW5Vmrb0lZV5Ob+
GjRS2hLq32en7WoeJoIRZtkfseQEbQir4okmg6Ig7qRJ/VKEWy+Z0eJxIJr+m4Hkc6Dx6FHa40wQ
AYii4lG6PRzDi0rzCjwAvlOLvPi/jUKEHyITp9dOMmHB4wBzlXjLoX3QKr+tzTccks2DvXUh/wJG
rECMd+XVJIte7dlcsIy6MNYZHcDSrzyLLttzHAenO6P7Un8g0ZWr2LS+6pzZzKiTgTorRbcEAiUh
ws9ENZVocZe9zUKLU3OUrtFyBOvwxRc7fpMtPDwl/xC6TYYvRL0MOhvYfp79MSbOnIClyedJNzpJ
97WJynewVYacIvQVX/wpnNIIDLTEl+mW5Ra/8eA2bHbuD/N1l+0qSS0KyRs2BjauEgNkovvZWwSZ
M7ezc366KVTUB7cm7OR0lbfq1YtkhWr9EnP7SVynxWuqiw9cQYZBp7axuRRDb7GB7Z7qF5cn8Y+r
ocfXLrm4LEx3oafnN8h/hZcZn6MFi2mAy85dbp6wVQgJQ/EGzwTAl1nbTmoSYm/8gFAc4nseOgfS
tObuTfFRak6QVbXX4UZpmEAbQQA0h1xl4aTdlW8cBsr/umaPRSDxM0oYkCRqiAa4PwJ+TuDldJW+
SmxYcizLpjqwfN167blcujxFbGAI2BwpJeXZz0CIJ4G4bRDZ3wFPsBz/bZVKzf4BJS4pZ8jphoW9
mbsPkMvJnzOYIV26NvtIyo3bW0FMQnYBgfQkPqR32WP3LH9vacDkl92fXiJC49M15nVP27wWmVwb
iquuBfOBGfvjm5wrmDwMSOLynJYrlOqmT3mMIuY4zDHkACXvpFeiQd4T6Lgxu7rNo8xfJ749Fxmo
YXzOocCWD+Y4V66qIRO6k5zr36bY5zriVi4ORaDLvoWLursSi46Mbfr5EDD5rTNq3UlKCmL3fVoI
6XXMADc/HSHdlB3JdHpqFAiNJ8Bag8kB6/N5xqRgdT2gn+2SMAc8YiBuYi+0NHb69k47LElhVv1E
AQEK9xOnPu2UUq/QZ5gDYkC9JJT4xzAB2I754dY+izhVAAwZBY3z/SmPlbj/aQ4roiv5D8saYZme
A/BDSo7+pB233GxECOv7f2RnKPIDAUQkvA2vFKHilQmgWrnHnCqmpEYbcDdoGneXkJtmrvVJyPeO
qeJE+uEbEGgOPWkAoNdMNB087+++C4VDFIeBMHDWgN6KyXCnLLYe76/srPBvmHKeMCyAFAtbQHDf
fF+H9O0cqEfmjw6911LIKIuhCp8NqTrMnb4Qo4nqNhyac5TYQQckB/rz8nBo//jCvmVSpuuiTKKr
q1gzAn1wPUVBEu1zANW+c00hsWbUP8NVi9kLYmChf/cK7Zyvpl3ICcgkgHAziafNHX2SktleigZl
7rMWGQSlgwzgM0akRMAvKYmc2iUCP+lw/ZiljCAstJGyTWrnwHSh4DtQr8DuQRzPVCUxWYWJdrWY
You7Bp8nL7pBKYSTFpzMbdhPrqor+Lo0gjZgRNZwEeWJO6ppcDbCVFPI3Ylsv+R+9TOR0A6WCIZY
opVnugxa/thByUUvzrv83Dea8xWUrqyQZSHyS1UpATn++OeNSvYW7MHYHX4WC9mkUQ3xTZFNNBNn
DJP2X8tCXTlQ2iUoMH73+2r0iLEqedew72oaeyLKI3x4Ul+q93QpY2KrmU2LuRAQ7z0LAM5Hd+PK
H29GdMSbHKMjKtW7W4f8f8+3TPzrGCbAn9PR0IUDNHA5DfQnxEKbVrKPa0IInhQ8RItXcWGqzu6J
PBgXCN6mkPTgdzD6Q7bx4Wd7rJKMhO1NWvTuy76fX+ZTOdIoWfqCFTXNXolb1Pksl/F5P4TDuHK3
NDRRz3jMwLvvt61uX8MEjCs25EI1Wt4PMYL40WGnwjY870/Jbyisoq9O+kyjZ0AN2CjnZamsTvJ4
bJYNqnumQBgR25nkk6N5AJyGS8pIewW/W79Kw/l9moTlCIAoZRP320jGYymHAHEzTquMhlcLFTx1
0KOMAJg/xJPxvBvneH9c9Bvk1yd9IKEi1L5/hPMFAuUve4RSdHA0cQhOnBPtQAQ3HMR7ULFUij7z
MUgVWRiGXX8NGmRhRZ9sx1eQzYK5EUeqTX6zjgn8xP09Z4ozEGCYB9kpQ0yJ/e7Xx/R29AEgzOeq
ZKN0K7Q46Tr5kO1aB006/cu/inmn0NgUIs1PMRXjxihS1EEf24vbao1CQqzNmC8w+SQQfhonR44H
BA8d2FvZ5CZg7j4N0rzb9uiThKQFTsptjdDP0ByBlxPNZ7AKie2/HMkCWy3l+ceP42p6ZcomAzHk
WJ3n6hl6i3czYpQunGTFyDhEDUknNdeUCGOGS74Gkgng34MH3JZxkNMZ/LxrZ0cikDKE1EzCaHk1
OA6pdE9wk7Rv9M8kyv+ZYw4aE1gPIqBUA6kDnaGWXW9mhowvdifnAYNWU2u8yXSKVE8vr5uvh5fa
lwtK/r3pxVNNvcAH+i+82QKn+KoxqH8JQSMVAQw+kiFy/vU3XltGu1ZixCwnS/8WvFyCvYJlUQt2
6QYCt4PayagXEskxqpgt5LKLxCTANIYNBqVI1o/hDj0t8MGM0MhgDyZffOhGQODuPY55N21H1d9S
avx17/+hUcrIQnVrerC8pBx37NWwf7fe6Bijip9IrYHn+WnpYv4OgCXYdqRPqJOVMCSneqejf2Cx
DG8DoigbE381igPXJAu3Xqv1Tk9tyAN0otJr//9O3JEOI9ilsYGvbZvtYFsd+pOvur+SI8e4Fs6H
usPjSZeIbJo/bkT0QOoR+cWYTtSJEVD1iq83J5ZsRhMiqxAJ6MCdXccy2tnwv0s6Y9rzysjB9Y5Z
E/IY4fpqWVAddaJ62zol6jxNOb9D1DuEbsBvhZdQOLMVpkXSRgX7FbPXkLylB84INH7LvA+mKW7Z
fp+oZJVHpC8Eep26ufIHhhKkH/x1V/fRfBC5vtf0QsXCd10MXs9ne4wnZED4qOXJCgiD0zrIU1sw
CcwZzfhXXb342C4K0eLJbMVdKN86iqY8Va84AxDYJFaJQxUK409T4wW56GvhlQ1Mv1u3I1dY8oTe
phaMpAiU1AQ7Xpp3d38gFAqjDuTi3qsV7PxgA2B5YxOAG/5ofp+ZZfmxF6fTSfVCrd49JbNo3+2w
+fPufR5oAmaV5ClYNHnUAfsgitCPrXPBudxuoKjv0xF8/C2bS0H15Zyps4ephA1F3jmBw4vmvD5I
c2Hu5ILIUOvZa81hUI+zwykMlGcuccXW7UoBtSN8Zy8bDIAkQm9gGpOa+B5sArsHg0ZoXN3v0euh
ElHv5gHMjD+Oyh2Q/zGzZOmIXjI/kqEldiKLf9tOpwsM/23czMQiqPkqwKc8p/+3YqHDTpW1z+JA
WcrA8yvQ/1HYU55AW4ubEs3qUUfD6tRmneAgtnQth8f9Z82E17q2SsdV2h2ASBr+l6IX/WC95NRL
szINgwG576Ll9PZhhRrFgo5xspEkaaoLjPmbDBg3ruCbn9HRvw1jtVmVMxxuwqYX69D59k7wfIl5
Kn7nqeAwMxeXpeifQf1Fxbu71CAQzE6siObhqVuoXJhk6DvA9SMmAWm8KsTWJmhlRXrchnzBoOQh
2R9rsjOqYrlfjZ70ZBo+QI+C0KLc0jTuARSngBISgnKvF6O4oJ/Ob0Q21BEi+zA9MxqI4uzg0Ogg
SfeoFEKMuWa0UEcdyqlb77ZRvWFTTz5IHV3DgMrcG36ouO8ATSSShabYSlqiEBzMzw24/awhJ5aK
a9sqIiHwgXm85RdRtWlyVldFe35uhWPAiIRtIVZirXt1XmC3Yp0S5IbvqKUJRke2Kxz0Ddgq+hwJ
cRRI++Qm/G7gLU09NlLJl/mANxD35w1wGNfsBfUxlQoUWSVunJLTg3+eYYbIBT74RGJXgJ1tnzsE
HhLHfXufjA1RCo31/1Svdk44RmPdIKQy7J08NC001FXzQRaudYNtYGIc1FB39ujOg0nwCL3z0l50
6f4G8TU8QWuF5ujSTw9D1eDXrQm1nBQ+ATxCH3caR5sLxXNW3WdLDnCDv37VcmbaDbTxZcpkIjGm
yig5jom13ViDRFj38kIgezR4ov2l7SEtA0ugM30UwV3RIwCjUR9GPSdeme7OeqXS6a2LbuUOM2Vo
mh/Ih0z+RjHZ22mLmN/jxKLQ3H+b+jxHSFqGxMGxURG9MeaaaFsPAZcgr8kmo/esSK2UaW4Baluy
R7yR446edyjqTGFKnqXfIh9TyAz+ddGyShk7Ce4yaBsU/4PMq/Ij+a+FM9ygt6ykSRUElbuN9upT
iP/M8NsFY3zDTFDG3ZJ+o+9nd3kETJCPP/rDnw1cXWQhudU2vh+Fv+28frlxabKwco0MDfG0T42Z
gQ7X+uMelm94gT/1Tpo1vlOJDLO7JyKZmE8QEhQdWKyW6gche1kqiZUwAKeNCzSnFT23KAarScRs
zHFUFiHGCuuEqijf+O8UyALpbmmQqc9WYKk53KKwID93PC4XGb+LHG25NyTOPk8IRSxQOL85Zs2N
aKs3BkfLOf69O55jxo9IpY6FnGfxOITOUS333FpenIiTJhBMiDURFsK5/qIzlGgiImpHxEVRq/MT
XgcYiBss3CNmt79ikmCJ6cUYrjRk9BgaQqxFETitEsVT5KX1uHMeD1Td2qfoSZ1/hzeQmf+IzQSl
NS0hbddWA54nao/RxmeSHejBoo2ZDSm6bpjmCoFBVCvMGHAA+DZvve7OjcN9lspxktJebMCJefHC
53O1rTXm+SHYIFlALtGU3DvD2SKInZDOSZIAAcZOeuD23biiSxnVL9TNLOHX6KedE2YReN8JWu9T
5vK+nw5QkCIE/gNfPlVlxAcXom78F28sI6+9VLS8U0+IkA2XVykbyEGkBEqz+NOer4hqMfJ+MCaE
UeGld61Eib2vvmTntF6tCsoTcMimipLipn9FdoP/3LwF1scOvVs9htBClYzcgktuLXSIQ0z9oC3i
4Bm01hE544pq6Emc30QybGf3+c0S2uJAFkGJQtcImUdDQ8pvCSbvnw0zEQZmQJJROjvHXG5LzXdn
6uakBvpt3gzHxqtuBXZrhQNHkjtxG93WVhJ4xnqA+lQXV+KHM8G34R7kVF08bZhl4fjqlnzm50S2
bWtxbdd7iuvpYPSj7VYh7Ef2snjkPf0YOk5CmXsIKCqVbBswG9E5phEI9CVSqe1GHQVNkzD5MN70
cVQn36Sx18+6HXDm6Xv3mSVugnlmiN+6rpGK9t410cJCVJzf2/ZSRLkGVZMnDDOM5wYZ6c491h9S
PA0OwY1eqXouqDgutABnX2X+wYdKDVMS/KcTZQfwsOvtvlh6IJ/YRg25I/YOI/f+QZ75JvmmTitb
FLFk69IB4cx9hBLlHBa9TAlGh5AKfTCx0adlDHcKwrODeepUk9ZgAdC91Aop46BghO6fqlMbFMag
8dewS/t1M2qiJIS4t6aUmCJKdXFSEt5HFFFvnAAOzA50QOW1Si4xRSr2i9B6gxtdnqphuLCiAQWq
+DwXQVNEA7/AGVmYxA+0u5Zfqk1EqhcafIz36r4/ngPGx/D+w7Xa77EBBzLBNcybY2HzwyYxxg4Z
hBuaB3LtbPa+XyvqvyoAtkl2CmDieizP44DRWQX1ylj8x51hcXnqFt3NjT5V2t5KmrO97Zl4H6Qz
wOgxU/ntdo7rWE94zSrR/F4oh2u6zOWpZgvBPYYpIYd26vksRXy+v4fjwRR/8vqFBMz1TGHvoYbY
k/o9IKV36tTnpJPFiM6wY6xR7pgCMZEm85AfMl8hWAcf9Jb64uPC1HSmaQ1QBE02OnLnT7p2oQ/u
nFCWWOnWlIS8j83OLFWgzOWVDDDEP4o+KKKOge1px59lMQNdXDMbtpA4oHtTn+yJZwieVLSlYABp
LZI/0vb4IgralDUofGf0v/Fv48YPKGG6VrInKiM3UyG4CmBilrjfuAMjNdqt5LUlH8PygNZ7pKSy
FKFwH5IL/ZxgAyP3OtdIYuZnmidNnqe8Pei5/KovAstwl5roiKo40YmWvxV6wXx1KPQDULb1HzH7
Zqyu6LXHd/SPW2oTJjKicercAMPObqOcQVyCQzrms8pwurVJXn5PqbXjhniFfuzckyGF8W6nZpVq
hwxUoAMHdQNRycdmy+MPDEMhhX6ErlCYsmR/QTJleQz+gjnU3Et3xfVK7+OIUufy6stM73n9EOwA
4p0dQLfdWa1xgiVhb+ULtFdbB/HDnIoWyFC0y1ZAp1tSKhpY44GbxFeuHnpTH8SS+q+pxFNx0KYW
1I1uby2D/l23WjP0zTsKVNJlAGMf7s0yyjXELre0Ud2YCslK+nxRGmbzEj6PI672A3GjiYyTQSK0
pvVjKvI1YU4HlKjlzV7jt3g6VuS8b2tCg+d7YTEP7L2HvJrY2j3wDYmYg2E2CSUSxuZBJKFdpLNH
Tptr1qH2n7JCJoy3Ls4/0Q4ar6LysybAAVik/5w66yIA4IyDUwXQxUu92OfmgusVgZEjA/GIFDJL
9GliaoanOmFY4WZI1Fwixbn/ElaIIW0/72/K3+p4FMOX14Qc5Z2MXV7jea0qPkG2hUNxiAm1DIfh
iTX5xnlKTSMz+INl6/wxVbaoMS+DlqVuNJsCKZn46WgcNqBlt/2838/nIrWN37rMatm0+VtxWNqU
4Zi5HWvP98/uevglByw0W8B3ohbOGQhUSWGJBm45OZ2wPqktvr0haJfrV6wVCo8mNCRstF6OIdBo
FT18M0GFeh5xsjXNnUeeUAfX1h7HtVpG6zfCC5UniRNGokRWR4HngTVmVDQjuWVQa1wXNLgsK+Fr
n4BtdPP0191gVuCJSu3YiKLxbwD90d3+dRQyHF8bCxYcvux+K2cKv3iCxBcA/SErHt1/3P6RJId9
O+iPRxknuH16I3T/T7OkLY0pZGDn8USZyhGmWOzzguWmYpYz2xbDq7u1gfUKK+CCELrnZ4f6HK6B
hSgbs6rEZz9TG0WToHqQgu49Ta+3876YdrMqLcNnCd2ti8EJbsxFnZhAODk+1XQJKHcOHCd93mrv
I5utaEAgoiw8LzYFCrpUWeFTGlRm7w33jjJjTrqby73sFMxa9FHWeLU9LfFoMgIKScFCGWBEEYFL
D+w4qLpEm/cb6LHM+82W0vpw8LRpbzNFuWUnfb/J2rj7QYOF6oBsoqJKKCg8ZAg+pJwMJeMbEk0N
cWg9Te+uSPf0H5rl3/x8XidR+mVamghW6dxWuV2LseSGAVRsNDRLGJ9HHdi5GWzU4ButCMtuGJHW
2OIyY+BKV37r+RG/0RlzlvcEpPAqgUTvdW5/bYbCx4Af2fmUwfMBx73NGkvBCCUpewbUW2Qg11z1
yA8BuAR4TN8n80rr8Etc0JuEVID/Zp7C8az/Xl3mNhgGrb6SgaFqb+rwehy/3YhAsJNBegAZddIW
AHJy4bVZPxnX61j/NRSPH93QahQbSFHoRGG5zUzKNQY7V8rHZs5vDFziR27GpWHjOQZ/mrhqZMCC
s99D2eGn6IZuPAAOf2vMHJ2vPUka0fzf363t7kePKGIDxoYBNY8vexvi1DT0k0By3T12p2g/cCb1
H6lS/TI8EIuIEeB9JnL+u5x7v7jq2drmkQYSCNoRDe8vXv+6KmV6qHMnvk7VY9RCaVcTOlK0xA2q
kVoQmyDHMndk18EIwF9llKNAB8PPUvt54fWJlfFsOO4go9pjkFyjSxNXoIgTW6Xe7d2b6shAO0su
fmIl0nYbTNbqRzdQJcqIkBLhlvLiHdIws7VX+vVnkCRa77biXuVLsctJ3eblBf2BbNoLhyEpNh9G
MHu5wWZ1eN9vgpX18IViX8zC3WHWQLKl7eaWSsGGvJvEOhLdRjtR8tWaGC2d0FaD5H/tPTHPAB/V
RKszIbvrQJvZ5JqWB8HP13oybbYVfgWEHGfTgZDbXcvuKnQKdtma/SjpC81PVQcmoaV2Cjry3IIc
OkpBiWX4kOrph42eSn05e1TQ8Iu3+uU0RV1kelC4IDpdclVPK1FRket1fRV1IXKrEllXNFq2N3+T
eW5Ocjlremt5K2DJGLMEE2L/LicAsgWKrO4d+OmQf0dZ1LUOSVh1FVjcQuKPJeSMAmwbJJETQu/N
oGmytBERfpsTvQEbX71/QXkKQkhQatEqjQbCqFETcRZPv9/+fJjvzeh/mGgwj3LC1QK1HhwB0hyE
SuP75wC1nVGTpFIc8Va9N2c/wJ48tnMdC1u01fB6z5Krz080ovKkWPlnrphSqwICy8Yf/BBD9tGn
VwUDAtNGjvVGDcNlwZW8cvxjv4GWw6H8xNzSexhOU25j3PKOggE/KOKyReX+ysdBC93NUUoMOfjb
mIFnxzKIzGtmYfFbgRHx3Qllxfq1EkAsn3HVNeVQ1W3mmbhHVXhUkzapv9Ic8qlFfEMhA9EWWM0F
o8yYF4PqkhoON6XFE+E9XeXiC74QY+4lliHaTaV8i5N8N7jKhWefGr/z9Z45eF6eX8c1OP/qe6PP
a/qVkiLqyF4BUlfv7ieCHTYkRErNhY+474NTQUnpj08ce9sUPgQ7HSW2UXfZpx8n5aD7puPQhD/B
OBFyp44a3nez7RPKDksEYu62WLQfYM1bKp7HtAu6Q31gX0dbn7jGWskt2q7KIJKygRnEmTAk7ZQD
CFd1V8Hfl1XABnrd9ayT25zJSj7BxCLBBX7JDWvmBUwXJixXn36PxFEv3snJgDzYs6WaJBbHUyrO
mN8q2F7vYuSOo4fqdn+mlXOPaBODQqN2ozEgvCeh2eHjIbBbMvds8Y09mxfmnSEh7CRw0+rPgrTG
k6UdYgGq2ZB/2XJ8zoc1N8spiLTVXBg4yHjbAMKzP3KR5lHFc5OX7IDCTOKnC7IjxmUymxwGrDGg
zniaDOV+Vv7z5q4dVPYRc+Gh6gLrdbv/IO68XWM6nhdB5T8Kw7nhri679HH0zmpaCMfSfSoP5kMu
jHi5NxEtPYwuiasBHxSjXSCEfNR2y2MFIY/GlJb3IdA+JSd+S/MXfFxUPJeM4Hz8woXp181QWzSi
YNFQ5SMQNYgIg062zh6WDbqr9lM2qTkdCYr+oJk7dIwtnFCUBt6FLQzm0zZnwwOCyt2SXxrLlt1d
Rq7wlLwaeDEsosSy12tPnFoGQRqxEm5lgNbGrRHch169+cCpETdsBrRiHhcKQn+IO78/+bFdiLeF
LwFgHVF8UJTlAI/+cARK7wh1PcuEQhKihVB6UClWJ6NRsTJdJNMVhVYX1J6MCPNE6T+L5lYROERh
AjAMHHeFV+Wo+UiN5wASl4PpFT+/x4WmR1nS1vysGZjsc5W2Huzq8SlGItEZ+2k3NRMg9BbhSZFX
jRJkPsGRFCnWi94q0Isb789N29/n27p4kAWjRhTBy4htMZ3++/dOzxjAR6y2Rt8H+WBI+6z/oTWK
zshcRcRKVJIMgHCFI5KIIxH7+5l8u2Rs9rhK6d38NSoFIWkmkeY5SklkhTw9utUxZuyvVfRb1K3b
AguX/PSijxbaPUdB5Mab0OY4SlkWc3k3EiZWV/t1GsL46alymSPl2LSZ0mSBJZgv/1wHds2uul53
021ViWkz2Nfjd3y9/YTQRcfYaZb/cMqndQ7b5XJUI/4Z0Gm9yTew1+74bDGTyzh9q2t5ptxedy8U
vSb6z3E/Z2tM7IdNTn/J4EHgM+rHNRAZ5stm5SGK4hQJ7BzkWg1BLn4ygDctWZjk+9nOIJiT1MUv
3ORvdjbd90Qa4ByAMf4HPX+H03nT/nSMUmJzWCpCuB6Igu15OT7VAE8USj6xcD167USFjDmzbkIw
xtCJSpji4/tvS0RxJpLm0/mi7hFZQQR8n5cLpOpHSuBpvfGjVCUKUtNWnEZaYbqX65gvVjs43wwk
37m2ygM1Jt8HNspA4ihgWMPA+Dlvh1iAFC3dcISmLGGET2b0qlXBWPB2/RaBXKA0srKw9Eshzm6W
xbx5cCv4Bl05FzvFeTVxEEgkbNEJViTOr8p/JERcpnaBMwb6TPOwh+mJMfd4t3E0pw+K4psn+aTM
hsenZtuKJCPQQkEnj1KsgJxpQTZZ91wR3/ClMSrrD2VkjU/kKE8UhrvqTYBGX7zFfrlaLrwqvdY4
FVdmAAdLfgDU90r24ln2DwetkDmv2AEph7mmEYlI1y3lQ82qYnh547Hx4Cggguc2YJwwDDSYkOez
jFDd6J3FGsBUPLSjGl1+zcp2cxdcbQT0kPPVnuqEX9B5C2EPkN0auMHO19DgKIKkmqTuP/KmCVkl
ebFgcbKqKdsD2kXb7jLhK8BNwySyVGZGJxN3xVDOKLejdGBf0H7eTn97mew+XwnyfMs9IMTsu7u/
3FKp+qtpNBg9p0KlX475NOLoAHNK2EzWKN4maaswA2LRFnAjtvIKw9EFWHMsQaWJioGAHcT1Jd7r
/cU6+cVYf+RcraWWBsh/oqy1z+uHLPNb9aQMnf0kqY9M5MYmhY94V7qOFTNtPKbkzhtaZbXH+RO3
rvG5rB5KO88eErATPDOn/H3XbZUSvUdgaM1upTBzXuEz5VQIWgwtR3j5pGzJhOiQASQzEDhEmeU0
oKlIu6YRD2lrH7SvUPeLzp1nLYV+a45H3xcFzfywArIw+nH90nNCqpNrx2i2nJymD7qpUwPCf1Wz
/w2DjWxYV+bWETHZzQ9F9gbW/3zE9MWtir1QPbhH1ATCGXi1+EZ5xdL94Cz/kPS2r6ZerMFlC0yF
fntePF2o/bq2XXHSoAazh53c8kklUgNLqvl4G3EWJcKaCIoqydS01aZs87SIv6XHR1uk39AxwidA
KFpk0Dgfy43VcW+tCf8NpM8GhWdX75EaE2c6l/kc85+BroTD+OxyGJVDMqass6KwFzGkOxpGYOAF
pdL0seXeLae0Yk7BYS4G/W0tLTHDg6pRpRG5ckwGf7gnnx9tyb+LmnTyDYbzpqRa8gT9kQ3T2hNv
0b+fll/0vfekJyQqEXXvQQWYVtJkhyiWx9OLYWU5zDvjuQrbkCVoj57xyOFdUeECjMXx4in7xiXT
zDa6trSKTPIra9uHJueB3idoDvRyALV5mSbZepNP5AF8KAeLICNenPIxTuxRigWPtpB17JhkX2Gh
IHi0ibyn+fWcZomYGnrRJ74ggKLJ3WPWCKjYfILVy/16mgSVzrxOvQTDTvUbEL+cD69x7joVzP4k
l/OGjeRgClQV7SANtkrePtyIw56t0f5uZsnGE998trLm3+nekQVa/6gu2m8nrKC9ktzXMVz9ECMc
fzchpOICCaChCYv01oFeu0Kxk6E8qWq2SdPTBpUNO69xbNrqzU1qOU1CIxPs0XNPvGTWd5xyJIde
+QjcYbPL8Oc1Bk6DbXVF1Gf8M6HWHO/qyQDuC+EgCxV5GMoqNWA3yVGamp06SLGhJrjozOa+Svz1
LB3BLnGCFJ15FKZIa00cPaQ8ZaABhZaPO/GT8cMUomgOW81/MTnljmSLYYdoOz6+b7RkYJQVy//w
tI3M3gjZDp0jhMpCo2DS2U/1VsnckgYeRXinXH/TGLTNd7DGJ/k1lV1eNH/lydteQ7hXovfm2TV1
GbGtYc31HUh6Ue2KHPaILX+tha3f9Ce7Ym6zMreObWwxBD3wzzCzgZwrEVU5a0rnM0Eu4pyaxy4E
l42xDUlFN3XJv8V3GwXaPVJ9DmraPk7P+sRqdzgN03jU717YlM/xMN8G8y4m9ognvOQCNPxC+qCB
Fx/Toqw0l6VNzUOTcfXLWhgnCSBxTA6h8gnEhJrN/eDkS/NBKInN/Cu6HJXDINdfrDzb3rIobfvR
ryGw8G0+P1yFIRTdAbq8a6k+8S6IySFMdvrTlcU2luv7muPgupvNotmJNwNF9X/gJPyFm9xzGRUf
LWlILaHqXyFh7CDbFHV4Ac/xg7GAgyw/xrD1quh9EYB6gJ7YZ6MSGR3H9ZxAaDZBguikgzCPwAO2
WfOMClc76LhHsUYk/9wVUgso8ksltt//LWDYe/OK8UsBvOYUghyJZTE6QtmTLJFPp3tcrRqfbkP/
Oy0hnXfqK3INiEwdJdcWmOe0k660XOUhrnuKhyz9braoFngfomfUf5RtQuekN/UszKcIhDIuoW4b
Y3Jh9ZTXIRUBwc3tAEzUhgLAgJTihLmBWPpLUlFu/UsLDZW4a744raUDEYuaSsrwUa9GUDygxEip
AAGqA937o1aGQtE7ki5VwJCLPnIvXbDozqOtP8Q+uU1ds9vHfInL5VVLAXCTdcjbbN46xxQhGWpe
54BA0WjjtI/mHQ2fN1ZDi5+KNE4U/2iCSw4WYLY+8X9/TqBzgya2/q9606Z4G9shgGXq7RzYPjOq
yJrcd/cIFfjZYTUoEuh4igXg/bCiozE5e9LPcq91EVqoSONwS/A6czRHeLh/Zlc6udrcdtX4qNPL
H57oXA5UVOoTyITMQPhLasF9j/+/LKHv1ZimNyK+K8s+rVpurEx6gyuoY6p/GxJRvmSesbWAlkMX
CSQqCl2I+IwZ/phmgQX2Hh4PzwM9DUaS84hfA4zH6VGi9FRmUC6DZXXCqfuUMinCO015Jmkd2D55
kx0qVI7aVL3q1xROi1J+iQEQDeak2p8lQYCLhyzkQtsApjD4EaHnxo9d3g+9Glpn4tYP98UeZirg
q767Rcw+kbY7nH14CkUreugF6oe+D0Wy4k+RJBllmXbAoWslzHa9xDQFj0nSdwTskPLRv6mbG8kl
+x4ojU4wdCKkjsTPvuQRvfp3Ek2k0qjc4MkCKXKfG95rAnLiE31yCm3Nj7nH9vo3IWKUG94dz5dH
lvsQwckc/8zedx6mfklkj3N5bVpJ2R/Y1baVo3yz1PO4az+pHVZrMfBb5/acoO7xad8nAeCvtMU/
6q64jfTOuGV1SC9vqtq7Oard6hkf8Iszibv44DMizDVLXvrpm0qqAN7RKLuUBR8+CbO19OgD1Hyx
Ajm+JgpkgqEC76rYvRr0oh6KPVk0kczofrVIeBi5uq5ieiXEaZvWu0/xe/hsQ9i8O9yQ0PCciNyH
8DJ5xLVRqGO+lRW/pGdY95S0HPRSJShQsnUjV4S7KBLGDddK6JUrkISYhD0U9bivbpGVJk7It/cd
VXaz1/DuqX3E2XYRPnhwm6jFfMK/33RNJ1Uvt515PsE3ppERVUinBa921/PAr6vWSirtJOSQILg3
bm7oDBMeX2bwRDBCG3b7aUCE04J1NvlxWqDZ9mi6U4EddoAInK4GHJ3U6f8kipTHgyaH307b2vps
9TiP705b2V5bkcwop0X+zf8hVg4SZXSJwuOrVdA2mYgs3YCYlMCcWnUV46VrhWTcVoqaeU4AKckc
p9+KsgoYBj1+bCJgwMnKRKC4i/szAK2KYFMl3lPnQ0Opuqk1Zf8EuiOaqzMBP3HlnQMUsSqY/cSp
BKq3eYb4ylMM2Ue3QMikT+twypqN5nVS9xpYJ/I6tZGTFwbdth4/Ds9DW0qBUNSBhxbgYg/vmvyv
MgVo/aMmg8ocdSeVFogJY0FEXDZlvi7bceFeOmXA8h8oAeSxwdwsa+EaW1Tqgx9cW+D28/8UDep1
G4iNf1u6C2iVokYfSdBTgcM6LjT7OI+7ZaRhrAwRBJAMSqa5iiO3ZD9cquUkiLVt8lcOfwS4UZGH
aFTcxbAy1JuVfk5IOXiW4Vnjf4c7Dj1MK6Sj8rh1NWd/85abjD7g8dNyvnfJBYR34oraRwJMMEil
+ghR9X2oWWHzlsvW+e/0Vfe+Y212+8uobvK03ToF8i8hvTEnfmussDKZRLTPXYtmi2H5+ombvClv
TpvYI1SuUIjzJNJqhMDlOdI3EtpBcAggNNHAbkZH6UA3nOBvkiJ5/KkX+Q3oO924WUaWxRf5AL62
iMnFeJmtkzghK42cBwf730W+Mbl/js40eFrXAWMDLNAf48ZAPzJ1GS+cJOQ2J55mdXbywzyCMSwU
Tk/aPwLQt8m6//oeBwuM8GoFnyz3ikaHSKthDnzNYBaWYiL+3/xbC/TFsF+OEajsV8w436agYjK6
Dq3A/pJkkGRHWmMp7iKg6bpIZ845NRRZS6w8+1mjHfNw0zpcCSoaJ+i+s9l6r3DQPMQZthZZlho9
MfjALkcGW3TohRu8J08ZalxmManbb5BXMeMpAAUynDtng7S3SO5GIDHW30/a9yHTlBT1yZMIML/n
tnZgBWRHVu4uzoKcdSIOtsrt9nf6hUA15WagfcorJ4YXRBpBOoffR594NcsMd0sSQGYId9CRahIq
sM293fvxhMkUTWOoyrMmAMYgYdPCJHG5nOgEJ08EI88YNP1prK7ihc38mKlb9G+T32VxjjlRwUVv
ixq5uo9Q9NF4TpCBr+ahP+Zhfs7992lUocjkbF5ifI4rvLfPzuuvJu+uRiSVO+QJt3twgO2taT8T
6pXYlqCd+TK3XXeq6LXNhsZXRZkzfihvRNAGmCIa1lANvQ7Ub0m5PIVkx0Q3J5VVCLw6Gd+w8WTi
H85mkOa/uNbvZzYjzKYp5Zj3gxOnW85avgrWygzngx5GfAwM1GT0e84ER+nwZTM1J56TQFvCA4tg
MyLDaHuhKk31btH9yaWmDhvJqXtGQhj073DqN7yFWDNnqnDrXDdUA8PfCQqYDUjSKNKD2ouzBjKZ
T9LRZHhDGuR00NBwXb17bY7lY5PZQBnYla1CvIWo0f7WxjqSbvCZCZ5gVvecOuLwhAp06hmRgxiL
IWq+7R6fNbevlbhPVAykgZXJffKNJ381VXPNpwgZZQ0D+O8FwOwJptueAzJFnh7xZ6Qz0lLrEf7B
WSV+0WQDY21U0ByyTvYecuTQxtfPRPNnzw2w2AbSAEqSdfZvwP/XWzr7ekhnuNfFMS1KK+hxfSGb
N06hWfNcEo2fcZWXSEF6aoHDmvjLnmLxhZ5JuWKyqVIKOMwihK65ILoisem96og5viGLmL0eXpxi
S7y8tM6j++sOjk1UZqSwZO7gm6wLzyW8qIBJRAaFB2B/GrOTU8Xq3V/izytdRUpsYSrKKKImo7Cu
IkVxmjRq49jZo9n4tsxcz5PkW1IsBqUOOu7mHLXQUh7lgKGDnIqoptBpGHQ7ZcU8CvEEHtAqsW46
jMkjCG8VX/aNytRMGhn5IQDIXCHYdIyGYPSDmasUg4EgdJYDAfwjqst4OfSmnF/xC1klDhjOcLih
yCMyrwwuE5D7nojurOEluBvFebNE3hXGeZ8ozw5XV7VyN6iroZPCdzEtlswWyj0cbvFlNtra8Zjh
a4YwjjazWvWTjlzkuv7V0uohVAwZPkVSdbusp6FUCpty0twP/UL0YN/stb89vrNRsslIbpk5WNEb
opcjuldXxrmjAQSK7enS3UDUj+CZGRroQpqCSyh5u/BpLsiKnknCZp0G4FG14ORR2vzf2bOwTN/H
sbSFfiL0Bw2CXa829iiFp8Y50hILPGDh20RN/0Bha6vXrSjKW7qsrn3XNQDb3SO3czq1jzVN/L/X
8R1KFD/Z3+QhDaW1oQytrIWzBiPE7gmvDiFqreModNkb9LxS7WDdsK3hsrNSKbFguHkbMDEsnosz
fMKhD5oBNYijHlTATHb0z6sJS2ew+LdqMDq9QSGoMqkr2S5J0ywlOmN1Z3VqI1N+R733zvlzB/W1
1b4v1c6Cm6iW4ftt7kJd1VS2yDIKMvNh3pQ0UDOmIAxM2IIWRXdfO7pQiXZzAmW20x9ONb6wRVKk
GO4TcMHL/2et0HTPH4buKyirm/ImPjQeww+yXfZC9SRXiYhucGdRXFGXH0V3CBnLkS3jDovokHe5
OxQzUHrGIt8ZJouAr5Ldld3gRmJ5hMif3LsH9NvC9YddQVkqJqnWvpz+wji5zbJevUY+DQLCLl4M
1SiaN8loYa70JS5VYSsEGZ+f9pdbMaT/8DrrI3jXKsBwPc9jPuPvmHWS8e56owxJgLdoxs015F2A
hGXZKDauEHVmL1vNeKnh4xkYP7b1EBytTrHnmxvkztMwYoYw77NjBVnvFElUjhZLNtISiy/uFp+T
lGX2+MNmX4rUFikAHfbtIKw45viUVQBOpCjyriZKLQpERBN+7wUtnEw/alL1dDcYS70YAhXqTPpf
JIqenwlCO8lz6eoeLJmnnYDSB4Wypp1iEzs24XqmgEs7SR/qnwRuuFZ8gQ5vk00Lw+IbvlmAumim
hgdAs0lqey2rcvEYGiyFWbYT2Oj5AiPxet46Gm0Lxe7SkQeFk8wvJUr/Y+g5dpEmeVaOyXLxjUc5
WGbpPva7UQQC2HXyjgyKg8LCBKiVuMxgJ7w8Qtje+/m2M12+ePbrPlyBQr4RxNhVsDHOlIpX9ckd
kRVaEHZARKm6kWNLKtJVmiGW8HKrzv3Of9Ip4N+NsGYpuL2uCI9/MqWACbnr+Z3Ldb4vtXTCPYn2
EmmByF3sjzsVEXjOcrHk7rxzGomQ+UMkE3h+KOVV49OkjTeslBYmMjyzV5fE95+2FgwV5xtXPFqx
MFXiVhHpK5GqrHvNBpgJbFr+hX2jqaJmCSPZA604806O7QTnZSbvmSltchHtJw9mMACBzY1Q4krn
TFvX0kqpLqS+RkGF5DH8qqtBsTFBpTugskFt3VRuojJo8vKOXMJY7gB4vq3DX3gSAYpTHbC64zIb
p8YIaKyS6YcXZhKYVR9j+voKeH+0c+xvE3JRIy1sDoQjxCngT1Q1oXWBbyAbUoTYL4KZ/X3PYVUL
GkypiR4VZleq0HFQJ3RcaK5FFTu7VX5ETZXTPUEo2KEIqSL7iO8PJR1vXqWduSd0BuRsy78FROwU
j7VPi5QJpvWCGRuhBEivOkA8mLFRR5/HaznWv26KdD9Z8vuNjAAD0a9I0N+URpOBN+/46aBB0WNQ
Ud+pbM4rd8B2KEc1SNL08X3DjRL/HDHzbdzZMBtMQna1JKakQ28FxHZXXtiEeBBifoP/j+hlN0r1
l+YpYGJaJu4ucB9v4WB5+x2m8Vd+YpS29DEbhh4V6XinrZDymkgblJs/ZHVzpQf54OJtXfKFco1L
IFka3tEcmGqKbaKiVLL2Oym6KnKDbmIOjjp3wCyWRepawDoW2a3mbccrWJ2saZiU4v3SYwMi6YNu
a0DtemscI0QLnf4UeXekicNW461KtwISfTEr8tHdiempwbA/PvSRT2sQMvBM05MKZq9JjCLb17qA
NtcAfnaeVJKNtpEjsv+7zY+Xdel4cNUizCyxFLp8ii+p7vFKXWwJi0H15Ecx488Ft1FjGhpL56WI
+su3bi022ATeMT24wnx99zpLyUUY8+wJagmM3GGLKWAVE8RJeLbPfiT1q6kvMAj23ZjKxw6rLtE1
q2tJ04dIqE75CD/undbL0BmZ5MQqQ+mS+9EqEitTDUc5OPfnYMcQ61/Kg/06m1U4MVzlge0wSoFn
49eY5JXCNnwwkF15jQecrCQs8q6JncEsf1y4qOkMhkM0J6Q73yZF/bn2fvbaQErM/htJT4OnPrF0
j6JleqT6F0Ujp1UTyZn12sdCMofEpU0tg+3r2mWvhrvo9dg01s0YtDdpWuspJe8WUkDfGDdS4n3s
Emk9+gqQp/dc0+JqmnZIAPCl11U9qrD7D8ZeupCws1QHcd4sGKJ9Qxeo3yYR6a0iMtZxCjQ2a1Ux
bz0hyVQMk0e5ufBxbHh2fp3/7uBuSKbGfa5tVvqH9vcOHRIafzGow0qg+hWuQldihkhCw9m2r5ET
OXKOM0r2nOJUi89Cjz585mHLcQeu9Hp04tdn4KOiZ/k4D3GtYfP93hjeKYkrr7vpvI+5H22DRbS4
K3dt1ETmXEf1zVHC3cAiT3O8PbVIS+A30eNy5+gdow7Hcck1iXyPeBGSKxM2LK+55jcJk7YwF8Uw
WPdoPUNw4dVLztIBVI6vUknCQHD23NkTB7o//nqzP5aOXg/yjcXWMCTS8Hm4nWxCqKewiblIs0Jn
TzlLQawgKDkfZj5hFlzVPH/j8ONNkeWF041/S/xpb3nnQKvv6pBN0PjUSwf0VbD1dwp8BaEj+RJA
n5Qca1xymKhkOKyQ/iC4ZYwPF21TC91ecvVV773gdQkn07NkpgTeN9yNL1cDhSZnnnpUE3L4sOAM
eEhZPAozTNVIiI1ZvSxwWfPK+1C1Wb5RTRKrAC+Yn2N1k5c1Gx4UTzqe1c2lFfQ//sTHOWNtdPUJ
z84yhSiWK4dL6wTX3QpClO36RZtnVMLVPfP9Vv1TfcQ+ikV6aVTlgCcYEQgz8FvUTQXYzylORaeh
eStJjkbu0vUmY1MFaitJMzecXVTuxDFA7w1gLJ166smgobp01ZYbxa9FswxwNhauCHxUATBoupa4
Hs84OA0qQdqGmkjEs54IRbzr460PPdjquxHfhRFQyDfNGS+rdDIqDcYJCYx0tD6HzCRYMS1TwIRW
UPhGotXTNv2oRHhKk1WcKqFoWKX/ffhIxj5HJjP83vLuKsfRcDqHiFHEUpxPgldRaUn0QzCdg8jT
qNPIjIJdpXbsg/5CbxUlL/KeOi0ig/KsfUPP5onbCAUJG+V2hSy1NzjuKfxDYnmIq3OZvTshdZyc
V4H2bnNEVQAURKDRcY85C/1jL1ARjdn6M2IHqtfIUwUYfEa3pUdHor43yWW0vAezkX+bzHDgdEJb
YH6m90Cg/UrvC2dB3egl4uOycK6ZUSkKRFROfaTLal5V6/EjpmwfrJTpq8o4T6iOS9x+l18ounN1
8aberFegg0feXb+zT+e5JT6MBL+OJzLMnNe/1/3WP5/isVP2Xt2mE809Vqm63i1AbJtBn/aF8pBg
w5ecH6qooMGqZu3sT0MaCN7M0Nsdq/+gLwoaeDkkxRzFrlw1GvsqQ4v3Q8WNM21p69p7OmjnQ2hZ
KaeLEBMl7JJPOWroKZXqYr6KIrIaqXl0Ki+Ro4K8puONye99PX0qEhjXlMjSOOTFCVrXt40OKtRh
bQTD0HDyv0JTdW+6J1ta/qpTeTzEraPUgcS25eUv2aaMSuciSz8ColVJjpteye7VsI1KIU2qKeGF
Q1EDGrMeYhpQwWuQKmv7z3N2k4JM29rVaH1CCbfIey9Y/Jn9saIeK8I66UMLZhkO6rZLYBcOKm/V
tWPv3Buuog1JZCdIg/lEL4kMXgfViCNADj+BYsqUuVFut08HK7keVuIXVdacyaZpFypCE1TQR9sO
KcB+9nAqJDQn6obEa+4Np6YT2nPpWGz+9uRSXdB5AWUqDme++BAj/SNZJOhKCEWNB2B8G+vCLjG5
fzNkyzJR21IOVUzy9KGkxnA7Pg6t3QcZ9q1DFh2joKqNNjb10TgJ8Yy865QBiJ0o1Nlb9S9A+MXy
FwTcHotGWeiaYhoPso36Fdud77wKRWj8+GQ8rp5bOmdVOZoW7iW2gx3VLjneNpOH0oTUU0vkvqk2
cwa0HzH02XCxaMVPK4nMuvIgeOqLcI79bWEaaf9aNyhazcwV++DotnW8pFJmjmycRYu+AJGXS3up
TYsbelTuSv8FMvasMH0WteLl+qgJ1Zv8nh6ChuqayL0i0wwiZrzHXTNgc+sE9slnO0gAd9p4qod/
Z72syXwzgb9WjKDTgxTsoAyauKzOQcP9h2QFuSjjSJdEJRvdYE/LeXJIql5meGbRJBR/P/bBO7Rn
PnONUz4KhYL6XsVnOsnJ9TkCnYQx0V1UoMS6mrBxPygJF91MNMQVc8KqYzdxBjUNZXioXZ1UBdoV
OkWzdP6CVaKDP0I7+2MKRafuiDe0OPTyLODi8UsExMwkqNmYIMepWMZftNGZmP+rN4L6VwNPyAza
AoA96+aIIXrCzLBcNozVGO0IxFk51JVGVTZsgxNbwnoQuEaNJJSqywPku86Y8sImUC66zdg5MqRn
jnfOohxtt30dOWrREGwN9YYlVCURy+5XqQAnhc3Aj8c06xzPi4CWCEtKGk12uD1S7J+4Ge5fBAIn
apUIj3MiTKUhXDfRpA3VPU0yqvAOp8IjeRlTIa7XW2sVJEjXlmBf5f0BxgRaOWh9zZKP1bKHlqF6
kTJXxqaQglIKDO4N1TcsSaqDHP5MvAp8JY9Yo9uHeSQXKwz0B7dUPo/EnMXzVut3v4Xg18/3iaTp
Hg+yaRiFaP9GfxgJIFkPVslYSW7BUsg7UTDrQFhfISh318UL7R/GQGKhqzOMbU2FIyWp8A359ZPa
AUaM0Giofn9nDMwCSIonP4IjCEqMRrYKXO3aJkwdRXL28DYKN4M2siNmyTvIauSVjztCxdSa5Qb+
rm+l3jPyeF5ThwbdY4Px0cL9VmJDhnoQwxeoCwUCgSlDoC126i8v8Cd8FK1PeKQQu4fdGt+dDaBl
5m7ZiOyVLyRHgqC/Mf3RqikNxurOhp2CWZolkQDIARlmz7EYHPHuc/aLJbknKKUbHSb9LOKwGU2O
NDhTeOu8WmTOvuvwc71yVnIujzAU9/ZL853kq351BxUgJpH/NHfKfZTSeuFO9Tmy36CMpTE+2r1d
b9Gl7pIkCvhxoQGx+9iVJGwsLNDamudbXlgZ+mp3aF5wAGWYmq46Io6YLJ3jX/KeAJBL6xsw6gjX
6PgGwUQDdqlw4rC9yMHuyo4sbecMaNaGZESZf2iwQwm/u5PBSLgSgyj284pYZdKdLWi6Yq0NJ8/W
ANy7rangZ+ws/DxtIV8L7FkYMT7AthHP784XRRp8iC/SVKvz/CJzhAW56xiKWyeTBsglzl7Wnhv1
0zetksW2PhjweL4FK/rwENlrxJjG0e36dTvP8YiXENs7pmZNlJrS7WhaPFfRvzGDrnojahEiW7nI
cF7bIoKAdeSkvUPmyJikZe0NhebYzySzaQz7bt3FaVJ3VINgRDd/+8o1I8pO1kEvMrJDLoZJNtmY
1VISwz8pQT9TB8/0GgHrkWfpbtfxq2WOLCZnhj9ZWwLrLR3wQGHXyNMJlWboFMoDKIukpdbl7R/o
xootx9IDxXs85MTRgp5FaktdwyWSXYf6MfLq80goSROWSg59ThoR4DasEg7WwcGah7gH1ZPivw1+
onkNkVOLZZatjONZzz19yYwTNhq8FE5IUB+UHdPESbpSOIfcD174I9HbhZOUScGPVV8lGSOMGkf2
+/wV/isXYi5UGViXhqGPZr2L3L2+nTYcOsKtam4RW9yECsnq1sFz1NE2UyT2qx8IsrtqpnBVEgQX
jLo8y6UG0YWye8T+g1G7XjfbHCRdaSCIVNZh6FEOjWo2pwDGSCfkWxw1vyXbtukZplJe760byKjW
O6Uyg38gjV9/fJV0mABG13LN1w2qxDpSE0fcoOQYLcDR7Mt8LdGhqGvM8Up2qqgYH5eF7QSDn6W2
kMaJ945g5mGJKtE6KUu1uLjJ2KKk6YTjEAFKohfvBXAxgTTy0Q7wQGcS6XgwmkMCqqmyDuaCFUJf
KPcL91kjQQqQErzNPe/vFYwLSFiy1qEplZG/oOG8rJhHkth5zJYtSSwvytnScV0o//9ue1fTzZ0k
P4UBbJ7ZIoU0vMhCdQdiPyQ+WlXXYhBUtDfrn9AWyPzrXJFcRM8pdDRYCATIfj4mjww82k6eGmNP
FnoLlJGcDKqOVVlPX63NuZr5WGrGWroTFIG7sSdFZmGo0ISmDI1WPuHpJOYy5C05wCZZnjRzYdV7
GvZPoX1eySOAg7kLW1k4vc90uGdebQPn/8M3aFWbPaITyZEt2k275dZjAWwo6X8D9OOcO/bp6yHE
Fh1xfN63q/KaonGtql4KqHWQz9RgDRhXO5OKqRhEAd21vEgQk+bdC+Q8d4t5V//9kw38Kw9hiSBe
gv+2fXri3N4G7rGwT3Xvymuajx4B5+jgxdJlz4Q72y40Ug4s23HT2r1L66s7WkdE++uN4U3qPTIM
DHT7mr8+ssuaaDTNcmoDrEIOv+jJD1JWxmGFOjxYHiV/ejhvoLJWuteZQdJNJsc5v45yPuxuDscN
8RL9MvSs5E46y3B919ZhTUxZp8git9Wz8sw/A2zVqU2YwS2y/pu2qElTPVGbPvo+68f/i5NE+5tZ
1ZeeXkXM9DtCWqJRbTxpocW0SiYLyQHrGHNMVSYCzSK6UfdpQpK5cFjjkJhLSRSLmvoX+YI3jtrl
yDKCNOWJjvsF9kO1QYqs7FH19Rrm4FXQIFS15N/5/7I58F5s4ufwTI2QU8ZhnBdQwfKsJ8rdc+k0
JdCHxx2MLqGEf2Wnc8OipuzhmIydtPXz+2knYE5x53TUNTVkfh16S859vFFkgJXldvgfF6qh
`pragma protect end_protected
