`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
V82h/mp8FbHcv3//3zVZ5VW10Mue/LSt5dvjsUkiSGtG5WaH8H9Fv7j37k+xy+3/pQvfXcpqBF/k
iaz4/vETUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n4WSOWV3uUjyMD/l4IGcKD1bHONRRplCKgax9lu4YRYlORLHEpckVBvOD9geZHtnlLIjTLNUcuHS
rc4oO2K5x66eEf5+m+hNzaPYWCrVKWQI7/tyX0imMAsD4JQXzU2CP3ATsQoldRyYOQZmggmbIMiB
stLQ3uoRuVc4t0kXI7U=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zgo3FUzRcS1G0FRTCr4C/JBs44dp3dv5CUvkYU2vM2fDyGtu9ekJcjDXnFGi3Qx2X0BV1gEyWxsJ
xqQkFlu/f/1mutspkUjOMtKZNCgPGDHkGfwBEPN/xT22fOBwQJUR+Oj5KSeDWe2U4t5UJ4XXcGMb
ZV9syPFreDWYOTWkkl85cAKcf/WXC6oz+tOUowqV4nSLA1PaSrK4ohf8oaOGNVX+4Ji/w6ViTIJJ
OqmPJQ151npm7Kbt4RW80tp1OmABkNI+o6h4rwtTS1IHzM6bJ1Krrp0V+2aEmmqoZkuKINjX5Pw3
P4Vi6iUmJI0uMpdsCPr3MEC8HH4v95WCnjh0Qg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A45QQ9IEoKpoNXpmniz3AuFZmGAAZIhtA2hP4/pi+Iwurx8nPI4ZkKpYXPnn4DfH42bSsec35aiS
Ve+A8f1Q00bmFgtclspinRe4YgFesk40ftn1mzy6g6sLCNXhUm/IIjCSNk+ie6jVQS7STfOdio+z
cvSm8QQePoJjzlJz/jkNhsD110PhDAevJWb+C5fforY6kT0k7ZmJmE7btahod6wU3o7t2HM6+XGU
DDNZ5E+RLS+IiJYVCOwsdqQFDuRaWwS0k8Mk4UuDiVWtU0+QLFZ/8UGJhy2ZDSYlL/8TrrsWcD/1
Vku2N+fkWCj38RSMWEEe5TmUHSSzP7uBI6QwVQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b+wEsHDGMmVXUM545W/2toIjDItLsHFsIOyFDid8Fv6KhzBePVZlc9t2c1LfdAa6UEpdqcx5kgIr
+oVEglJG3R/fb6dRp2mvlu6+x0AYh7FK0My5t84q7uKZ6EPBxHnDds9FLGQdMDUFv8E10WtGrG31
lkto5q+L5WLAzYgiD3//MgdbP+aqLc/75XWIRhw/PfRn4OqyBU7xSBeoK9TDxBwOscUv0cQ+dauJ
dUQ0W2ZCXwF6cP5c47k76Ikfu69J0/IO+FTLKMkjAB7Wzsyqbpl6RMVdJ/iYscNROh1xxo2k+52w
4l9VnVKN7wTWZdW75B3V/MsNTrKb2I6dBdveDg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyn/owx08GdB/M0CwlYM5XwpK1DLRGgNdNGvCa53fvz5ftb1LM2R7yhWTTXlm8iqXlg1S70wvPmw
WVO2ZNZ0csmDdQcX4HNMiokrI2gpR08Dk8n3nzdOhqyFyh79/eVJzQItyKMQmJZNCvFfww0mtX5K
FbNe2x6ria5jEBEBp3U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J8WwILioFJtk4e6vNsFHYZhWTjvAMbsqHcnvhYKYzsY6fpaoYuWnjTNNNxS6JYZj7bKOFgPjdnBA
rKaGPLghV6UU9fx6UcBVLjNOj95AU3CZPEjWGC/GqjGRPxOkhGtDka91PZuOBRTBqJT8F+5qIgQR
vO7WJHaKezpaUm2zbeC7+ShM5p4Wm9L4dzJ1OuUGZNm39p9FbORAZNzAWa35wpfJ6PPOgATFMi7Z
sN0Hg00oxMFCKSg1bxvN3p4iC3rVT+wV6yuzOecq97B7Fu+tfvP+shqnUhodTpF0WYfGWHeK9ocM
Mg7nt62XJybi4Tm5rgYGMIIM0i67934etK5Aig==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AF8EDKLpUnsf5U27caIfzjHsL1dKCT4FvrlOxjBwD3ZJ9vsXwbWO+EJTOJOFymKnoSSFnuslr7C8
ZCAbkJJLJrLXJwfvC9hiPRksxuYzuxWrtwsjJd+5KWtue3gL5kHClD8Tbo/V+Dnr3gvKzMRNdFRz
i+4p8dC6/32xR0/NITJMYT1uOYu0oBFDHGLR02Wn4PqghcTR3gQMVeL0RsDhJibeNnf4Q0NsKqCF
7OscDpis6r9ZAFao+mdpLGI93rreTlZvJBUPh2RcpqOjL/8IUv0iM922KOCZ6j1LtvD0igXehvHa
5hOx0DDcMjOoejqJiwIqLij0FB13lDBsu+fjWw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10496)
`pragma protect data_block
BMP9G5RAk03qFRu5UmzfhNOOXDwKJgxZfoTYKz/V88UZr3fa92qF7rXs7/eckNewUxlzrNjvo1zT
4g5opuY+vW3a88R8mQc1x7I6d4Naytx5g71mwuvh6KS0mH/P0lIxy1WMoPsjrEIkecYZzfPCQOv0
SL9V2E1j4mMz6Vv/fTMBhGTzEqS5xhwamjThXm4hSV55xmB4og6Vl8ekhdw5L1/z/HHhfHJTZs42
MF9CruASJbfJCc01fE5VKNIV7hPMacbKz2v+U6eNGECGuwJF+eGpVomN710lvDfNZSN4tX1aOeds
X8oChKq1OP9ZGUvsHZGArt8Dvu67gogQtqel0gB1LeshTWWPPzfg1McvXlF0NNcwZWsi6y/2wUdv
28/p0OaQtIi+XvtvLYpQjMr2LSZ7PRMyszToi4L6J9lHdfRybq3dj3VvU71XEFrWm68KkMX/YjNF
uPopoL23+/wseQvdMabzYV3cFSEIw2sP3VVPIvMkg0EJiOgwFQm05MYF54UzZRTRlEr0ToSjL9dw
mByxNNiEF4sM0DT1QfnpYnqoLxc8+aELOUjMqrlpq7/nq/dlB9LQVOCYHf15SldSE9lsXQ1WsPpW
xS7JpgqN5Q9Fa0hZL7dOLuD82FuCv5mJaWe0EVmqLirFzHp7tHyGMGNI5M0TmVl8SIZvgadK8l65
QZYBs/MZb93DvdFHtfVeKprjHKHeRN3Mvl+RG53VLPXysG55A13fisAKdLTtNWiIvG7FSTft94NT
xaxlcydUg1t9B4EF5nlQixYOho7n1ea2nY6nkqxj/waBqebI0qMXr9aIF8scPXyURSRlEh/QuEdB
W+/uetonnXn8Kkq0OzJK+eeCd+aNL32nGdMSrvoCFibTRFwpt59yeFIzAmf3yPZFU1i3lHzEOAWJ
FJODdJ+Wfob5O7+9RSfdnvAiC3c1gnuY2YtW0NJy7JNEtY8SM/iIhjfTw2fdg1J+U7l4RZ3h3uic
uLzBY9h2oEggGWeGMrhm/0TNMS6hiPl13haDZmCoWlLDLJHnwKVI7oM6NPH9OVQC3WcISZCEHASI
1u20JoHRLkNr8DhilPIrDkcV8FljF1fKG/xtBfWyj5UA1inxgwg5oKayHN0RYGO+IUczZxj/+LTq
ssLW4MW2+oKvt0yWefXNVQ1DBIOFe9G9rWoBYbSQ1eEy/KWxHIaVcPUrthxqsrHtG83haU3y4x5D
iEQlklYrERTmm+5O9d+5evOUZbBhLlOfdZttlvityrYP/x9XQjMh2/N929MuvGSxJwiPVSK3Iujz
7wHnp/gGTJSjSMNJXrvGrCdHYopnRn4YsYHnDEJDLo5V1z9eaGXiAaNUBlDb6cfrPGR3lXhT8n0r
MKMC/hQiB3gYrLgG4mIQ/uLAoGUNzVeZNG9nJRhmBehRoNaW4FhSGMds57kvJyuxIYB3A9MqOIo1
DFowdSjssLICZFVboDojMlPM91g/+ZjrvwdkVcxlEnor8KtVtLFmRyqOkSuv+dWlaSZzMGlgGDXi
D/oq9gB8Qzvc2uzEV0yooah+NxBWEr3WYVaxJa60cHks+VxlFQTkf4rh5az6I0o+swAxSt4Y/ynS
i5u/KzgmIfqNOrvJPTgeVlgyp1mzU/0BIb9Ug4oxtQd9ZfIacNM1kUVWWBVGerdR37TR8Fm+IoNf
Pl+GbRxTqti7C6bNiHVxpB9NFueDtGEnrx8tx7VfXzHEErOwVjlCVb2M3Z1deLVP2EKt6XiKeixy
UDBBmKSGHj6ycHAWr1vqggUKsGM52y6vMG8fI90YWz0teWUuFnPX6KZK5mEDufwZN3RAOXWyzbjI
fkdzbN7FNGhAXsjJk8shxWccqJQ6hZfKVsCxk+WVR6adXgjt/nM1gDIwzUd7nuZfesyEW1+1rQSb
uqp+eOpCAulk80VWeaPaec+Qad6UzarZ47ieS9CVB1myWQpOrWELuaQv1iy1aMi49u6Gtra8b4uV
OlWDfR92GggkMeyyDlorzOFTEK2wkkXhkCuQf+onIHId2+wrUaGeJ0iqRnEaZKGIIV+24jHdV/QX
P2Rxmq2NhXUOTijTUUXGngZ2BprR/t2FMi/PJWLQSHkeA+RmFa3+NCd52LxBV9lcIXcyFw8Uoqx1
e128eEkAFL2ATcYNQ0alkaqhO/th2vVS4Yk0fD/mAMLf0P6OmSUSxhmdV1neHc80T5QAsadQNRfB
AlAqs2TCKgfmECa3HTpdzkwNWyIa1T9/lcYubd5rddC58vdsHtP+hOtQ4t4lr2UILqb3UieGdwCq
9QGosShYsLwf1fKMArsiOhx450fhLTKGd80MHtAiVhpUAbXD+7x7mqDjALZNfnofb8Lxs8KqzLiI
YIPIbO0JZZXdYcn3nbWL2rU0/eQwJzLgdI8qu9CzjuCjBavdhn9nb8wCyCIdIR84kPN+AtdEH3mI
0tSftOlaVi288hgIquLDgmQXxd4EUzPDARkHyDSFOtXPtY4tI2lwG+wRCGYcAiq7Sv+r/+uEQZ71
pSW6FSDo2rXwLQmeLaTKJEOQ6VqaZxC4ug5/BKkxYZgZRM4BQOBD4CU9dVez8l6KeNQLBYs71XRU
2dKErh9ik0MPP9Hnz4KzuAeshtvzrkeEBDadTu4BMNVvzrlCcQAIm/Et/rddllXiAlGvRovXhq7r
t5I6MLzRLhm1ix18Dal/bBTtIeKtD+yz4XFEdLBLpW40x95wGX0fhPyRT1SdXphx/ZgN60XNNh5C
hwIb0cVOgvhkwab9N+g1nBkZYWZ6T0/ZZ6VnVNHm2TXM+OTRF7ib5I1ODQWjHdGcWOH5OgL6PQEQ
1pRUFuKcaxZxxPW42rIF9GJ8OLRiFD/Fzt2+/m3dl4M0Pi6D8oe+ZtaIHLInFCUM3N0IHeM+9dDR
MTl4faMBu5m3s73XMswKhpqa6sdlAK4nEQOMbELSABPiVrdcBrHrjZ4HCa6lL76pgKC7fcnolwWQ
jxLG4DlGaeJrWJ5uIpSddjPuAjOVoo2cK7yrzcPabMMKRm0UPVgSd803tgL1zjKaYwaQ3MVqj/tg
jQsQSFvCh4AHv3+c3+qoBNiAgjSaZyIG4m46NWh0QYHoocLtGPf+Tr3QwlxY/vUA9FAkngPpwzSF
WtGCLa9FPbqCyMr9KeKQG1apM4s53II22vp3AjkbT2pj1vyBWxK1L3HCH2VWWfuLm+0RQflV0i3B
3+IlwrlaYaLgomNLpKM0hmsUHsgqo/RGzoa0ald/OMvcK/KlMoLY3XdTl3NQyRdY1kFAEOt9VWy5
1je1QkPpd8F/IPE1x36yc7a83HT7Z1gN7/wEW8O4Q5mSw1lTZkQDIQL//n9BTNH46uhgqc/3+gob
IL2Rdc/vy+Fc3QgK4ck7KppLwi8A5dot4XvDfxyV7EK9Nn2s0QMOr8wEZ8teV2q/16TRukzuO1/S
TSCWbUVHP6rCSuocZTx3o0SSGbUmzQf9+iVMlPPgVYZcemv2NBPySQbzofSLmNHfzuaypstaFvO+
DP+tCrnmtL3reMCQpAocfTAKygXaYGd2zxr9o1Xi7khmW9SSLm8NmSe5EJzK3HIBhqJG1bQzDyhU
HlVG9wkpL0IXnrVrF2VcrXZ087VRKB0vJVjNuqaSWSeCmZqp3cizJXLM6PvV87LRadY3QUI2Kyxu
8g2TnAN7OPFkDVF4Uf+R22O8Aov10HoETJPxabtvIMMm963G1v0YRz6HYvvGG+6+dukC4ZW7IlGu
QksDNngcf1+joECL6bKovxPWSmB9FjQ5l+ppYp7WanDVevLSamx8H4pFgiNJbyNNaYDtIKhMUpwG
0Ft1u8mcfJ/0WWBOESizEM+vrvvM+Fo7Euzk9e9CVI3oIcNOIjTzY46HGM/zi4+Pl+5i38i7EbnT
obdUkvsmb7EBKHI5PWlt12rUYF15oHv6ypsW2nqChocTVhN/oF7n9klbQSGsAgY0BAC4IB36j/C7
sAgQOKt/E4YnOUIc9xsHjLD3tN7sErO5OmMRiyrU0Nrjbh/BTUb7voqMAwykOpzl/d/nkqRwkOBd
wWGae8vHmYEOk0/I7s0hAtn8lmBUhyCtR3bSUxnvfpo8s5eRIfbVhOwWeuu2a4TgHjM92cxDypxY
DTAB9ja+8LwU5qrjNYa0VKvn4sKp9JX+7LcCPctTS/ggSImTnVMVvqWp7Ki+rUALrtl8p4aYr+HE
rYQbylOnFrItbtFHavL/uZd/vJVPZvg6cN4KRGQsTm9MTlBVm+PDHMuN4J8Mo+mTOb1NTPiK+wCx
48uitM6Kbug6zD/ikyEZiJSAi+JFPIASw4ngiaBE8zcCuNTndsbt3txbJUku+p3H9RlzK+jeEN6M
AJaQkzWVLW7bXaotA/JXzU1zkYUKFeWXTeJCxt6CkQpyhN7ePPd4djJhzGO/pFeO3ujcRcl4TlE8
1/Nore0DBox/SZQJP3dBpL1lBIFG/Nr0ZDKyICd4A3xo5bA5kIoRmJPylsfjV2XkYUrYeUnQ88u6
e45IDahUBIPb9EadxPfsawRslB+ENf1MT/Vb4nGknBcEjiNYvxRVdeyd5U1T7FvpnvK/0bCMsPt0
1c2YjGKK8MFDKTRyvbWveLKfTzBofE/2+TgqneFjn/CRG4ScakSTk0jKf8YcGfy0q3WwT0q9ZREP
rxor+TDdwA43lo85u0Z3+DuSmscfWROVbYOERYByvZnLaraRvotlSpyA2Vg0ZfiJCak09naE14Dd
pg10eLfwh/R/T9YRB/j977dc11wut15aZsnl4JidzG/YPAntcM5XoaBvUFNVuargqGw6qr8nfEIK
ElPQ57OCsJrNUmm9E/u0VJxDQp/OTUM+zmTPx991AShGIy/LpjMWFgif2dpO/qN4SzYTuZqnlc/a
7TkoiMM6xs1IB9AHVqk8dYtPsBfQBktB2bFdl9uEg57YhnwD1mg67XFHfI/jyx5HyYnbyZADxyc6
ZDYQVyifV4CLkhRIx3ZCZPRYjpW0hQS3mxrv0UQRIL3AYNBbGBPJbRi8B/5PBDTc0t2hdCPsyGRj
cDrywf0d372NuSqh7pM9SiPt3TRl/8SCFZT1ILf6CNhWJ/uswMxKCPEqs8RqtgNGwP4dsd7ceeca
b6/71Z1b/23jO5xs9BHcEGt4QG/s2z1RBsdnS8mOmZHzasT4lGV/QylFzX63OomcrFv8E/nQEhie
v8B5LX8WBMo/nr9NlRwQbOVi+2s2EbZ0o6OTN4sN2svzszFAyGyLOxvoRtRZ8e5AZvtV6gchfOyu
RX1xLG8GTGkb9gwQQ2Dcn68MsgLSzlCisXAsZnSkgGIWdCFrwf4HW/Q8SeuyGF7gUAPVbfMrbQj8
FaF7fljzpAgMR8w54YP3dsymlKgj/XN7HlXYGKcIT+gQTFYgHTp1g2LUCTeZrjQphu7+IFvIb8DB
K3f7W7lnk1X784uXwsHstPgmN+L28NhA/F717AJiTP0dOfRQ6e9AOoYuf1tzaovtC8Mqv5+1vc/c
PH5bPMyVUJGdhfjPafmucQVUIbuB5mIA7PA4jlnm1RxhFsw1ggiyFd4JC0EDvTE5745WcH8W2Dq3
CGPZqQVUnCcCsoQdscrekaEsJY6nsmGgqFxEGqhYlF4u1kjjt6tGf8RenNrb+GbpFtcw5fBgwYyC
rpqe4oXNfazJtQffVhpMuhxpucmHbkvcSbPeowpACSfOIHsp/aSVX9vTCKd5Q3XKeM3HIDFidCoG
t++Ct+Bms8NJPk/aQs2pHc6FtcK/8jDi4+s+r9ScQZ5RrMgM1XHJNpID5UdjR23MGg7nvNetw44f
d+qUPrzx1jiOE6/EPUk7UtKJeTLZaGOpc2P222cFBdPLXXy3ykj7zZx+wNto1rUZdvcVSehIIOk2
cLXss4eWJncyaOOeOMTUmHCRB4DQCuOxjsx9tUaGWqsXNgotj/3qvt2Vmhg/yGONOv5OQkQfUJGD
TVJrHBPPSnxGcldGKTmXV6hnpD3V3s1J3u019K3inIlfsPyvGNjuhWA6oazoHMX+I51MNnIw0tol
NkI1+rejmOspbsyvTA/6imYQPqkp4yl29RpmUbyYv1rMSrMy/pw4uxNzEoZ06ryXbfon/LnL0P0d
l9DXS/XQ72aYpteP0PPtlmXAaP4NYpxIkkYopGqerAaGX6Z92E4KfA73Kt8CqXECtwF8pjYoa1T9
u4dkbx3ejinKIclCe6pM5lhnc9Vb7P5T2ckkKI4r3GBQJuxdk620zWTH9Cc/M5N3qb/jdokc4R6q
C18bpknDjbUzsRzwbB2wpuHRg4opmM8M+gwgFLeHqY6lg0UdasqIEG4JXMM83k7Pv4E25qsjkxBe
YV9Uh67FbqFOqf/GVy1E8xxGN8w5RM/6+S6CDzSBFKm+U6XA2kibK6LrdmeOYA6Ea/4dXzbo8Z56
8nzq1eBdFy+BlP7BvyhcfWF9HqjXuOnuSAaOAx0t4ZL668sStBN18T4dDa7prJwJWC64M5gOiLtA
5Uspi9nvRRTgd/YU1H1m2aHyWFz3aNHyRbnBhl5gu4l+tGIAwUMcB50i28uu65ccu5SljooCEJFi
kLYlzp8wDj6XmjUDmub19Xx5coA/VjMuupMuUE7KGETSseaZG7/eCrRWeM8UoOD0+qNDk9tSY/ea
5AUcxjY6LnlWsCUIKCqYRB+syZadlam6MdIfxo8bcRG6l3xZNmISDEPDHQtFL44jP/BjiRc4/HM+
GCUAT9Nf/2jPCmKj35VCfhnki/W0zr1fX3HDqL/W0LB8h4z91tXJsHpAMwSj/0pbXgkvkfTmnL3K
j+vdlKp3gHBMa3mBpk+DafH/hYOTdzUS3RG1+tIX4mBKESdJ9XjEUO0cLC1TJxnVrZWxEEdRK/R9
5w/LK8GEPNDqNaa+kLvm9HbZID6wKrmjxYQEfWfQ8JMAS/tI+iYYNc0enCR0jDGKKdBBuL0WPg1J
/zdZ/NqLo11AgoO0HnNmEHW6uKl+jHvhLjezCzhO23j15l3oo+J9ralIIFwxh9vqaOuLBCtd6RB5
CwHjWpVmooLIUXHlbPQ0783DYowNuUhQ6dQUhAZ6aT5bvNmrXW0vrV5+z8v0+QHCG0ve4AKiB3w4
pN7hD/lASoZq1U2jpzRYGxljO3LQSIZsb4i4QqisiOqfrORImeJfFbU47lJpocsbG6OTy1RDvcvN
ijDcl+OCtO9LtqHt/ionef1nl8ZWO4HgdvFmgvMFqTXn5beY4L4sQy2TLQXs8g7Ftxnk/B4mBLiy
GP0B/PTYEBuHl5rCvf9Aesom3yz7K6sBwBgbHb//CG3vo4glOLdZboWT1ZSJk65l9DZEsSuMoRNT
mWx7N2FAUGX5U6Rfy7uXN4R5ksvCMkprccjWSJLyJ7bqB5DlHp82S1quYNYkDwMhaINu1Otp0uZd
bttS+50Ncj7ZW8cl8zh3OyY5AJcQlba1UtIPDIjsEJhJtpbplnkwuGgZdZeDddsO1xz5WN6r7YsH
j3eYbJX8fOgsho9YBUZ/qIwT3wVWF+gWh4Dc78+48AOKK3lqNMBECUn6FLzdjSszARjkKA+HKuPu
fSBSOWtExkmwDZF2mRWsXywB3/cmmm+swKiVhrQI2mpWd0MJpe0hWFe2NvJDtrRKrGAeHcAkcDNf
n6FS0Pp7d8QImhaOsWwhATqTYtC7VNMO5fIWvxBUY5io2AGluRsIpkW+nOL5xpvY9Erpa++BXaVo
UHj7VU3Lc767q1RSM4cZZMrLVQaTRNM5D/QxTTb401e6mglXq9SBu5Hp8mGM2l1hHNkFqLOPFTi1
yOJy2bhKhkEo7uic+iCjzmW0LvQUOCXxA1OwBpRBTJmBNfCAeTmSvVpeRiiYhgYIREhUxz68XCKq
mD88+KQKdSfrM9wLSp7n+khvTc3xZCsyL/G+/Oz7qQnNYIT5d9NXtY5UZWSNeI4GKN0LrLFWYivN
QLI5FibTSVUTDhBneDILGfFjkGlQ0tVm9UywM9P2WD7OgO0uG6hMkKOV+pU23b+gdKYLkZn18wZv
L/VtxTrBNwvcgNR1UJ0fjqm9ygr0Y5rKerBzAQK0Zopno5e9Y/dUR9FUvjGPUr0xzbmyBivpBAjk
GhGWlgJJNITp+kOXXoSVop5nKz2taOqxvouJAyVReHGsyZL3ZYhpJhfb57Gki/27tbkQE1apWack
+PV5dBkSD5HT4WE6oLBrFpYNULJ4okd2SBUCay3alcbsuDb7/uYH4BwKuh8sIHg5bK1QdgYWo51u
AnPM8CO9rp078i4S1znE8KOvGRdwNGBKpt4IKFL0hkBvdkt0dUCY4W888HYtVW1W4UzGEDssUj3r
3uFsbpG4T6Kl8t9Qi7eMtGKoYhX49+ENk4iZ0n5UQQ0++iRCZykxHjd6dDjahVtfs0fQFjsmj8Q2
B/XLMGDSZGjWHA/+Ss67tUkN7XaVww8yw7TbUQkoq/fWGI0iA9xR/Bc1mK13+sPCyxLksTlv9XTH
nN9PU7PjR4YwaRFCM5/BtaGIJgC3zvQnZ0Eutq+v1lYds5nFnzrgqsQrnUV97xxPKGc8wdB7b1tr
4C5wL9FDrKSHkj7quHPb4a7strXm+9FkNzyCQuRiezi//JXEdhx9UaK7SrNlPx4jDmwB/XI02tRN
TdWWRgmJ2VSctYWGEaBHH5HIC5OsRexgCacKjyK/PJ5OirvXAzNu2YcuRrDu75r+6+YstT3Bss3u
DwwsS3lNPMa1DsINzTD9qUTpIZrtuQiGxd0Ii33299emnF1JK8jRGvbqIJzb0/PwFDc1LAGL+oQj
HhiPvyQr+ofJZnssIWy2Zu9cicdfxYQN2Khd8la6tPY0Yt6DdGASsatMyZ4YsdZHlUfUw4zspbgK
gjUGNKo0mGYlzVmzR8/CPx3hm76GBxhslzyoSF/pSrWIozq7zGcaWCJ7Ls7V9/2+JeibekEJzt1Q
acKMwc1egyZlDF/mCWNYWpLx9VWFT0ByuxjtO9jp34+S2y0l/+GYeYKtrfDVvT5JVd842X/cVbPQ
aSXxkpsc59cZWtqZo+fFQ4xzlYfqpFbF6xsyxBFOwkrcl8L9OWNT+89a7zMp4oZYhLylF2l1JalV
cwcy+B5yEJkBYFXZDKrvuPQqNlgj8Mgy+5ViSrLChiH3vMEgdPwNsdV3ehZ1Qn/04wyC89TbR4PR
NPuLina4CfkOJOE3QL7MjnT24APs7UL0ejyEgQLUCNm5gk3u/PYCk2ZTRsd2L9vCjOgr6F2FotAu
34gma8hnLzzD6ODaK6FKZk+CBNFRE65XEdhrPiKPlXQN9JjK/LxcPh8u36qFLDGquGi7bZ2DyMN5
j7dKZxCuRXJC2KocqhCt4kjCymxYAcV9yIZndLQS5SqB2iBhK+9MyjwscZ/ewgZhVH9J7vdHW+3P
LLpFV7KkRtQ4VyXxReYYBjsECbsArcD1/2vqkOnXXzol8j5sW5AAV4FS56BpdW/JchWtCt+w3Kxq
EfsvoJ6lsPBNkO5ME9wMGKxkWA2Xm/Sodx/Ko9X6ZXuZBcjib8e98vc8DEQuJXcDJ1mcAj3Nv42M
wS6Gay/xFgFVl3yJr9bWUmN+XAmr1KjsjqPJxaA5EOGN+GHSTnJiA3w/Sht0UidYLMD0cwrtja1d
fYlk6SMNgnfo5sUZtGvwSZE/P0X7g9A5J/LzRrNieh8dr4zjZfNrZs+vCiMwNyNmtD95SiorHQPM
ZZgGIT/jQkfXKEFvMtUnRT65AZzRXM6lGdo/qduCt5hGrIv9cRL/L/9cl/7IEhkCHiOFKJuiMJB6
xwVuqpnoPnNZS9XygmSMPPg9lYZruJ/fu/o4R3RVsUGZgZo+nYH0EjRo4vHMtvqJHDNoaWGsYqDu
sxl34t1e0OpVmyJp2OxGmrF+vsbWVEW2uD7qs7d/yvcR3IIfCl8WGXHR7J13hMpLWGINcrNmlAlu
FrWzuOOFZLLa9HXxqgpsAgh/IHitGmYGOWPFBb70rRGd/4gfosu/Tr5hqEjbvsjlkYwTeha22hpE
jcNP90+CMsgHSmYHsqZPzMsGEGg1hqvHJEMm/wxDoVqsTB43BhyiEXgap/rNk9fO4/Y0ounj9F2y
pihfsyisZ3V+NH1RUq9Ag7/6xLMvMLcjzEddlHS209OIg71i46/uG6ugnZjVldss8uAkd11aYTNa
KmANmCrRK2ycLiA1EPDXm4SDBjodR/G4YzPaya/HgLP/tAY98FrUVwmnbE3Sacx3LMfuD7rMJaPp
5FU8rpeFQb4sQ4Onif5GMeC6+EeUu4eJuf5qKgJn83nJfMA9Q4zCwd+kyRqdNxZpIHxlZZsppCPq
GKHYPHOoBCbIrINOabK9TU6lbvVyC9eodhwo/T0EKYTLPKsV8bdxSbf1PXo6dtVbapdlYWhkyhZC
U8mAfGsvP5jwchjlTUAMf64ocSfPrE5/oH6ZsR5rVcFTLTbVm9SsW5lGAK2PfpgmM9126veXlQwc
RtwmhgnyCmOwph5Y1s+ikjlTUBITIXgWTpWk3AJjgcP7YzoJJF/uV43Wke0GKhCW/yOvQHGglhAq
LSNIBAlTuS9t/+ndMlZ1abASLmniYUMZd5lWrsqTQhpXpryrX7sfK8r04fUDfJmuOvY/OHzobdbE
KdO3StrDCvKaaJRlUvN6yHZZDdeueKFFR3h/4jKpYpwm864jXzF/NdKA4EYxlKn1x++CxM8acUMx
HkICfXMbOn2547syUswFYXYS1yAFhjqMryS/gR3lgAfWcH8rq9UINJ4I1uqCQnbhcrJ7MugZ2eey
l18RhTY2jkI9/ycqFecNELS0yEL7r0Sv4TWdtjoOogQOqmo9JExhFUIERh/Sqfui9v4tamJhgWrt
/uqogpdAdn1RCLdZx+lB6HjLPFAb2/+s4at2zeN/RAS1LU23/6L4Z+9hmAZPihdGXhxKDO03+Jvo
ZI88NWNeGCi9wSONnvoE+rZeZ0o5GCJEsMie7CCSjvIvgxQCVcbWdl5yw9NtECRMhL6jejI3U0el
5bTUKCAjZQyXqPAWrV91mjEoc6j/oGoXSraeMSU2GVFjpZHANc9C0/fVWUZ/po7TDDRvflITgiwb
XMcYI0FLi3Gurp89FDom3KqMi1QoRl2fDqooATKeCGAxEe4Xg6rh70BZQLG+S+TnMI+tpfJnkJiF
D/PM3yHWm1pske92qlmYtYfL4OGI1eRZWuEDupGAUyEIFkuwyFTryTYUTIz3v6xfsEAYaCHB/ERR
ybPtPj+guEDj+A0A9etRKf0Fpq027XfMxOWl5DBXIFbTITBPRHR6n76lmrjo8WP+ySMTwds29y9f
fn8y/APYrys1gFO8HqD+wPClw1MV91d15PDyTgPRhcI3QLp9K9g3z0kqd0En93vrZzP6MUQrIoa5
upXBFDBwytuST1CYYD1KqlCX+ROuw215jNdbbab8fxeLRroAz1Kr0pWCkvu2u9Aeh1CFn+kOkBO9
IEvqfni0h8m/b8MhmK0k47uDwelmCfJkiHIEpjgaegusdoHxvB8dTm+k8oe0gAKWo6lewc14sxFw
9cy3MDh6h33V24gWHPUIo8qljrbH+iyFYWfDRau5u5Y/LDiQXHdV4DWid3co1p3s+b4sxryv2V6v
nlVRveT0eR1QZe1bw1jaKDsAvYhxOBZZs2R/ULkYe25OWgRkxtehv6GoeulHuk+9oVlrwIILBpnG
+/Uwye8+Z72VpFf9MQAXk+87N6+nfGbQq9bqdoFQDaJNpmzZzW6ltSy4lY6HbzHTVqrZhd/FdX2W
+yXi701R4KCCX1MJF7qopD8IcvU/6MHhZ1chK/ff4NkY/ohuUxBfDyHORVypMnWTOc51Kk+B1u3H
7Kf6EwFlP7OshrHf3u3oF7A5rJ3qyPv5hCrDS5GWpLxujQ0oopYf1deHPV/0fFIspgfn0RI0Y8cA
YuwbQ7CSWX6LZ5HArtrXu3VURyQOaKvwRX9wkko8/u7W5GotPmn4oGakQofXp3QYKoN5BzNPYikB
xrtb6lbUxR+d3fQpZ/uTK1ZOP/EyI3FsSPd1WFEufB8uLm8w6KnJ3ehhUspdV9zBa3ymBCmJhguu
bcKE+bNZHW1b8YYMHqptzP1U/P7X8K1K/NPTKNgzRstwIvHi4qv7/WkiFJ9aRkk+pMHa7FXLDajN
q6nGraI8+rsdun2mVN1XRy5eig3H7W+GZLtQNt1aMm4dxT/at1WkNvmEegf59RXwHkITYJxscrS+
ues5lCmy6ewCtazcodk1oE8E7B+fP3FgcpxDj9kJVJDeLVn89JJNZUHZN5YQ7xu9VXOvZkwbTxyZ
r9NYAYIM/UgK90AacKeVZ3jKtB25PidO0gM/So8LDj6ZsMpPRBv4NTJ7Ne8DFiCfOrRzaiF3OZmo
ZWXx5xrt4Ws+ipcTlg7ZK5KKSmZedIhpxmMVMJ1KqUUXX2C5m62/GI210hPnnhwEY74CgO55ReHq
maKCmO2TJZNOGYJUHsAampt0g7LDippI4SNA6umI7XLbL/8g0zcwP/tXd1aOZjaCQYl5jhi7+GOD
ep1bvtnMQM6ZhV0zuCXB1mkvtcutgHktPxMsFmcusRfkufqXUqTJuLqXC4cH4lxPvvXkIsWpZvT/
lVCxlkZKoRgyxoGrxy0hJKDd/2rMzhCmqbAsUIrDZTh13Vbkjj12EOxkYy+EKUhTSbZJ32lejot8
SkAxYTgKjD/VIpLilnY0lNcfUua5NpDrj5RxcQiQHiFwTF9EX897/1PPLUhkzY2IdzHOI9eKnwlT
xYq7Is8WRRQjiYCqjSTDDtPPBCAQ2cLyKxgLMicD6ipiy3p7kwSPuiXQobs84q14qxyyFm/+vXvJ
aOdQfnvu7MiJzDAQaf/3kpzNEBInT31Ovy3q3Db5adMsninAOY7/WUFH+VeqCGiFYnqAiHi2hrya
kP0kYlDMBh2/eGF/VzGpFEqrbbA/7TOSmgop2WblNfEVbqxJlkjfkWBVyrbRyP19WQRWD/7qZ+b7
Adp19GX11+w2Ltrsv9k6juNmVOo91hvpXdKUjBYDXgwp2egTeUOO+6iKuqtGVCa7J5nYd2Qu90Us
pNceA9AKJ5kQ8ujHO5iIsJIZjgS2dk1cFvxZt1GDGpPtPO+PHtXaf6L6YDYda9gByr/JXp5gvTWp
B3Oo04B3u228OuD7NqU93aPiqCpwK1tVbQYzvijQ4T6HqUA1SJUzJHEDr0uyhc+rJW93OEEMc2Fv
2J/qMcEPKKqvcb86TCD3B31A9swF8znd1yU4AIrXBS91AIsPVvCzDsF6Lwd73lKFgbMwCnJE8G5i
xz1OVa8IOTw/7XWH4ieuo31DcKC556I+jUGNc/JfN/qTuseF6cJkKRUAcb8DBkix+gvp8PSJsjOi
2eSfxEgixyd19WbfnoNmK3oUEPzzPTENKCJ5JKXNIrvU94exfM9UXHJV9XnmBH9wOD6o4fGQ9KKd
w8KVTkG+Q4+1wZp1yxiEEyXmUFkyFHk0OTzif7/TmzsuLDgqjG/H+6SZDE0IyVhTxC8qvWYhxEmg
GNKn7h/DE59PD7GqxgQhLKc7MZ5xbU0TIPo8JnCfsmiNEqSN/HgsCTYvWMhJzouHFCaLqCocistI
v9BcrWNs4gSsg6nSJIewhUrfTEtk3kAvuEBt3YgCKXZpS6i4W65XCR3kxzcprbgpG5HGMhCFkif0
rbpUBunMPp3RM2mAFsuF5ypi2ZAptnzzasY0369+TsMBedit9YoqKIn1OzDUPhJneO9tQez/9T3Q
WNXNtLqcOm5PiH1cqthc88w5zhw8ufOaM6+IRpfSy3T3MviJ61L3gQXv+AiRBBOhUgnMb8rpdUVd
+5cFlgo+3xppx7BnMIcj+OWu/j8AHk0HDUPq0nLDUodDDp0k2Qw2EdeVHo/gD7ZJDR8P2VSJODeK
nu9EnvElGEKuVuUk+fY0C6XdyplvqoBKbpyEqihxqorT0lKF+rEiZHOrlieyZ8yO8mN+GdtD/kod
MippMT6t0BCcr/JuozuXgaYSK3Mrs3rznnjBk6nkb/QZ6Poke89GgeeWQvF2RkM75xm5v0MDfNID
jeFLLSV/fvk=
`pragma protect end_protected
