`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17696)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5LHnVX2pn7aFXN7sisirCtQgw2EUqGnr4BEwd45PDpMHIFNy6gf7MF+O
oCVwCTFleW82LEUdayu2Nq7Ejf+kfnFzalK81vBHv/xeGZUw4T2uqrGcQxGzV9C8Hz2iuwXYaWvZ
pD5p6+Qa86zKWB9LCkI8LPb8/sQ555X5/uoF7bkknFrmjNgNiNTzU40jIpoZTCAUJluwS8SGo26w
EMi4d5ghNJFRfVjWKwkXWAL+x1qSuFe1UhUz7fTia77o3JJiidqUjgLsXEiwlbdkTZjlVrnNLhGb
jdSpeyMa9gs6xKHyEww73J2AiAJ1roXC8w2fGCvTtvYi+Y+O48PnedL2W1FhAgSRms3CFkrLV3JN
EZIy01fuIwx043cNhfX9lq4y6eJ0ALyfRV5IjgIYGTJJTqdDlPlmZcceAoXGz7VuDXTDleHBnAXX
1CrIeSb4BOoVgMbBIae9bjrzSx1hVV84WhFV0dXg/Z8DdhbEaPHJjaUM4MzzE8SdFYrZC06YJy6/
cp2yZ+eNyGKUlegB573K5j/rO6/dC3caZpVv56Y4eTOCeXW3KDmTEhqOZy6KHOptqL4vx5449DMl
K7J+8kIMtMJ/NLYzcRs94eui4XYyRd5jsZsVR4CQioEHlQZzjkA3m4gT/hHutYrSaVP41LQtLqoP
0VZC875pawEugoRHUZ1v9i1TKYltt4D/ySeBfspcdcIfbG/l4YsUT/WArhi6lITsa+FYnP1JidYl
MfNlrjTR0tFRjLYUk7bG0joa2WGHGd98EDpxranwD1rQwf9MAxbbnzRws48A/nuYH/EmNFJ3MNAu
bhsvcENg99o2ccQclJVkgSAonP8F8LfcY8b26h3BAjpfmrljlsw1TeGoABMGCtQpqkpNGWxq49w5
rB79860YvjojdvGh+zXWxv6lUucicfBGL1h1xxi6GyfpF1YbBXCSG0ja++UOpPp63v3UAL3hAeW+
aDm281aHZ7XYHdKJihahCSq2qcbXtRgXOl+ipCfHXZuU2I+7QQb2SONmwN40jhHsVMIofl8eFkrO
FIGIGhvixDLGpsQQDjD3QVyn5U1aol2JdtnS9qVE+jG5IPhy3EaDyhTNQ4KfYFHgxLag9tveUiTA
9bspaQVts9UbF5fMV22d8soVIBRrEpg//Kl62ixxMZBsVqjTEKdYyLAz3t3rbxUR7SV2HysIcUz4
40IRLbhtwP5PY8N3AKC0hKabpGcV7p7Yln8GcL4MfYwhLICfCVsUXEo3xwXPaVer+Alx7SUqiVIE
0yYazakdwfNyRCa8nzt7pHAEx/4IhNyo0zktm5djNnN34EeftC8Wica3dpidHPlVIKMXWEP3uDc2
1PsGtVU2FpYyzqgsEY8M3IiGmLjdnVfoyKYc6OW6HVNZcpr8VGJtvtvMlullteKxEwLRa2Kubg9T
RNJV++cIdAdySs1pkd7I4MABcvxzMRNnkXJpEEgBZHEAresifz9pkQkxvFrZ5XTZKMfFo4nWYwaI
1SaEeSGNiz03CFcZglVJgCU0fADuK8RaHfPx9/fS3ocux9Si8+qwZCeqziolcPqe3Hth+R6taQum
fDAf2yZ/lmz/ono8DJ0YS9e29bdWFKXUl7jZ/a8/EzF6Rai37e9a+yv/srNO+RbivjOhmaMY8c8W
zxT+eQArgjpUMlbTqQL24vFWura0IgdQD93H63QGhiNp8tsSyiCNGOpkefrCHziXveeURq92YmEi
xCz8efAeNhxwrgS1jtrBDogYZZSafUR9YQLUOkeYCjID9G/F6t3Mn2ASyUCANuzpvEyueUKumOYJ
i6y3LA3jZyCDuKTszVoFpU27qXWEgCpcLHfmfTEeveSBHGKW6Z76lN7dI0u+W1anNOgfEFXLpA8y
ASJ4LJ6seP1dKLy4Org+8/d1bWlVyeNg9S38U6kpxxDfLubw+4t7ZbO8FqEpEFxX/GMtAbeF60Lv
OdrNmA5UWxO1dUJSPuLXz/oQ3YP7KKtUPFVLnTpcXCGEFfqDjC9jN4T/LedE7arHly+QzFSd8grH
Cn7wP1v4bpYPQuD/Bnn2UPajxmEyC8D32VxxpMR4SDp0zWvi8Cp3AKQXckVjKxCg720CxUzs+mWa
qh036RjV9mtyKFEmvu822yatOynVbw7WTM+bt1fkrqF0pnzGPhCapERoF4HfySUskpVwy5fzDZpJ
3hXc+XPqNtrKxWNzReB2GORm7LVTBU+UuHgI1aHX5A9J1LWZUDEvNp4Mf7Mjnr67eH8PhU8pOyCP
z51eX29gsxkLuIWYHHxAp9ziFzaUXuY6UbjAY1phylDInq8fQJkUQoVME2PIaYOcxs09slKcob8g
YXNsViyI5RufossFAL0zZqW+H2L6Gu+Qpx/odYgUzmI1oqVJazhtxw46+tw5WS4WW856CF5t13ep
g2GwlxNVjlfu6Kbc3WAhieeoHLVZA/lLiqEKr270v82p8PGQ7HXg1JYilC8TIk6uRbkL21ewv+KW
MthbjjM6TtSTzW1Fs+SKMxuAz/egsKQVB6jgSrFncgIRB9uaW34Neu3zARb+yHVXVQ2CaW6oc4Ba
Up1nFIuv31n0Tb2Hb0Sh0l/Wpl8EK7PFvQLc2e9+lDWOem098I/kLgHoii0XpD/6KsKX0fxzMsAc
hx8O/Do64RXGRY44yx5TuH0T3Oaf8ZOSYjzkPT8Gmetfi6atIlVpw9en/zutIuaYaDrNDql8HRB3
lGb+XLvjsphi7yDmUS9N1IMGp9LXSdnJ+k4XMah7EBFwbvHcrQphcm2ViCdSYu4pIvEaQU/d3jni
bQjStNzS2K4yFtzaUKHER/jXx8/u5TjBKiY9CHG+V/Pc0grRp1SPHxxyJEOa0IP41sYTqK0Za6am
a9vi3zeeQ+mfQq0IFC2ry9f97x54dAf0DdgGrALon47j028z012VxsL6AivlYANRtQmFfNaeR3n8
CWkHydgw6tzlt8hVHg4z8cVc+nAPZtnGWVHxHQ4qjmLUk0YmAMaOpnkYmoX7AoeZVUMgLl7URjx2
Zt0ZE4wJyz8EAvQvvwp9mL/JbRyAYAxL+zl1/Wf9EVvBNL/WEPoYVIaSLY97HJJOrLQUdTs4qszb
P5IKXAaBDewUEhh+WM4uSMsRbmU4Cvo9OgU9yyA8s2r4NuDEVE3XNhUGCyRCKLnS4wsNZX+dUeUc
/V2xeWmbo9njCpwJy73UP9SSLhkWGofRR3V/x2bskkwDd3F3u+Tkg9m5Za1vWSDLqnjwEBSUGE6T
t4/BRZagEia/bBrTy5jivaCnwVYeSqBO2RLPg7/GjseleiVQf5eIlUx4x+8xuOVxmRyfEcSpaI5B
Ja5l5HPud2TN5lwmzgGONKFR4f36MJTEuyThpu4SV/RWjsGXHzZ/ekb82ai2A2a+nTcqg63ZRAGd
a8k8PKefNbLsGyyIXQYMYn6NAkKNcJwW5nQKvSAMIrLWfUm86QV6U4gtreIPMmdvnwx+R4UNNNgE
/2CxMUG3ezZZjZD0/2b1WqhRZMQwqpBaWQ5bGd/JCzGz2q6EKTU2tRNJQXu/an2xZ52cRzJ6HgzY
8g/LdmXJWTnieQ1/HUEI/XCxdLK5Uwe9EuLGbLqQAFk1ln8e6mxSO2L6KQTmIhOWgH60ZDh49m2J
RiiC+LO8/VBgjlsDYmP1J9lyT6xFvDE8V9c39s9Fh4eU/VzR8LYdS+tZSItLFQz8xSbpgOuFdzw3
ltCYagBoENB2XnSYk3eg46osxUu80X9dE+JAFUpkeN7oXDe0qOH4UvN2X8WlNDy9JXyDgpCxRiN+
DkYqRHQFzLmrn/qeWt4n/8raPPR+NJHaSUkEx/u1FXg2cqZy9DbIXZvg7T7QsXtEPcyuZfPMjg9r
OIDsur0NxuNDdZNT1J/sSUO2rDEWXhd05fo2wLkLyfJ/b7W3/r4amYdHxmu92gI83iw9YJYEC+rc
cJUKaIB3hoqDFry2B21kQ5Zzs3JRqKlwAP5zTixxbI3bbxf8pPlGtehJ9OhFFGvbGhq4wbkash10
sn8l6jNi6q7Y+dUFlPeXYWLPyfPtfv8Ix+0+GpPtCNEfOvz/vJpFH/FCPLD8hvamFkmBmo5gq4qZ
j5XHDR484E1gB/7TIee/pyciyjTGCijGnEJV8Uwjk81QvmUVAIoFwwIgdpwgeCkrUWxIKqU6kC0j
wNcXT+/TpaQs1K8SLwf/HrArR6E7VJd6MJobvFVH7aDVGpKwCoMpdmVhvjJ48SOSXcz5CRQ2s80q
S+01c3KAYyKvqSNKQS9Se22wCAWKAoZJVj85Sh6rf3Mfjv/QGikLuYpgUcmu89ZRtqtd5Z2820pc
UuAO1F+S9ClUV1TwuZyxS00/mOSdB83a1G1I7jfRA562axPkpF41X0ArYPqgTdsZtIc/WqIm2t4y
IPvxgRT78Az1qfRk54qeqveSzrybBXJMlP8gxMIpAU9MHewpGRCWySwM0smiiIx9yA8QQtSANFQE
XEHcMvFeP5kQFhPRHpv2a1i9vZwk+3yG8TGAaCUjUT5v+Oq4kZAxr450PldjgBt0FTMSFnK/4jHl
pXHBLZBs+nE9rl7mSNhK3ua+esz9YcvpUiyYnn9VASgUCL7aKZOUvehrGHK/XBoSoA6WtUfm7fcc
zit/FkWbE6ZcA8YJMpf74IsrQaO5ifNl2DAtvYrEHljz5o2/QVcbjYgGWmx2732Ijs2S5u4j+AIi
QvCWJlgu2FjVMcdnIJecdQbMFGUd75OTT6qyq26Wy5rLRyyneTtv9kbI77xVnelOS/VXMqvf5xUi
29/P6tNtGkl1amVHAscO6nVBOHOUWPjcm/OoyNcLZCTE2WMOVdmmiMFOCiJDUDLDDeTtON4/UfWQ
f/cFnLhKm6xKRf6KM+MWwPMc7ct8+158Chs1el48cW+Ve+HIYFgilRlZJbGlt4X4z4ySSc861OrE
wrE2zYiKSPFwmzYHulDewQXyCfaiJAKwQlgzFkZLamFdjDuiM4A8mdlketuzhWEkibrpzMDD6G95
K1hPHch6NiS2rYwFN9Bnlkv3+lJe3DJmmw5pAa6URDH6lQXnjgs7pigdjSJIc8NY2wlH+XIo8ZmW
3LTZsAbOWX5hVVg0IfQYTDcjGKEr0PyMoxTp10AkIeP47c/mIXlHmkKQLrJcekJVCdvlvRSkjX4M
XWOi29KK0hGoEKk7MZujXxE/w9JUZb5StwMOpoNpzyPoXieDInwwT3b//l6s/uXHhSEu7DZAaBmE
XokfvNBjTkXSCMHX5n98qvrYMMgZ1l9Rvt5/Whgv3K9zXGYGRBArWZTxc3z3EWIyvAeHcoxvzU6T
L/9a40urIXombdMuxvAFpqPY00MkemfXgxMDqk4eMPBlBUqZhMGwZILCTFz3w8Fw/S/Dyu/vTeJk
GXzRvkJrEMPsIt5vAbO3iQdT6GoXeNspnIbJIAxVSuTFKkHRUgMRxneylUqsQ+3dLlkbJfyu3rSH
YkLaIhIl+9/9ppf2kSPUrGu4Wc4rarIiMRKkMFWEBg7GgpurEUz77NBvMZHaDWcDO2F6nWn2AGOh
y+4UHBUKpMrwV9xef4I4KPzzBNfGG8v3U4L6SGOX76uqtIL+9Z7TgdhO8SEyWXJBUVD2fVlJ+r2T
qooTfssztEzEchaFMDnoYgatpwsEXKcaLjtcJzgfs7oJEPmPDke7Ni3uURvMORYLrmStQiel86iT
a30BrT+sWYFBYz08iO9icfbIeZ9rqZuROD4bSAsr4u04yZ+o2Q6iV9amyutjAcLwt+Y6TM53UH5Q
vYX3d/Mq6KRAv0khz1i8VP8aPgWLbHwYdxURImwq+gZn/DSoj4N94+1ZpdfR7dVgVKZ2js7T5+Gc
/r9m5Kzcuv92fk7DVz2z4W1z+Inf2K0ndnj0Eid0ktatkhKe94sxx1aVw4v5Kn4s5FCOouD0KQp1
j14bN0X1xsRMLJFBRxoQ/1rzNF43l6s4430IR0B5IKKTHSvV6iO+cZChiwhyFnQ7neujRlilXr5L
oi88hEM2alS8WA9hX0InPJYCITwDuSSvBasGPCk1fHSnj4BiG/449zwGvBxi6B/12TnjHwmBcR7C
qNL2fZ35+pr9UjivFwuvare15/PaHa1PWC7DFlhR548KbUBZKbH58BRqyiBaMo0xY4FGT4KW81g0
finSzSzt7MbjGh7t1beVYlb2afAbGTWLjGa63M3tiQoQ5T8EM9rAbl2hD95FqUfvpVEro1qq1TSu
hdqaO/4HdNERK/ERotaz0iRS4KVaS3tHRCXxlNtlqX4LO7bz9ItwK2DHEyHJ4HpLoNd6/8U73h/f
5e34VlE2pFDQVQNPVT/JJmMCalA9nNq7o6ylq3sYAvlPYIjGkBaySn6hqKKlK1+CRti2OXol0XDZ
HKm8KM30i53DPwWGVeiMyY+bAAOEfi+ukkXk1pQh9dKQhueXpjq8JpbEbBXIL1leFCbgemIZ7GTA
khZlXE3pquLcV0O2O1GL64wE/y6EM8bPdIqrYWAvPIc3xFs3ZRt03L4MVkUx6otW2SKDg3XFbnc5
t6tlBDu1FFvkzVpFJLimLe3qnvuT5ZCJak+kvAYAYYOqWIZApyXWjUMFPLH65C+5vWGurGbrsI/a
FrCUYvpH5i63Vv9dDEid6OfhGxgqvyucVCyA28BEWAHsivyltcALAD/GZuvaSQNjzIQljscaIBdg
uxd63h9RsujfqvHV58p3BviKJ7oT9WyA8slbU8ukxP3XmKglR8apeTqg6S4p3GFIZJnjd+ztno74
tXH8Idtg1BdUdiVLSDLeOvlsLCyZ1ckIRCIfWiQ/FXIbkzwp8d4jvLNLiqGxXhZ3pAwI7MAnjIbk
vNde2x2NLre8OS9e0k90GRDWMrbrEA61spM72jbE/MIS7lM46OWVsnRcYH8FSB3bfe2Q2AfFyYvh
gx92mVQjWCouKg61Vyf8yxCzqcj5C7RnEZLwHNLMloBYocM8yEJC3hvJEq/sVASuZRWi8QdM4uxT
XS6jtXMGk0m0dMC/1RSU9WAzLDMjY+uVeaGPhVfsDta/E+kjNsDTfIKpL4qHc9p93SAEvVtY3hft
KrxyyMT4aMEhUbXte+oHH2AIikJhU57LRImf50G12ej4FtmkOvnNQjTQp5RLav5vZuI4gR0laek2
oBpAIgkolDZYFCiYs6MzXjlpdrPGj5KnB9n+eHG50UbxQKcFPDSnNHc5Eu6PHOAUT1l8WoDE+9cy
vlKTe8uf1GvmDPOg/WxGtmprwdW7Iba/2K0jTXRHo5W3tN38xeGX2uvfx8QxvP5FkulCLtU6deBB
Exg/E8Ktwret7S4sLnSXr5WsEMsFzA8pl4BsFP0JWFmdY2GDGG1uifThMh3u7iZXBGG2KMtaYQN1
VVD6Kh57fVNjL0LT51fv8XWj7g3teafLTG0kwVBomBqdvmKBvhkWACfdMqqjJfZqlGlrDXTrvUEb
Y8mk7QtMBl4lm2Al/RO8PT+8yR59pEtw1/H3C6GUiSv53pLQYxvF1E/Qcj9OajWmthP/8yyy4Ov8
521kqOP6c1+cYEVIOc4qFnxt4yM8P0/rabXk2Wwg27XcoTp2qJh6ZoqTwMJC4HHuHnj6rB+MaFA1
G9qXLfPvE2UwefZighZh0mkbQdWQgpJczqconUvfOSkleA9vDx/qhQda2k7Pt0U8hpNLWaUqsvqJ
jvoxBCRPbhWNCmpquXuJPtY+YqrElbGnP03BsNWk0FVXyQOYFtlgh6vw//AUS/Q0ZvluVStkDzke
nx5Jzs9yI50MZ2pddzOIgDbbnYaeuRB67xkJxwYXN1WGnujkMmvkJ36JQ2IlKZAyZm2A2abpVC4e
UHZkqPuWCTcZSE+XRWvoQdrtSnEw3F/L0Gs5kJ44FYOZMktd8Gljhu9Q7cGCnY/Un81OcDitb+Gr
WuzCl6d28dPU+Q1zaHS+mTLP3Y8WHGEniowpjAuNWWEO+/SXr+5IrIgTGN9si0HbosbghYvfl4iu
Eq7APl79+efqDWXkiegfn4aYpjyfjQ2Ztp0/dDeli2PG7S0BDSEsD1uhE7bws1safxonX07PELaQ
uWNru12AIAEUUw0NAvgRLhM2wRWM3FwWfYus0JnkqiCvW4sqcBS72F1TTU9QD3Q4fz1DUUvOfqnF
TScLTV/Zdgiaf02L9CSeGfwR9iwDuqVWCXuF+oPJ2o9e58QiKHCpRGCSByGbphrI3x4pQc8LTMkF
4EnLRyOH58vQ22chTc25ya6VxPspuAzpm6/22UQvQONxsa4BofmqJzMuQ6HqpHqjUk9YBuXpOcjt
3yBJyqlvDQ4HyPIKjgQdwQjdWKakF8+LT+XTN+NLKcSCeBuBbo+dmC5haFU+dNRIHIRGlBLqNNyS
SIvyDZ2RJULMqb2y57u1139AKSWSqsNH9fQF6x+T62LDzxINU7P91AOdBoVLsHe4VHAF7UeVClmO
SWytnAxYF+GTXqhrH4ui59lxf2gtI84pF/P2QOQrlH80ZiEQNQ6IM6fI7ro6WdeVEYaMIM/CDEvm
JzL439psO6+2Q4x1u1xk52Zu3T3GXDlNAbMM7KIAbwTQNlYYNCp2B87v23ACVP6RNIgUrvZgQPK/
NJOibakn9mwidvkJ0xE4CK2hMb4XMKURraQxYxGGdWHSiLf7kL1uAs3CwlBuGdY7Ogr7mO3haFyl
Xu5yyv8QoT2JcPlKtIwYA7II0FaMuf5aIWnI3l8Gd0YWZ/5MKEJBuAk5fK8PHHoROPb8z3ayAzqC
u+j2hoyGnE7jOrSD5yLCa/2uDroS+aGbwQ3EpW4oeziR3HDCSZvV49BIaE7ZAVgv94Y5fD75FdPt
EFse6YJmkKRXdPlsrxM/LDXXaAodgBQyNH8RVEOEUsnojdHEsPiK8JaLVHzzGeo+/uQj8PdI6LFG
Yyh/YapwTJ98fzqUn/qUaQm+8nYddw43rQNudbAr5JTv2ReYmmN9MXGkBFy+HpqoVSNRxObqm/5a
yPG4yJmwaYAyOxbYAhtK1DunefIR2UGMTCm/2fk/dUPP4K2NWBVhTC1wliP+bbvKmzHWdM/SbXXk
fhgJp1s8Yj3ezCAGYcN+q6lUwNzo7UAaJ3lrl9+W85GF2+dA/A6XKicFljU5WZJO5XzNogYf8NXH
sRU+ZXEO76Ry9JL+bgiArdAn0ZoN6zX96ocjTsB+Gny1A4pnuAZzOTzRPK+N+SlSv687FpfNZQK0
lcclVzqTF3wrsq93ipCj82e1kzSx3XCgVGXqsMCcoFqvNAdeQ+Qxhfja7cPAWiNacNtk0XwkzBnw
sB8YO2gvlrFCD+XJMYR2PptS379IEv5/74U3qk85IMjUdtR4uA23EgQKZFyTv5ixMxCet3891wUk
UaJgHkeQ3pvJg8+bOZOs2wOMtC89X3ezSwUnj97MyBAOHNGTOaSaP3fLPlxN2O6/7R12LPQvq1Ov
taZMyJuPKX0umwo04q1msBJzD//UX+CwpZd6VIEVwbTx0UscxHpEe76cjdG0bh/F1pzLgQxM5dG7
V6oPYEWOnNpujVU3M83dbD2A7Y20bfGfeDEbKEjKPq++mHphbHH4Euws2l2p2sKOv0WN5CSqczl5
c/MVH4HCYaLhKfIfKy7U2tkghXgmF/y6HL59JQkx6JfavDl26PVk8zjUYsz+XDshu+TmltC3LD3E
PKz99vXzIg3NANdHx6lvDhGcLAeQ91k5rgT3zRTzZ6iivylM58tVeWoyE4tvSy/nl2U32LSrYSWk
eV2z1npfX3Pq6mwqis4+N5Dg8A8iOzVKbIzk7Fz4jawrB9SDgdBWx4xC15COnF/yObWVZ8K3ZZ5O
yNrQQvqmPwwAeneTgDjXZ+bIy5tltILu8kZaWk2rJ1fbHhJvlF79SxV3LLK5R00XdyjJaUm7RwET
CIkEzpGjOYCPjbFkkHEEvBIFsVrLCv+j1eRNBvEL/tukBcD380AW0kyprfMMCohhmiAU+cU0LyB2
YLBnHornR93B/pTEBSSJAoBKFceOKBE/vQzaUagmRR+J/hxadO21vj1ZXHKTgm4DO6yQ76nue5Nn
+Iz8kkDpvShdfgwSLP+KCCYEkwVoa3jAznztSN+kTJ7JWkq6bcIk4/PzuQrKbUJjvyv9Nf7Jftw8
KBOeqZJ3W7nDb5dAt5+nAVGU9Rodk4YISB7CQW9J921J/1vWrj5icH9C/vWgGXd8mm+GhRuee61/
ctxpwmXAShrlou1NVV12aWpnyFeJVLmuMqthgA5d1PNuzlkcLvOY3Hc9KfR0xnXa+7M8ysKv7As9
ErmY5LFwHAbucJ/5hLpdlaVTbM32kxQtLGRpbnu+/PLaXnntyfKIevShB7o9MAsgeHFK0CyBubGt
eZo3SPLBxj2M7nTEsjhEgaAJ2zx5xiM8R1z14AKGR++B/voaEZvHPyDg8s7IT2yax+hjiqidcqD+
aRqXDY6gK1P2N8QTdbYCz8ItV4TNDV2ZX6rBGxd7eWhhO8Gz6fnlvlFvidVnw0OOJASCbNEfKNRN
D7H39YuBRG9TJv3Zy7pXMHdlvyn4IjCVxSOxh2n0XPkGZl9wNTbOiTE917nybhI1lymlcCn2wKg7
hWRiwO/U2zoVb3gqTay6S8iLsH4Gv32+lMC36UL0908rAr2qlGiAr7QEfJ8/6uR54V2QAxjEfe/1
Nx0/r3TPuYaKOcpAGLowJeOjRwTZdYZ+y+xrrYCVGRAc9mTwI93WdCRfrz1xazcaCqLechLHebj9
tJXc5cN1JlFrSx+FlU2i5J5EKi/CjubuTV7ZsW2mqAr23j0JPx6UUUinphBSGOxPTPuvKv9Vem90
NWSWAWJ/PnESNqK1tuLx9K4i3OfG8Mfntg00I8bazY95oN15tlIjdOtDkb6VSNjW/GkdsECUSf6I
tybOpzdSG3++9TMqImKAFet0ZItYOWceyY9pEqNUCpXZQ1BZohR56ZY/nDX78ucWn551zCTjRt+v
1a1YFL4Afg0LV2kY5mmlxi479/p+/EXy9cRomVFNn4RLa3gevOFDqOazlcK2EJPPFra1FgF6SXf7
zDMRhcR1iiNCnIz0Bl919LhFPsLSVSiy0XKxHCbpypgzf/1ApQcFXUqTW1a/N0zN57gRqRP0eKIE
SosLXRMN8ouVYLMWDJbSUrD9q1z+cgrbPcNcN4VJZgpsrUfF6w7lzMmxraZxMmZysMro5/Bo0ta3
7QVhnqkGZnNYmUbTowr2Iuec8G4VoLVkvM7FmFhdwB8uOFtuoDVaKwwcZz68y4Vpwugi+2K3Tzpu
T5X58doWDtW8f5S95Eb188u8wJvpYkKZ5G2VSvVSd+CCzRTcwi2+eTNNkCnGufVD2vfXJSCqViZE
IKYZWtubptBNQklOaSS5adG9qw4KtwGsFN59znWdHmILFkvlQ/tXTgJc61fRYFY1HL8WH9N1I0eX
PNKfksY9qf3WM0hV5/OnYWvrXtsLLVXrmC1Spdj1yGu0sBsuOUJBu9JV4pYeyhajx7VcBCC0wemP
2Tm2id9t2iYCL88JyYDtjaSH5wIcqGQXm3I5OVAtUzRCTEWDAXm3ad4E+Mfpg1dmhAUnYaMTYSpH
xvUH2SvkYOq2hUdIG0pLvBRdIKIaHZhGjBqBHtlUjf78EX24/ZdKFLzIA+BcnUpn5lMdymz8HCWu
BqpJ3gu8gKsaFU5F8KOxdX/C6Zxf6WiVB8QMrbZUZD4O78H4rXO4bYRREDiP0NhlEYnxwBnPxsPI
tMv2V57KIAQjNxgQoxiT0Vonf2jtlG77bFaIVA9dZsT50F85AlMmfu+Bk7mpleI5VGzxucT+Numf
1BjIvv4/jqMX9+IazLmqdbjjWT6WMFStSq0xRTZBYSX0DulYf2LUU1mZjVwanREpMYqDZutmI1Pe
YCB8TV9V6JXQXsMm9ygEfX3yxQmiS14XPzAnbOmW7XjXPK1YKwJuZOYuKv4dacS4QsFS1XoUEkb4
genAJK4OsKXBHJOu7gSfOtBVRy+dgYQSZOLlQWJiVGD7WAPxCr3D00pHi96T2q0bRFQiA/bLu0Iz
HqU2Ah2ZWcdvd8sRQlfbVBEOTJDtiyTNssY2T6hxC2Bo3cahwx41IIJx6xNocbKYxG5vWAbMKei9
XMhUAi/Cw7vUEX+jxjcbzW+rp4rDXfh1kyBgpV3RrWLzHA/oKPNn6LNtW0/qrXBzCSH4jo9TtEPW
iVGejWKDiQp6xlJdfkRiyhQAkugE1S040jpLyc2f1S1cgI+KTwMtwUsD7uFuW1iylgooZPMYSIpN
hr+I0iX/ufoKYps4Z8HFKQckMh5qMDSWrzxnsto46pidVy4VmySLEHUaoFzgZRDqKC4h3XMm11pr
crLop9MIM0ZDshlQP7fLq8Utq07GGV0wQpVqi5gS84QKXar6RP9T2ppxOYIQgpF71eG0i2O9JOm7
Ge4ea92NJuA7WM1CTBYcfs6vTQH253egIGUl1a+TAMJl4tInrDUwCUZEt0welAjZ8o9b48LA5P+Y
urQhmTlYKNjjZ9M/QAlU7D8dSN3R+kfKgYDzh6IJ1FpeQXdowQCdPP7Ua1kpeQvxSqTHQN6oT1zO
ahG4RvDtyPYlTRosVUbSSTHdg5iVMLluDaPVnSkGYTSHiRpKbydRsZPrXZx39DXINs5J/q69rr4p
sdXqt9PO4yrHkvRSK+1A8IIh91s+IQXfPyEJPkKCYaFc+KZ5C5uJuS7vG7V6L6Z+EY+HkXs+F2Rs
kClOvOcl175DkZakNEdW+bsfNXduzLrPUNeeK035/H6VSJZDuRhBJJtQJ997MDo7ycFPKm7F46Ud
nLJdzQyyPEscG6MDGmiTVIeYrkDLK6FdItPBLcWPVFDHkwXRDi5nOQFn2b/rtJQx/HXY6He5cz/l
HXWD+99x3OWYfOHx71yS2xuUTTMCWNnrHCP6o5bJ1qZn2S2Mav/yZKWcbnW4Nzvz77gjCMXh0RZO
U0xlEj2gfUYWowM/h8QHvoBq2KTcHeFxLOGbi/ljgW4mP30G+YlCN+/GR/n7e5giwZAy4n202329
Fr8LThLGFRtZ+TEmBAAyOzWZZ/Cj9qU+c7SgeWGOZA3nqpFpqeXsXw/YOzUxYoYax5gUFwtALOCW
ZrjshlV6WJGvItAZJH+Kx9mUY2EU0uGUWPiJtfXK/0HKvBxkgDOKDCQL9ZV+8bplxSUKWesMXd/G
6B/gMCAsm0FqxXr2BGpgXEA/9ZivGETTSP9ybPuMA80ukhU9Kp5LGsvv4yaPJBOeeCJZ3sSgL0xa
2O6rj7GIPCrXVwB2X+651Aa9LrovAcYYl5/DuulQwR1tDwE1LjXrC99TkJVGBYQv5Z14UHWG6OpA
eY+brAWM1mv15zqzEtMqfkBrGZJH2Pm42H6SSSBhfx5mVxzW1SKTSm1W//1hvmwxl7tIgSVYCbeo
j2dagyt3YOOI9XavamDvrsUdrRvLuUDH7IjT6O4TNR5dI39LebjeRglbFHjlzltC9QCTUfAnSqdV
kZAjUIS+/6ttOpow/BhSozufcAWyCXfRUyDBSnnFmhiHg4ntdXP94siAhO/3Eumw90za4NH2FpMY
f245xpZ26qT7RIeUnap005XO96Wzk5CVt6oE/m2CwgWKoa8cu/3RrhOu1lQ5NA2QcgGr6fJwZ7RL
ju7GlHcIGWEpHULRZOpBgSwhH29IPyyM/ivkCl4pPVGpUX4h0avFkVlckltQvQJvkU1In4NK0BJv
XXtCUYXbhVZDQ4fCquhdDhCBdFIBDUH5fiY+y2Q/FhcTKDrP6CDjdLcXvYJdHXssoru2YHSyUsik
tZ10tR4EFxQoFe01ZChif3i/vPtUjuMR7V7/q2GO/nYr/LnpobAU3TPuB3jy8HgzR+oXnj5dGPI3
JpylHby6KVwzP/g2Gdyp0Nb8zyjxDmIb42Yh8I9KU+sA7NHPR7MpXT+2XZgEeqzW57r0Dl+cr4Sn
86wtdHxxfAaVgb7nTOibTYAb40l2CinTM0nfSJq2c5tiDCndUymDI48LBm3cqhShwa6DePSsm3i9
VIANn4Hh5cVMnm8q3cyxOHex6RhCNN3g18Il2YsoPc5kGI7arNU/fPhc+4/vJa4Jqd/ayUwRSQhK
FskoDYRr13NnFDSHNNxg3G71cxhvTAoQJa1cl+T1Khc0cs6N+ZY1m2nCvvPKPTDCbO9YPjcOIgiH
PpNdHI5MaNhm+Pgjf9/YEOumpO6+hcyrhkM16EKro9p/dv/eCvb26RLiIISsUGkQG9Vi4oBXB1kx
uHBY1z8TTGT2aVIu+dryz5fqkmFWyEYzq680ju25Xg3FXMe5/qAL4AB7SsiLvC/59pXpVdfZE42j
Z96Nu8xexOlx2UkOw/7VYGGajojFxbUZwQP7fnUpA9hqcN5L76Ve5PfzaluJOkhqAaR+WrBmly0h
KhZdUBba4TSLzMzLL570pfxBd6U8gGP9OL3AAY37bKExkH+pzu5gXM+Z5qeZ45AQObQlethNEOPM
RfOf1882WXD1tjOnDxPUpK/18g3Qlnmv6jyXG8jQ2QjvMJjpKFtKl6LZkPh6LMjGjop/kJgZlT5O
DqispF87+AqjrSartsSh/72vAz6t4a5CBx+858hVh8rQtjpskFbs4dg5T3VTJ5srEXACk4G0p5mM
c1U/+TlpYfRS1Cv9Bzu5RjOKcDFfdz0IVLlfXLsQxNKzTe22CzLa0uIUB1Nky8bO8CxfzGGB2xbw
B32bNN0R1+k4R7/YQTRV2XaW5logvzAfqPRy9ti6DiSFgYKSGBmBU/5NPKA9iWFxnn511K+snk4V
7ixGI+x6tQOxqrQV34mknNXCRtJMysKY0Cxg5Kzgbemh5Fz5fkPEjWv5saVEY3qETYaAwQNiEsNb
5AYGIj5a8PqNGPUrk1nxM83d2QYZvCARrUVmj9IZjcZzP1tM5e1vGh0L+g8y9YgVr5AxnhScavqG
/Y9cKxEYWMonm+9uC5At4xTXJm9ziAOCNGD6cjTGJFtkvxAFWIlKKgGh26Www3DwAQUYAoAp83Pq
LmMPMZ+8ejkc3/3+ALGSYLIBECNikkqiMjWwXdv+QZi+QwmEKSbb1NcjpIYYWX4I5ugqzwfQ534z
qg9My1lhCxriXVbmLVGd6+VoapfXuzLroMCTAtIJzHH1us8GMnOP+kjx8vQ4d0MIy3/os9LBI6iz
twWMmnTWxL4tST3U4AEimhmjuGX9/NDJ+LITlBD50emK6oUao5eTxEWXixcr5mBlemu+BQJR4sZa
9oP+RzqkFiTe3k0IJCsMjKGC0vcro9VsJraHYJojpJBe4hlnSZYGFlnbVFpofPMwolyRdg65u5em
WiTIsaCo6gDPZVBTeHcM2PbWe9vV6ZU7A64VTvb7DpwVN6a4wGf3mQhAOXSJB4v4kVF7il503qkd
Jb37TANPBaWVtIXFvnJ6l6MVzFTvnXxLxvSN0mwVp6yS9DK0VqbOJ27otYOsi/aUfztTHPquv8wV
Uz5f5aKglkb9Hn0heMXaYm5/YK1x3glF0GDvnvhPNJRVYlsNCmfh6qix/XZHDrF8M2+KQ9+Fnr2Z
5oLPTT5lXtzFgihOmPTw/hFAYC11V74KUTHtZcEQl0LmZXlWcd44kELzl7S65AAKwLxO41/idbzy
Dzk4JVnAiNr9pc2OwzSr2IROCoir1gzXDxq6vtJKgOhfLTwVsTunDigRwUE3f//2UmuYQGGF+PyW
P3Gy2mLQiA2WtGftsHPDkHQoboedxPps6UuR9YWEuAYk+/U4HQz0Pe64VCKXH8hL7DXCXbwojd1E
mCIaqy0TNPcsRhcF1n/XoVyXGxSiv6kc1kfcib+OBSXi05aPmjsLDQzJRTxIiIQteY0S5MIha8qO
Rai7BJa0P0USWNE8EmfuUfMt1isucJUEM3DnC1Z4QO3EYbwL841sIW7FuU+RTL4BKgC0jfzQZNwz
Sv4x0uJSIU8a+MYUujy/8+B3TqXa4iS9LtLwx9Cz8PUS3TowRe53feJ8KB78R3hkMwW3wnwMXuJt
H76wOHyvOV1S/X/RhsZEh6z/TxiT+eGJOelBYV5ZUAy68IPIfvLyFN0Oii2dMGQqFB84EfxHAQik
K5JR/dpiewKuV3Lj+IHh41+pQArn3ewqOI2u+huvrCDfOE8Z3mS3jzSqWqUun15t/kkmz2c/Komn
O5SPlOfmEzYv6uWQkWuW2CF028gEgt9DuWwWFXU8WpGULjRRU1XRDbrEKP32A02K18IlTWi6AT2X
qJfUyed/DZGe7N9cd86Qroe55jqbpdA7abNG5w7cFLzUi0Etr2DpPeohEfEXVcdH0DyGCnI4qsz7
AlR862XAzXTcTVZXR9Hegz7Js+C0CvM7MwG/PWGfUOl8xJAdL72LoL58ccez50TTtkPTPA4Pvmie
bxxpL/4AS3zvV9iv1odQ+2ua3JcVcOjgDIGSB8flG/zkgXIfwY+lPPXr1wHAVXQ+5yKl/dPmZD6H
5cgtEIq8bwDIYk0xWk+MjonSgfPjYtF1fW/nEY3YQ7Ht5Qqh6a+CGu8HC4pNW5RmaGjZyN6jxI8+
rSxm2Y0krLpeHsAY4gdTFlhU/m6sxGVR/Wo/CP6jZYtSjTTZzuiVng+8Xuyz31MYX05O5D/1TsTM
Q0IfqOUINCesESlrCVdym3XFI9y7OHuBO6W6OufdjpqI2OJsAp2MPjiygZTAlAJ792UTNlY1a6bV
Ml7b8fb2tC8xDWKblenrb7o7vng9vDH4zuAcTBr3e2KQhyMw6YvS9780mzvXPjRzijwbJJFuGo2M
vcMox9lZR7fqsrTYuK7I5+NWJfHLX37696rN7tGIizTByo6UHAM5YXSdJeqY6nplidAwV0mIn7aO
B2ZnEjngdpwlkT7Qu9KDV3mCoNrnGaKpA+XJwp+pi39fE6Z3yobkNUfg0aD+D4urDfezmd6uAjLm
xyq7olojrADH1Oz91cWeR+z7k7DJAZaN8Tu+Q6B/AKkqiiAPFT/TKx2uKDMfDD1dHq+BwvjF7dS/
HOxXd0ShQI7nS8PE1wh22lh3NxKRy01YXpd2IPzDYUDn00Jn25mba1nAwsRXS45E7awx7r5ro6XR
UM+ho+GZ+gzNO3+Ht5cLJ7A5UZXaZHNAQ1Ky0twvHtiV7o9hQ/tTIYC4fKZ6J/Bk1B28bN+zF0DE
nuTM8CisXKSqqDs/E3gMCApF6TNseTDm0YgY7f4UtNzxLzw9ZajBA9Xfct/KHaj37Eke99xep4mu
nZqfyT7gVHAjgkYnPhMM5CI8XNzJEJOWFAy9G/Uu4GvtbrZax3Hi1uIYfd0HsEWdjpXmIZ5q6C+s
fliJRxf5qocSydy/V+AGWbJMfoswaAxiyQcdgZNcizvSyaeG7oNyvNsAqm6RQc6omn63OKmmz3Cw
fsszI53AgSk3a9CymteM6ABg6OSB3GYU1Yv1fniw8LWnNMAJwx66rXgcCwC3mOGEWN10cqodyQlq
6szdfn+u2zbHdHcc5CsshR45bp0sCWb08SWfqQ73KfRNoHiEulU9LOpTPigj3NQ7S+EpVPgll1Ls
34NokD1zhtwcX40l/VavJT3cEqPj1uqfFToscOLfJeHCvuV+UMxYEzTgDp9EcZZ1/Q3sNNsVgjxs
bNjV7U1C0iL40yROP3x7wktKowOvBpRYa+X/FabuSJke/pVgZoiR/yBzBiGEm1+XSWv2xi0eIVl2
V1mGnnUinr1xjSuZd9Kz4b/pSsSIFIk8BDSbD4FEOoMUZvTI0zXmCefdxiWGwn4IlFfC8thf3F91
ppjkYyplTfsCWF7KIzMgXFxKeKzZjqKv/MTphJqtuvdd+KbdNqqVVFhp8Q4VkKaPJ2k+JtIoWcCu
zeLzON7vXErM5P9U4pnHh5nofD+bFa8ETOc982QFHqh20bYci+mdHhFIleypxyfNkCVVB+1Dh056
z7PU2fjMkuYufkl9XzLKKiAfu8EIgQYgE1XgtBBs6IR741GEjlP9/NDRSJJDMZU6UxuVKrMUAI4c
mCAtlfvVZuQ3dx9yyixVvXviDM/JaOxSLCXeabpvrEKCfZjKYV8vemKMOZVRvSbDf/gv1VRkgU55
Av3knp5EbjTAnyZwGaUjdnj/XB+dDRoaVFiqTYGv86c7KRgQdQvnRehohb1GchAhCQjQHGWVZefO
S+hZ1DXup9Au6N+WNEKGbpNgt9FeZYW3WAEQ7RoFKvqh9wcsvYHqLhfnOC5KQFf+nVvffzbbFGcT
nKMdcv5BfxWlY9hwuxsvMnhUnXTNbfpArb5pGb1Q+R+OOhVMTvdUenVoZdAinaMFt8OAsvi30fea
hprPoUEUzscX1aZ6jCacHjUkTFpvLeZ09AkNzjpHnsMDJAJZ3m18esrKIm5Er7/Amd1irVigxrso
NQq9WU0TH1MjGXaqLj+sJMCBEIslNKufd6PnhgFNrg58TIG8khMxeqhNtQ8tAXMH/dGn2e9Js4RM
mnZROkizKS2ZxsYnfX+UAy9MOsjaXsDXmCswAnfA6Yckz3ZiT5eGMGhXvuzGgo9N6g5vNqfvm6He
8zCbT+BywZRXDtYwcRE1sKrcKxTOQmET+FSE8MECUtX3MUUW25Rsv7625lDV4sguQv62oaLRv3IV
lXzWeG6ipMcWkemfdNilfkeAeB5syg0hEFFPfF4G6zRm4OhATQiLf8FEW9HgSE6HgxquGhnFmFcm
FCZ2PviXoqTE0YuBb5/bRVOG0L3lUvb8yvARK10bVYjATJ7GSkXGLHpavGQT286JTN2Yh2soGMc8
hVafQbp2SvKmvrmZOQoTpuSlbxjk4HGoNp8/TIHURDE8u3pA/poVYE8AeDqqVi5UkRyR5Fvy3t0H
0kKFtLc/AhSnJILy8g4JmzunuU00KtQG28DS4BddDelrZ7yBy169iO/tNK5N5MWNC3APLXsBypNn
58XMP5NLpeyjfYSouXnQHKhSEkfUhI9aCRrAZUDLMql8gEwU4RtyjpKG1YEMq+3DepZy6giSus+I
eNatEB45gmTNXkhMxUyVkzx9GPUe8n7uQgLtxlmSgndn0kvs+LddJiIb74C9NcHkB9xInn00JgmL
9BigatvEzcvrIf+G9VkT4h6oEr3wDYaba6StH6GHMmucsAVdtuGNnml/sztjUTnE93jwWF1iVouK
BtCO9dsYeBtgqN+Xy1PmePtSKR+RZiLTgCgDlqehYO5laYIft+DEF2PlE0NRDNVQXgykQdNt9Aft
O+eDdzwL7O+LPJRg/XuWqlcqmvq5Qgykbcaia/Tex/pG+q6SGLjtxANZhbWQ1OvEegjkuJsCYdZ8
2NyhVwnTJswk4WO+T38jA/4mQj+bku/spXFDbTmDpr+MrlTqRPh47GwBCGIM1Vbn4rc9y3I/R8bJ
KhFqWfyEcFxc2t6YGTvYMm8s8IqOKD7HtZgmcuNclTIPhHD4Jnr5yqBYlEjl4IPrSHMDpyHuvjaZ
a6dejDWyo3k5dWBxOe/LJnvqJ0cSp1ek3K+lX0yI/J9lROa5PjFW+e4OrDFRCfFWuC3N3CNlj3tk
ptWFcc1GdTXeg1FVcuQSciYQMQ3YyC4WQVs4Nv0ZWJOzXfxLEr4RCgwsf/yx+nXVRdw/PyJvGChm
mePbsA0sdjYG0NWUQzHsqLeZc39cdUDAQJVGOCoaUWKE6wd/fztsOBk6bcEgCkT2CLcgJS1VxplK
VA1Dz4XtLsN3nWn9DEmMgVAlOfVxfs9rkV58TFpi2yY27be0QTnNPPxiL/UVvyQLpHDh1GZpcCee
Yj/F1VqLr1xQ4nHDJBi0BatX5YFTyE7mqk11zeRlfRnZfP+sulyIPF/Hh9gaA/6qQgYu5EdMdiBR
tVNjptR3i/7zrn9V0pjYEiOSrGcVYcLQ9ectbN3yTELs6xLh0HwBXLJO3eVnml9ykYQ2cs4oZkjs
12RYlQ06FSkKIveUG2WoTj6JqryXd7n8R7lhhUERj8XVE1hE2rD8hm1itZ9de0ia5yX0gZohuyXw
q0cmNNZuTa1sDCjANip0u5TRKxkS4Q0rcHL5JPCsmSa9w0xLAVlJqsqG1FjUuvwRVCSUMtk1+UNa
cF0fceV0G4aKVIwF4APMioTS4p3WeSjHk79px6tylCt2g0nHrnBcw7bIblel38JGLU378aV6CRZW
5KsDY5QYeNTU/evCEAQCq6ITBf+C/s1b9hwpkAYX9mAKrww8uvwmIx7hrWK8GRYQRUZrYfy4lLET
46VgdT8c1MDQda0nFQWXF6a69s9Elnv606lk+TsmtAzzOcFmRnUZVNW73BiOmqwI9C9grQhBd2Cz
bLk1uqhfN8ffHW6R8ARcYYHx2UPZm0NKpG+FBCp8/KZnSBXWzwu4Un7TvuSnYXWDEY2Ib3ijT0oi
n9xzy//e5r9+slE7UbLt2TFcxBCPuDk2dtq40I2hQR5wLkZHMibeP5dZ5WDMyLy/GHXBWV5Sg2Ex
j9tgJxj2eEL+gkX5kuRpTWWgsYDNh+xgJSQa0S7s79nswwaTFCQz7YJIFdPwND9pa1BMa5Wi8d4b
r9UvXC9tIsDXoZPx6Yo0GqTnd0xz+X3mmPXfhiAJWMdMnXKsIvfZ6uyUTc80sU4P7nJ83RxKtgN2
aba+2uQtLIsylKLJW2NJDAaKqy8dHCbGP41+lF/g9Y7P26MxSS/fX6JZUOVurXtawRAd/sfGobK6
iJJGeSaKsZCodzwGD+xP7IJ5tyW1zQ1FXnFKPQs1VIcZGcgYXEnXMC/wSvm3dX2gTESW5Y9+s8pj
sYixj/30IzSFrMD+8W4wM5FroXKJeM5HwGRtt10Ko8/I5pqLG2OYMf2mZKyYVu5sCDz2fSuZPgZd
B33YPpYJOaqMttxWIyJPkotsONHUmRpPuAT/aLb7+XMBSYU2D87T3scrmKmi5KkwNlIGLSkGZBiM
FlJswDeGXIChKRNobyOjxVLQ8qdpdyq3mO2eK1LrT2EytGsvoFbtT93Np6vHy4uE8sfoQzroRfFS
jAhz4IR/hdBhvJWIA2JP8tShfdNE3x1J3gxVDyKDQhoM0IKaC2cOZ8D1n/A8rX4uOE5fSTvtE0Gt
XUlF8BprJD9+yzYol4UxSvuZB0q2t7AVVVUJAcjSk4Y9uWQP2rbzLXhFkp3AcCtrzj7bPx5evlBe
fylsvn4tElZvbecaG6jpwLdXuGplMX2iYV3VTxAAPkKtgppVrDzy8dCJPAScWqvIfP60rg2Dv6c5
E2wtcbV69OuvdDGnIhrzxTbtBTzJp19YAcVpVaCDDf927qUKXuR97VqT2A7mujVKiebF53tpdngg
+EXDOC87Zm26aalEZFboRltyYOM5CQqM49w5bmb9CGDvBuG5vPVDhqqfo1a9fbV3b9Bkk90/TLYG
iaAHlXi3SbJ7PON6xbY+W4H346zmI1ljOlKlZfomeSI1NKbNroh/gNUE/iuGkWVGmgZx+c4cYiN7
lxi1sVoceUCUACtcqx0LjQ2S6EphV2NlJi+yJT67MmUqkVJvTYmr1/5rY7InEqHqvi2alkn/FI4f
swHGY5C2nGbGMCv566K8EdUZXITQK8Kxe9e+P5u0U3qso/NkiHptnNifv4CSysuhFsCFgGCngBid
mlCJ1V8wQawcP3XKO0PzK4kjwWZmkSvUNCxFRCFhjyKGECIHP5iQccEhC2dNq4iykGM7KcNujxfL
vsXCOggBqO+4GFC/sfEJ4B6pI6Tepj8Q2yWY5A8bW8IyUkiGeey5CqUB37GKX2EBo+9OkO7hyHRm
f12K7jGmohcJJzMrltldXLDcKt4bhn6t1kGY/dtC78vdlYGbTxKSm1wh/x3y+aC7C/CQpufLCOCQ
RJwLRoqaPgo8mTbP+ANhn77Kmn9T6dFRwJaDNZvM++p8gCwoSr6WslfKAHkMe+5GheTw2UYyfpYp
YCsCyFvHMSSImTAoMcXM1JXj3W77BlQV2qyqji1A9Fyml0Ik7a/JSJI6q1u7wY3c+f54kU/i3tvm
8WBSraAXbMkNQYCqZukNbQoZt0NI8JUQetgFnykquJ85B8SForqsQJJR/oJO38gSMj9c9tRnwAh0
2SY1BlpnjAX2r0rQFdolzGN6SceVpV4touAIJ+tPAo3j3aZPX9JM+lIM2dQcH+Iuj2ckh9KGO9VV
ZtkydCMBQb8qIJiiyVGcTkh9daKnCkxUOcwA9gylXoYHlpzqbZQZnevi8WjqU/M8pOkGsSL2e73c
eRpopiS2adfvYA4pLbsWKu/VkNXISh0emAcBv5z716m6dvxaQfEKCal92C6rhTL4TwFHOhs6lXRo
h0cuhS59oYf7ngi/vOzOckPQl+ggsPb+eDN1Q7Sv3LzTG5eygggTWZ1b+kKcL0SesIn3VLJvpug1
yOUJKumiZeSwfgJsmpH4l+7uohGDvSVelLGRPSgr80yUOJIxqowcm0C5jQfsOzuAmwkTwVF+RoUl
FSwkauikoiPMGaIpWSa0nRIQJtn2HqxGMNd3QZVpzggDGH+5CNthwGJMsT5PqnZUdVWzohzJeQ0h
+g/6vaWyhiM7K01PPKOJBFzQuVihIQ7hOtneUc/a/m4JxKdsoEc5fEK3fUVJfzK5Yfu0Gtud/1Ts
LPgaZzlwmJoIm48baR8l4nxhJ9P7Ihm9ohlOOWUKnjjLxDCCx9T2LFNYRDSGN4UM7XWIX9H0qonT
Qgz7tx+pSlX5QE7P7ypn4TO0PTvQJp39BP9Udoxtyk6bHRxRHTEC8EBtTwwLSNXnhW46jF25h24Y
HjXrRNyRAkfR+YItNf3wujR5eIlxCOaiTwL3Zp9MUDxsgmMqdk1uRjJ/2swDFcF4TtTBMPWuprkR
B9AEF2gZXHmTPqTl6qjtykF0JNjGXit+v1mfTdPK1CTmjh4B5ptVuVr3TB737ifi+nQEsZH27Un1
nGFzbisZPTI8nesDPvg7AN6rkt6Wj2n/p6zYBh+QEyzzRDr0XMhLhHqiLX7/DKnHdDrGrNoZaUjd
/LN26yYw/LsWkQhOUiaF1z8RPYui5OKZGPipTzGliGADi4eEqbymrRrgCp5ISJ8kbg2++Hb0y7Mb
eKFNDBuJqqENpV5Tts/DjF2XM6jsNEhFkjQ+HcPXLIVh1xv3eK4HeuUumT+wFu21MfaNYaZwdqJn
BpsGAo2P7eTS4tW4F2sK2lqSZm0uleAzEGFUM4qloIHhb1DiYJaP+wcRUM0jFPwe16Wxr7+obKZH
fdFO3TW6vd9pFRWx28LRnaE75AGXNKq6/VaW+mnZHxLIrc1pMKRRrnBOys4LquDLpM6JUEgFR43r
QEzmFfIISguNwQxNq4AkuXYEwMFoRBcxmCf8ib40kuyAFwMpY9FVjL1P9nnuOBlDaZ8WLBHp7EDR
Z17l6SCUZqDbrt2OkzEIepKNqZjDkLN0FkeraKWHW4/jQHJkpSkrKPe87sNQ9trHOcHZrzbUBJTt
jdBGGkW1SEZWetl6xpJNWaSRfGw1yAUdvxIcfuEc9egpHbrNxRj+H7hHghDZkjtIfGsAVzHLTxUQ
Iw42ZgT14215roqgyBzSGAaNGvfuSvdhfwxgTtY8XYRb1dZnrp29lKAO4zjljnc+WXKY34hlNWFL
C3TZ0XCNU0//RhNGohCcvGuMEOfzzbCKphU5kaD9S0gJYcbF4XTonyPQSiVGk6NX8mhbLM98NIrE
EDeUmnleq431CDsvk55Zh2RfUONHBF09LwI=
`pragma protect end_protected
