`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11360)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5IQJj49NipZ8M+awYasSTozcfV13fb8oyvt29Y2taL8+12Jbq2k3H1oA
bU1EhG8N+DKBn5aBP6ZrxX7bkkWMc4YWNJUP/bJ5IFOlIFwfPmeqY0xidrXF1z5gL9v1iardJFZZ
TNcs5U2T5dC8gcdhp4DreRxr4xXZ45+gjCb/MKvkw1ScwUL3ToYdz+w8B86IWutZ9khLpNvecxyb
jDRuX7uRzDlbyUyQDkCpe9ExzHuqFLQaeNKqWSOpRV+dn4NZDaHqb4Y++n9oAStF07N7nscvWUiG
gZDQ9+VXuIjeI1zUuvo/Nc71qfvJCIJgv5uHfRrMrm1Y9ZJ9cYeV3lXVrLbJnuS71Ma4fk0WNJNU
v5WyTro1dqoBzGeEeCkLH7I6AHQWnXjLHxwiFNMIQzbZPYe7cCvfAaxbxUIsqxamqixCxmf8BeuW
erLZultpq9BtueOqAyO8XIsYZVtwEcsg6Qidv3pgquO3JWPWfmTdIfI6bNRFqKOXs/yjm+DdGzkW
H5jkCU2pZgUL2NhcXLK4mlRukv98Zv1pb0eAIfETxIEPr3zdwWgTqfzFQ/5p13C12KHKaBuJ2G/6
fYxa4hVWnUwX599/3g9Jqa95F1UrVZrGitkSYYIWUnCdpBXoV4GA5avRqqQ1w/b6ejHca6e//kgv
iKVffmLe3NDpzr6T4gFo7pVueF6sQUULwJ+f8qDQmrw5LSWNc1TVcXPr3rLRnWYBbhwqDzvkGhJ7
EkG0BrOriGD2EIcQD6U2mv5E0Trb5yK5h89wYOrNdYCenNUje3JCTWSJvHs7N3Nqi0sv391C5aWz
WRbA0i6LyhZxRthkftHPitc/7mBjRFE44g8qA5gQUtgQjzgZrMnwZyk6zoVO7nDOZeJuDBmCpr7F
0DE/tHsKFDQYnQSDqUEdqn66skpNbR5bEZ+uUU+HUAOj8e9YqYufOpewkcT2mm6TjlibGLHi/Ith
njTYIUByfqbUjbltq1mKfFlAQUzPJCabfV6YxBZFBh4HLwiCu02eWtTCm+t3Ae9UqeQYm5QCI8Z4
mtRJaczCp6FPJsWg8ql5tJe/TCgju7AEDaWzSQBfzLNdCeSVk1mV7Qe4EHgtAe6uIRuf204VTSYQ
JiCi8jggWGjUwzvnOUewVjiIIb6CiORIcfsqolmkq1hg+ddFZ34nvP8DoJXmc2R8gaL1Aqbmnl2b
5/CcW5nXbDYBlVyaafVLTu23HySL+ezqLcV8o09NsdtuAieokOA+e6aOFh3+gn/gO+tp8jfIMxt4
YyM2pfw60LIprXoZrdOlCfM4XHNsM/p6eLxrYJf/tAjZk5pkUdLnr25Mx4e9q9tvbUms+0vM0lHG
fVUAtIZyC7FL7abiBLr3f369OC+NFj21XKtUODVuZLisGZFBrxTp4lSwI4xoWBCaWADo1FW12KhL
RQc7P0Y6IELkxdxiVQxf4OMPrT3YHV9ZMTke1hDZga+C2F2M7D+k12ZfhBRNG7s43GhMxQobmIY2
D7PeSUq7++QpplnQxxAvfShoflRvRDpzruaFZABvRzjlDaJJHSiGDfuLPXIvigSbBwcUM5A1YGwV
4gfwiGCEWyGGdpYLLpDbJ85/UUxB/YFFuZ7nbE7/0VndXo4TcS53NxM+jOtJNXuhKxMgeQ9RFBAm
AnmErvANStVAIaSoSg6MdfPjqcHz3rbonrvWAXVyVrRjXFc8g2nMgVh2dC32096rMpIp9Y3i/Vt8
IGo7Kr34DRh1neB9Uu7hTrDXfpM2yfeLrRIh9zqp3c6M5h4XVsq3QMQUkrkUIFZX/5m0WjW0mJMB
fZDrXKvcYnYa3AhSJh1cdQ3Fk4Tl+JbacsEuDFHCeWg0vubkRbpWE3q77n0dpjFOg1oClHzVDLXv
/tgQkpAEePUJf0G6hzQVY3piKc9c6n7SyG/Gd3MSrcq38j4P/5BOz+SJ/BaGfk6oyrdzYk8uYJhC
xIWsxyPjXI8bAis1oOjogXYq8kdyBWwjsY+h8J1bntIkSYBdGsusaN1oQPASsOT5N11Y2IRGPslS
ptjewTK4Zas45bJDrIqNTqtrZhuuzl03viX0AB/IxWQUQfqnNI1ck5ZgDU2ZXlLFd+IrrQiZYCGo
r9FqPXXw6ju3ZPIz8B/wDoymdRlohdETuWfWbwfwWd6GC9v1ktD8BkeehL5Uqj5TQ/ux4BVB/j9o
yLMwAu+uFbmUxg8wGRkH60C4iCdi93v5mtlJiNNJZ0DPydYwMx5x4MqH8749p4o4t9uVTkQ95BrW
+rbz1uzDRNn/89U2TzYX6NGqL6AvRWOd4yfbIMemW0qhT2AoQruM4y16DsSdWiLJZ/9ukYJIpQKp
7dKAX5QT9Q56+n3LWFoJsbWa0lhshNny62Ti8HX4kd44KN0J7IgDj4L3TrIfuLgr+X+FF5mAPMSH
yyEo9rC6iJ823Wg4kG+M+K/Ste4mVEhH+He9kAVgl9tfhsEU2kIojcI5wJA3/qjyuhiVcg6TQ5aa
Wj5uy/j+ZdggsiNqV2NpBfIrZl2VZpoNMMRBj52c3dZxuCNMLu6sk5EZoaK41d6KQWkvRFipkz/K
T/zFURYt8hpW54MwxTNPbYzDlZyKtgPQ4SLr1c6rHl+aMQg8vDXF4xtgn0X9C6j3zcX31jqTso3w
A1cp4C5oLjfT+Sj0P1zYGd260/3S6Ir+r3yaMnDFgI5+r7ElQxglNHM6SquY1N2jcDmgJQWtk1ZQ
0FfskoYjNdKpV5lqWUhai53auAXnCKqe8utriD7oSyqkOBULSYGClRUGm7w1VetCu8c/o0oPlrGn
FNv8a5TyLftq5f53fr2MWhvCHRg6pAGImeHMdJdKiFBpSrRp4AFmAIzyeFAbcKvNBqWh9J84AkEB
odyG+wT8tCwYyHiFkkpzy/AMHTNPfNUvS/zokAo6Cozpe6vL5PjSJkjlRSB36BS8BOnC3nfE4ahi
GiuMd/fLSBPOiMOOMVja3NRPHX3JDvpPl9IEJrVLKDRxHF8fVug9Db3E8BE1nxtTg2nfiJiE9WoO
bCDKh7aeTgjwrIa/uUez0YiBlnOKhPBMvN2B025xFOFG1zzcReqPtgscFdBm2GTmkuKk+Spe5BO3
4anX353vcTGvTdGWaYHkIKVFSeYpPjtXtFvDDsx5QDBXQoCJJaV5Y/EFGxs/JcT3EIJzs3SbFoZi
22j+72QNJ3rxUT/8ARILW33j82qVnjFcn9wRoy9irc1zpi7Mil9dJ3dQFQvuRDhPIyGtqG28rU07
GGH3Z3Ron40325D9XE3P6XYFw96wOZIL7VpCgYkZU/ajftbLOJwoqXOt1VjWn/2QTHEsCUlWWm7B
Pp9skvvufu2rgFIR4/2Afbc7klaemuKZNymBRNjeE+tWK8cf/vGRST+Qu4B33kn+5YziNCUewFUk
gBdFbk2BMcrVeYEVQ+ZNmPqpc+R0R+cHLiPUssydVB6tNJniP3sLFauSGpNvKn7TJBqoimjmkX2e
1Vg1R5mN2pIa3MGphavri0FRuyg35aw0x1rJSTYqwAGrbvR0hnDx8gmDYZarF1IE4ORMqs8nz9mg
gFG5zUOUSbo+GPi7YByaELbxr/CF78RrR9w2zekmviQOaTuP5zEDD7MB2T3xxQKG0eZV0+UOJK2Q
quoMhcp/oUo+hjYMsjlYrOcf4jP3Quk8Yd0o6jsYUDYQU9sqlMrdEmcbwJqyIuBcMvzd2ZpDs3sC
nwIc0yMLRpGjLhwkE4lTbOrxdwKq9ivm8NMuTdkcBqCy9JMHlFN1nbByYju3OSDjT0lc8QZfvGgt
XBYd1/N9ECSA2xMwr421N0ImkBSDB9lkxhYgPpqdl068nYkxO+JIYEhVM34ln5iPi1eNmjROs3K4
DRbqfRyBHiccKPjhbitd17PdEKiMtySP6kad7u+pDgA1IyAZMCh/TzOe8ndui/zPnOpOkKvw0beC
41uLYiQJWoYTfr4MZXgSGaH83Rla2SFCPz0LGxJMl7wgik5WqBDaKEos9iZRGPTMhbGDmOkAQzrH
i6YQ5HTOo+DYy9zC+od2kKkZ98QAaEEGAf9pqGBUfyN+VPHwrYdtXWXeDS6cFkV5Lc8pTbM+cfUU
HNwx9THKBiJf8L1oj4pXXLrPsZFC1hJU8atAlda907c2X04ipMRKRRjg6eKKmAwOUixxHp8So0Px
JpYE16Hn1sekrgQ8MdhAYHEmuffiFGKmH6x6d/PvpOS/OjLZwoGJFRKaRLbFwmEli40qPEleTPNL
98iFkbx7DdRbdz1ZMkEsqVsrxRkoCLjyko2MRS1MRmOFekC7/Vk+aLEl4oUOiTaRk1JVMPeMNNlf
5P3wamKstEiSfXUOMruGpHN9yAXnsvTmtwG40V9CFBzB8dgKnCl5cVvYCWNdu5x/2j3FJaaHEmTB
Ny60AKM1n92Qsc6c4WqvVTa3Zv+PhCJRx0menf9yZTPrWTWUcSkJsURYA5hLII9TcZ9R2qpSzF33
8VtaqNuYTV27OQlM5NJRkI8nVSEFxwSzJtZE6oeDGqOL3YwU9nvzoq4u/kvR5MepTVIcJoAI2mrS
0EzlMnSrWvM15wu7gO8U5mj3Vw0mZasfL9TEw8UbweJcwjwFg96X4TrSnkJJP6CCGbp76CcD0EGo
IC4HjaTBUmIuKe3A/V7k3Jq3Bc2wWvnlAenygaW9MI9CKQqigu3bGPZabP3GItZO+eHFv1p6hBiM
0lI7Yma5PBUrtfG2gKbqkWH04e9ersdASOrQv3RFhjIvvvEF5DzzYd1pKfOJg0zAemTSepSP3d9x
SIMefV4glklXNJLoNXO5J3cvdA8UAWVbo/PhMV74CK4M0VGuAf8n7GYSP+CpqndcW3S88TvzkXhv
L5EpVpZPnrw+gsAMCJtLVKcZ6xXNOYRTkuGzAe+Nrj2oQb/dCFw9yFWbGxxsV+zfZG2s67TKplyD
FEVsKuA0H4G6PJVd0+TCaDIlafrcP8D0ZqjqkIRqBmjM2cmAd9zpvap//v812wPj1Mab5G8EP0Yj
Wn6GnvuSOkoRLrFcQ1D5l7witAgDnQEXdA/YIf2lz0Jtb5moUrKftvrgTqhLmVNJWmykSflX9IrI
ujiWDMu8XTh31MKnfR90wLvM2xSo+FKGNzzMV5OfrDFWxT4bAezW6zx2I7EyCQ+YjtLlNFWlA50m
Ht/V71NYDrfM9k+npL2hkp01tGlGOCKjKsh5/lVJDeGRRf2Gfg3yGxXv41HF/IYNtnVwn8LxQ/7z
npNAm7T0+5njaEg9D6LyZ0Vddu5wZ1kt0kFfCCV7oJHgG5OHVPiLRIeszJO/Khv4nwy0yGYOYwxL
B+4ni578+FIjLAEV/VMRvY5zId1fwV1nDyrDy0pDaTvs+lFKPxpTZP1FeigVNuAIpFi6AuevSvRi
waD3HALpb3lHXnjpSy8XKJhIWkZ1XHY1NBNq5c7Wy7Ajq1ZwrZn+q4vXQijFYPndH5MXQOtUS7qF
x0p+JZkkS8Xsd8SrQ42JiWMQT5C5MlXUBGjjnWTZQEJFiSFLWjKL9qg8TDNpkTAFrXR05ULkYhjJ
Ad8gaxxehFq4oKyzaq5WGOSThgmc3JfVsjBN+JEE9r9WLkyC74p2P3UYw9x5qUrgBXmoJ+LNBson
JPdFMPM0nFuJc/LuAoJsXSDr8RJEU4Ks4qBxJ3iDiF1mnJYQPVuskut7rwYtseK66VHTl+eA2K9N
wo0rNThnuPDg8N3OjYHDCITl2jmLO/QsBE1UsvmFIJ9cxZhQYc4Q2fPaol0vIIJQasZBZ4+wcUAw
4nI5g40IdyhnmWBa+i4En9uvdz6n5fIaTCcL8tpLqqLO14piykO3KnGb9U6kpVqFJWiqIdoX9s+R
Mqv/dV+wcGF4qXk9KGbHzWvNGwmwUfU56HZ5pDJH5APuoLJoAFx7vqde3BZj4qSEgESzbbcjshnx
qQAPUSoNUWD3VYF33UO3fpQOlKzOYg4vZN0fh4bS9hiuCTsYQar/fZRWsDTmse1ZkqkW7awCANKG
SpVlLNHstJQHM/QshVlXTQaMidH4CjLM5Iz8m9zkltjyajxdWp8LdIcDSexv2MmMqmbvoxBRxqzQ
lwNqEnKghakhQgSdwBGcovC4yN2ywvpWUVqrxPirc9dHK8/AIbAikNIZvfSkOWjrg/0/I7RiZ7Yv
9HlkiFcrd9wyaHjoENQVOEDgHF9edEuCf34qGyrKjKzaVXKwW7W37GlwJVv1iLqGa3oXPoxzsior
gBotBo4h1B/KbxekvfFObtkGt7J0evBrQkw2FTCciSt62k7aZPc4fhMv11ti9QhGlHkZxYETgTwi
uoZUjvefgXkNMHx4nZBLkyoVDQRJc/GrSFdf92rNqC9cAD9TQNTd60f8ULoxsgsyYOxUZA/a3KCi
wCNKoE1T9YpRIBR6XO+qOWeN8owqAOe/f/B408c/fJjGmRKkQLQTe8JZfRv1lzPNRQMoNORyluJv
3nA3fzOKud29+GDzaVsj7MX1sMqKZzkMdwoF1cyUyQ6Jsmvt/qvO0i2MWFVKDkwRXVI629XmZ+S4
zsK4HGgytlc9AHz0T+tXXI/h9j4wZhYjmepmX8Doq/Ec2QixANpibDk6fzPFhjOYyS03LsE4Z44L
mdOrCmQURGQgDZ3OJXakddGOwciSIQ/dPLapStxV5obZiTY6asUU/VVEEoGDMmNTpYm7FMhAkUAM
BzMOnbCTAKw8+9cQEuhdC8IYj4tcTJR/QiEDlCDG0nz/NA6tUVCXQEmtSKvW3idR8423Ijj+PZG5
GuPaPpmD0gqOQvURCDXQiKxtiY+6yySoTAOqWne2C+vi0IvhyTMUuzjwTxSqCrLmgB0ZKcFgv+Fk
ySYimxSR21Ua/NzmiFfRSoNSPGv/p2a7NyfGncTXQzi3uIzrJtey6r2c5ZxTrfLxVnbVpQ7xeUzT
h1R5LQcAiWXqQka4uLewi9R9QoKwGkwEZleDSMKoycpFqIl7uUe5N9u4u/rDpsoYMIyusi/qQ22Q
P/5E9YNpkzHIQS1OzzUlhU62CkQaazpGe3adQzqdT33A2lpDeOgjz2DUqirGTrPEjI4HgoBgrYV+
XQ/lG44TnwZa0dN1+Iuoliau9tFu1Z4ZXXcVgMtF7NT5yjNUkXz0JYVRCfyGCYjuUgsrN6fU8GoP
WglIZqZJqjVD6ORlyZyUFeDb/I3kW9mGvhyRcFBbNzAYFYaYHRotdTs7rxlycvq/maHm7UZr+3uE
cmkG/Fpa9TxDDsSXCHwwNCt6pzBOiNMa+cneiEGARl6GHaDLMok3oywLrD4EfM16e4V1WvxaXYlC
e3qDixdQoDZuFSEygnxIACvQWwrA1nZNqxNqK/uRiVvpRuLnCpZBOAgeLQfI4Dm4qe0f8o5LV254
AulYlWauXIJoa+3PXA2Nw6862glX1g+n+2yYdWlaB6nij1lkiUvPRL8ENGiPHTl37pWQ/cT1fDRk
OosVmCp0yd4GV1KVmlnFQfBcgmn0ThhRyrAameMSlCSKcLxxCzt+zWLcDzf82oA4hCE3Jy+qcNBB
ELEfk+AZr7dHVjy8yu7w2wbzw5iWgtpEc9jNGkudTjcNx/b3jUO3nPZ1Nsc9jkU+44azezFs4tax
3kqw5zwD2g2xf3Hw9MV8RrDoa+JSXAUQat2fTVPTbwcMpJ7O4c4Cvbs3Zu9Sf4GICa+3/AjIUnfc
lxidQA+BX/uc3xslq/hTkTlyRelZsICVh2Q0tCtyEjlxUxddDSeI6PRBKXjBX92Klv1zSoNzKi2P
Y8M4mBf3N4Wh0rNaAURKEf+oOzF7niaJXglPQlczNoXPMO6WKAqpwuuRtROjVyOzlmjkoTIo3gUy
OoB5K9XQHp3/aVSk28htCVqSFmsJOR+Yp1IDvpLzB0ep5yfy479x9Qh1UTur3aGj8pbSUNi/PlL8
6raVBA4smhKfJtcxnFrc+cQtnQ3tHxudPF7FTYXk3cYkbf/tlBz3ZVAriG9rryj2hE2K3Jag3XVe
ZWcG/epSe1iAdC0yoMWpP7KbobbFQxu2Fn/FQ2W/UP9CqyxmBKtB3sJBUkMcr3HRQ3gMSGOi5mnh
tTUyY6Aa2RxH50+L74wano1fmmKq6TLujN5ASloDv/bpVRbGtg4Mu0MeXcBD395scqCOIk8zhXT1
GuWB3Npum5wycgn9vG6cXu4zixkaiDsPPHUcgDhQpAJMpv17oBUxV35xicFTJvgZXLV0iV0kK0ml
qqnR5sVDlUAlsQKZu2FNtqGvvnZwT2KjBR8KsBVxKxKCRHqwt5WpEI0JJbaCJPwEmh4CBlFdEMJB
+KLOLA+cG0/I9i3SKlPD69YGLEM10yfdRQVX/UsAmcy6FBKdZNpTqWGGDiueSkF79BS3sKVHLuDk
+/NqV4C55u2DqSMhFSV+P5jsqw6AdybQBvcp1ZRcFIA/hHyAfZUpcSIuxK++/qHh6XPlEpfJhogy
IaiFXnZLQbIVOmq36NhpC9wp8g3nxLU/OkdecbE2BuJkKLxQv32/R8UhgVOebh7eiEFrIaqF0djh
8EAivhDlEZVgBhlut0XU2rQRe06IXjSR5E/3kmDbYqQ1bZ1ZAr0HiQJsCfD97+U58lHlIoCVE277
dXx2DUhqaJ1aIbCt5t+AB8udK4LWJHwz50ho7DSeWE3Ja1SCN38pf+I1dmGJoScEXjiKRjSm4GG2
KfhKsbogVXJUHwfeyIsMdMEJdPg1UjBx2XbLydD9K4ehm4xqQwuuQg3AIgRTrvl41dO1uYiJNRSm
tQnXYto1sNRGpDWpsoDK+ynD4pDNjuAAWOZuiVK1DNU6G8ncrDgOw/Rypj1NmVykqtQntnBw4Opz
sbbhF4LIcLNH/tMpnonFotlccvP6/GHRy/fDyY5/qBTh6gEjc+qnvch4NFS7swQQucrthqzJwXIk
5os86CPNLEgmwcYPuJarvNKiSAdmKPN1f+zCagGj5ew1quWdlhFWRH6r6W3AAC3P4AHp1s3nfzDH
RBU3NDeuPsYl8SqND9C42kkyoFmvy1+Tz/kngrXgQ7HxWA3oh/DI1/7BpiT+QzVrApdJ51BR+iBs
AgxQNdrpbuDoLz+zQsW1lRQ2ybSgejItJLpsQmAMYPTRtqP2T2388tqZuh2CGoJ+DjVuDkVmBbY2
26c8aSQ0gj92YbdkC879xiRiS3p9jecGjsxdlVRcCpYQpcl3AMx3X+oBi2BiAqz2oqrMNMW8ETFL
x/ESBXHwqC2ShEGhyYvOGBIvG1/HnaCN1SMIX/F+8bOxLEyDrWPP2RziJXNRtqoXCiAdSG4UcKdm
+Ivc68Ote+9geyum2Lfzha3vh8hVZtFbhhX9eUkwvJOEaRBnQX45MV+3wv86ZlWnua22YhcTGoNH
SzkAvYM06Ui2sqVp8AfvAjPOWNghT6fKntI6ASwYrjzvVdv6nsQk6uXWKMaCMhup3/JgIzgSOFfr
2raL1OF396DEX4IR+DYfquuCqrJHdLq4P9v7ws4Cztd7JHK0InAendyeptULGigCoO8AW8NeNO2O
U7r+iSMCnb44gmOQQckT7/nkDZ0yc6meV+Ouj/FNDmOmk8oGWyfGJiw1F3P7ys6/y7Ad9wrUypfJ
8HGeO6ALWFDGQaCEtytEkdLftFm2P6/fcGhJtl2i1YovqX+Cx2Llr4OiJFcEidDP2oXQn1XH/hqM
38zYSrE/xzMT3tlgk6a9pLGqvPi2MjSz34IuUBuBo+MCSzeYT5K8H0mFNwPbfoC1Mp6/jGnIuB7D
yovLknJ2uts++53BaKzD3xGE0MfO70jx8ZZXKM69Ccrmu8gy5ySpxgv7p2mjiOZFXLws14p4nbDw
Bs3JwgCXBbHpmHJ5BglayRnrwEMeoWUKtdVZJh/cU4ID9MyD/VaU50gNTfv7PnQkxrYnfhH9fWfW
PcOoTHv18WruyR0WQkBfaLE9i2MhOMS/MT9blAVYwaURKt7sZUuhlX3cadnOxJXpVDq/Sr3sQZUk
0xZMd3nOjYLb2lajkwz7vdp5YZ8juFlCkOJssA2zMjsUX87x91lOrK77HUeb5qHvA0hbhE7nm52R
mCcaxjzbrzXDSu03kaV585Q3SeM9+9Pmn6zacHooMtayJ1KkX9uzgwLGdn4EvXjoWCGVeqtjKYTx
0DwmzZwach4yMdrp2e9ifefnSy/yd7rxpdkxw8vVybnFCOqTCvGojQWxpEFWrpZAx7x8Gl8f5yuf
ZdlG+eeILRvA0iXQf/Y2V8Q3maP/YgTP2Fo7oaD5iRz6TTdhj7ROX4j6zAxflBtPPZa2a/6zfe1K
rlcIppT2OcD02Zu/UOOqYn4/mRJgA2HpnDNowcwKDYLQU3v0Cvr58hlcJpGYdcq9w0mXNHrb4Lz7
34b+CIF4HEeV1ixvQwMeOPbpNRlxrnSdiZjpxefbSdot7J3oKJrVpfLv8ppljg2txjYdZYmp6LEi
1r1MbYOh0jbeuznd3wRd1ZLzkuQ4PY+zWQyWWhUxfy87yggFqMDYJrmHIZGhTcyzdpxK8osfqezc
rj0Atg6SgM9Lr9YtNVx1kkHUHd/4nvYubY/99ubYRW+Z2aCuaPqPpri9rsyNxwHkQ5qmuzc9mTdn
sl7M6UAajsD6yyh8j1WtMajk4NcIu7Yc9TslDnv8UOlIOk0vt51lc6JqUQ8hRwO4YE8b2WaBQCEQ
18Zx6PN1XUUQ0a44eAv0A/dxnSb95H6Jw8WKd9EB8y5V+80lTGDzVn1BqaSn/rXvuOFhgmkIZPEl
rJnUX3P7ewoVcBW8CrYtXuB84dW3onwdDoCXzHk1jmU3s8LjFHkpaiyRGQ9/OtEtKPXAzGG2JgNS
foHKF701MgBaIfVNsXN5Mp4yU+HO+WbRJdmJ98toYscwYbdfTOZMT+OluTVekzLIkh/PqHltvvp/
RjURXeUAGpJiXcLhPqgCUS8b5mvCIhNXeEiROnpzbn5jiVjntoLyMYHKtRW1JUHup/vKrjdqayMh
0Oa75Mh1PTWCsYgEEr8D6faGaffMCZGLXXWDolRAn7Tpcyy2mrwn/jtq+VnDID59t/JIzyRJStbs
zcQI6Mh3QIQJX+lxlvOr/mBDL9TZQgFsGH4z6/x1vYfMS3pGD8CrHeKUofA9EaPApzC1UPXt81Be
9ucpg/VnhBVf/a/zTBD+O23yrS4MrN2E+RGTGQZOnBiZoBsPvFonTAv3Hg67LPbhDOBBkPVF3+eR
ezyxkBjdLAZsTe3VrJdFKykCect9O9P5LgmV4X1lFGF1DjoXR2woE/d6n0uXJvxMaWRTxFzqRqU6
HEY9tWO5bhUfFj7aPHgiAnzMXfLOHnkFITC1TmoVONUuEVtEvmGCFiqYOYGbuFJ6spOjsA09W/ao
46bjFxmIp9ecZPiO8kVXbmNDRmDmQF6I69TdGgM4MNX/tqXBt61Y7Y5Gr+GIshj4vIiWfhdTgr0Y
fkqEJAFC62hOUENa97DcWVicEixiXtdcv0cvcSQCvmxGW38g6d0VMp8UPY4VXSkLJujmqmWOL1OS
f0LXiD7gogh7rW7Sn3BfNf9+Xaofau/4dOfrSfv5jrWlrx6v/wi1Gf3vNUd0689zvKhzCuaYEvLn
q+xEhfxKpmpqOSTt0UqIBfILnctAKYKcRZgSCUWIlDLILCC+51LIAjUkzBUb2BCYww6MuuApS5sb
KRuxHyz59vBHpCiqNl8ZsOmncU51y2OzL/yR2HGDDd3xRTMInrbOD5csQa10MTij+NSEsjjVo0io
5vmsMnl3Fk5LRKnVd5fyet40nGvfmxn4B8MDSS9q7j+DuR3jwprv8Z7ggigTA2opEI/o8Rr/gP12
7XEErcdXd18U8EPYcXzxVyXf4H5JQzUXjt/Ygz5m0xAzuuv/0HQEVkQxdSiHumtBjNBMolie64Gr
RgXOAhg0ZXMozpwepd0TcauuerZwI3x3FaNnkyrMpCdHQjyyR/Yf/+mruvbNVzgtFqr27pT6yLl+
MI9Z/l1cV3jfYsraGLhLmwwUExG+E1zSfOY0R+SgXZebHcxzlHSGtGKzGHUEGdOtwielgtS+h4rm
yWh4ViyLla3SnprI8F+d32tgvutyeu0JkSbMYpIMBjIf1O3gzsfP5Ghs7bEk97UJ58lcXF76T5/9
o3fNMYc2EhkGXLY2ShG2clW5D0JYK+YLdD+oRtKPGwHWV/EkjOm9gzGVcINAKgrIPpsAjD+qSHWu
QxQ3Q3HplFMYebJFrpf7VdxazeBfIhHoiGBkN9hyCOAfSPlCIcC9s7sk2DGNQRm8Yg6+L1IKcdpz
X4Q8hHAQMOyvXzrp0pJBLGX6hgKvjhQd4KY3FpZtwS9kKlG0+B6VTBU498Oj4iyCqo0dwj8gyxgE
l35NcmyZ81L/kUMbCr6j51DSjrM1u8p5mRPEhhq8N4NTXLCU7mBuicKPiSlqgfvtku0A+KMi0I5P
GFBaQFbYMMEMgRJQkbkfLbdcZyr+dldbO74YsAw6wZQCe0FKHQQPHuCZZDKz1QoLUUp6gKxaKG8D
N1q7l6ES9jYRwlDaH05R7jUWksDH8CruzATQRHhnseD4vyVlRgwPHCqLnGVm4Hm2BMpyh8fNJNhK
4cW2Pe/sTJym3Xc3vlEFy90PXz5LsQZvxwGI7OpcLWii1qyYuHdqUZdxEPofj05xo8riuncu8xyd
u3ZUMqxMZ465RaJhsxHaLU5K2uKci1fMKw8Uje18GiOKS7AqcMhymS0YPdXd6oRKK/6/My8W41Z5
gmioj2HydfIOkrHRfiD1ZXewTPe8TX8tsSesGIKZSaTMIwfEUZvcAFN3VfLEHk0Qig11gZk0MobA
n3jxha0KKPCKjwtIgbpOvpmHzElJ6c+38SS29Vb5TPPCKxVHRh8/p4LcE8OhcIfdaKABncRKwMXU
jwZkmHgr3eIpHisIpbrVqH+PliX9vkoF/YNkcgpdabNiDJYxakDGChukqph4duTYWr3swWv3Ccau
b3WHGurFsx6qu2Ke94plgtHUotLmc+AWAsDa0tMOvnFmQiMnyhJY9BnOibLkk3oiOXJtrAFUVwEy
enNLQ+eTD7tRqpItF2PYSOraDkejd6Vkq8bIE/fybkGMvFGzpQTy8e+ppNKku7xlKkyAWGizSb/i
ksscY9bzaTrKzKCnljvrclguEjoK/Nkth2Q41eKJZNw+rxx2SPr4wDpMo9LScH+Hmdl+TxvXeHD0
2Hs/W4fZGSY0a/AB5YddO1hDEAAKVJKi36B51EEIGSHb69/BQCtzlHD58+11c1S1jvQabUjw8+E2
T4qNCi9gSNTUuoPCmaexa8OBkUAKUOD7bLYC+jCxIGbqIpBdinv6RYzDBqJ8viekej5a/k1E6Y8S
f+oQW1NGCoO2bl8h/5QuwZRfghGJEMTBExYNw/wZCLMucV6q/Ac/H0AkUz8y6OizVURhTTgEBn1R
B75n2XDmN98RfQWYuJ5JAUn4wEWd+FsIyjfV+ITnJrD60cqInTgp9o1ocbbmoRFSAaAbWys9AO8O
XaKbyYg+9u9cymSknDaX94SQq21+B9Z1eU+NkF+gVlecYa2fgMKAdt/FYuYm8pQ0zQMc3C18ZaqL
isB3JlB4g9Hxiho2mfNfC4wllBcvStFKyiNv04MtTjlCZXjRSEGy5WdPc1JSVkHO5VfluIJwKzLJ
NLcvYPVdOx6A6lWtJXjbk0n2YQO6HZjhAyz60naXutBEUAyAas4HngBvoeGdXdcrev97tiRaASec
5q+L2w29zrFMACy/bEagJhVcPBAAjillGammnEGWGbOsMthKvisoZzRYOZRpX4LyFKCl/SJ6SQwP
tdJ+q0YpdT1IHb0ggbh2wvbq9IgUnSsBz1GwYK8mX2Tpg8KWsVgzMOPtS9gFnBIlgkuENFS64J4E
i1LXGw9gzp9l7vxQjwc1bSvQN+XSxStSBgNuchrf42bu6Q3P2qbWhHRuPju3sxowIgykMTVbdIIT
iZwuQWddpRfPMhUsGr0Xlk0sIxt/vByOG2nMZT/atpIcvuxZif59KTsABCT8bPukpLbUWjkbhQxw
c1JB2bDG7YAld6nv0sckkjQVMqHT35ot5CL0UNnn/ZfpxEtq6jvjHJp+W/B/wYOeZk8FUvqKmUsf
WPJ24BQGCyC46d9gbwctxYSoWSsMOTlVSW9OTw/p+Wmr7WLpQ3zd6h0sUJosmJPAHQLIkiPdqyzc
9ULMHAZRki6lcnJ73t1I+lRPr3Y14PIvc9csjSxqo+PuGnRzzD2mbnvaEAvBQICF+rrNoUHa4dQB
cW00nd5x5SIss78NM6tuFHGzeMy+LRpjLMibVV2J5Fellf3pBlGyRsxHVRaGmcUmmOF/uJRV7Njx
JdmzeDbEi7waTeBCIsjdBb73laNjrPPbuL2a+dc/hEFOCnhkgTlyqJTph28W4U7sFzVVZPdT8HGN
hDNptSh74m9+maNLjjUf37owz5JYk/RhMKE4tOdbe1wfnEarq6xZ0EZfn9Lfm/QN/A3+r3dr1OSo
xvavZk2rFg/c1aRxXYlQW48luJThPX7WAFrFtcchJqb/xeQUBsO+4VCnOfQ3bvoEIoqExl+SxhT1
bsFwEv1xnAUWHewHtX26ddgsz59TweMLYgnIkE7a/3yjwXmveppxKG/3Nv9Oc1E016tYWlMcHya2
1RM0chofCBMZrHnb/tyjnAp+tRkprR6grZ3SZ7Y8nbu9iMdMR55hDY+txQEV4CiiwoxVQC0Uagk5
KR3/MjmKsM8p+/2aRpdkB8H9sgl4v+QlztM8ng0x1aW6kjw0koIPFdOxVmRnv1qkHtF8fCj39IU/
/Pv8y8PSI5JEWobogYIEYWonAU8DN2SkMr2z8zDTiOCxbH7MHlMWgsfrKlxPHnpRQdYVhUr57kk7
AKavxvHyX0cBQcVAPCly1u6qKGefuW8vHc7k6qAq6AOYfqeIOgNrOuhEMuT8bViQFRKW8rrPH21P
0f6lx3JzfpZZYIqJyU14TY/htOLXB+rVPGwa+0ckD3ZNAH+JFCZdZZCZ/ZnMNa9Fu9IGDtBwSlG+
tiEAqFamGmuJ6cwUkbS7x4XqO88tWvsXDvQXRZRqKSCdDzMw+uq4Lxq4CJv6dNOyY8JBtVTVuBAL
K4+Zb5/1MU9ZDDLhn6C/jM6yNGe+wQFBBiLb8VPTUy+nDrdC4COguOWfNmEAoiNiU37ae4nheAbT
vcZ4ml2uSIGn34w/5VtYgSE=
`pragma protect end_protected
