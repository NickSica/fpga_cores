`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
V82h/mp8FbHcv3//3zVZ5VW10Mue/LSt5dvjsUkiSGtG5WaH8H9Fv7j37k+xy+3/pQvfXcpqBF/k
iaz4/vETUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n4WSOWV3uUjyMD/l4IGcKD1bHONRRplCKgax9lu4YRYlORLHEpckVBvOD9geZHtnlLIjTLNUcuHS
rc4oO2K5x66eEf5+m+hNzaPYWCrVKWQI7/tyX0imMAsD4JQXzU2CP3ATsQoldRyYOQZmggmbIMiB
stLQ3uoRuVc4t0kXI7U=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zgo3FUzRcS1G0FRTCr4C/JBs44dp3dv5CUvkYU2vM2fDyGtu9ekJcjDXnFGi3Qx2X0BV1gEyWxsJ
xqQkFlu/f/1mutspkUjOMtKZNCgPGDHkGfwBEPN/xT22fOBwQJUR+Oj5KSeDWe2U4t5UJ4XXcGMb
ZV9syPFreDWYOTWkkl85cAKcf/WXC6oz+tOUowqV4nSLA1PaSrK4ohf8oaOGNVX+4Ji/w6ViTIJJ
OqmPJQ151npm7Kbt4RW80tp1OmABkNI+o6h4rwtTS1IHzM6bJ1Krrp0V+2aEmmqoZkuKINjX5Pw3
P4Vi6iUmJI0uMpdsCPr3MEC8HH4v95WCnjh0Qg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A45QQ9IEoKpoNXpmniz3AuFZmGAAZIhtA2hP4/pi+Iwurx8nPI4ZkKpYXPnn4DfH42bSsec35aiS
Ve+A8f1Q00bmFgtclspinRe4YgFesk40ftn1mzy6g6sLCNXhUm/IIjCSNk+ie6jVQS7STfOdio+z
cvSm8QQePoJjzlJz/jkNhsD110PhDAevJWb+C5fforY6kT0k7ZmJmE7btahod6wU3o7t2HM6+XGU
DDNZ5E+RLS+IiJYVCOwsdqQFDuRaWwS0k8Mk4UuDiVWtU0+QLFZ/8UGJhy2ZDSYlL/8TrrsWcD/1
Vku2N+fkWCj38RSMWEEe5TmUHSSzP7uBI6QwVQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b+wEsHDGMmVXUM545W/2toIjDItLsHFsIOyFDid8Fv6KhzBePVZlc9t2c1LfdAa6UEpdqcx5kgIr
+oVEglJG3R/fb6dRp2mvlu6+x0AYh7FK0My5t84q7uKZ6EPBxHnDds9FLGQdMDUFv8E10WtGrG31
lkto5q+L5WLAzYgiD3//MgdbP+aqLc/75XWIRhw/PfRn4OqyBU7xSBeoK9TDxBwOscUv0cQ+dauJ
dUQ0W2ZCXwF6cP5c47k76Ikfu69J0/IO+FTLKMkjAB7Wzsyqbpl6RMVdJ/iYscNROh1xxo2k+52w
4l9VnVKN7wTWZdW75B3V/MsNTrKb2I6dBdveDg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyn/owx08GdB/M0CwlYM5XwpK1DLRGgNdNGvCa53fvz5ftb1LM2R7yhWTTXlm8iqXlg1S70wvPmw
WVO2ZNZ0csmDdQcX4HNMiokrI2gpR08Dk8n3nzdOhqyFyh79/eVJzQItyKMQmJZNCvFfww0mtX5K
FbNe2x6ria5jEBEBp3U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J8WwILioFJtk4e6vNsFHYZhWTjvAMbsqHcnvhYKYzsY6fpaoYuWnjTNNNxS6JYZj7bKOFgPjdnBA
rKaGPLghV6UU9fx6UcBVLjNOj95AU3CZPEjWGC/GqjGRPxOkhGtDka91PZuOBRTBqJT8F+5qIgQR
vO7WJHaKezpaUm2zbeC7+ShM5p4Wm9L4dzJ1OuUGZNm39p9FbORAZNzAWa35wpfJ6PPOgATFMi7Z
sN0Hg00oxMFCKSg1bxvN3p4iC3rVT+wV6yuzOecq97B7Fu+tfvP+shqnUhodTpF0WYfGWHeK9ocM
Mg7nt62XJybi4Tm5rgYGMIIM0i67934etK5Aig==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AF8EDKLpUnsf5U27caIfzjHsL1dKCT4FvrlOxjBwD3ZJ9vsXwbWO+EJTOJOFymKnoSSFnuslr7C8
ZCAbkJJLJrLXJwfvC9hiPRksxuYzuxWrtwsjJd+5KWtue3gL5kHClD8Tbo/V+Dnr3gvKzMRNdFRz
i+4p8dC6/32xR0/NITJMYT1uOYu0oBFDHGLR02Wn4PqghcTR3gQMVeL0RsDhJibeNnf4Q0NsKqCF
7OscDpis6r9ZAFao+mdpLGI93rreTlZvJBUPh2RcpqOjL/8IUv0iM922KOCZ6j1LtvD0igXehvHa
5hOx0DDcMjOoejqJiwIqLij0FB13lDBsu+fjWw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2432)
`pragma protect data_block
BMP9G5RAk03qFRu5UmzfhITiilco13nq5x5Dy8jmgQySOFE2blZoaaR0UpMQ0AhK38OO00NxhR5o
xqlvu8Td8bIfia2tzB7jgd4AUFqWbrwfcXO2/Q+Kv8Y5ZKaAKolguS0o4n+oRfUSJYGiIs3BdFt2
cutjmsjUGaV+FmfLI8KubWGbOVkSA4ovh+XfjVQs+UjpW+UOsK8+RJ2XN8J48llw9YcJ6+DtlmwY
lelNMZrqT05MQzZQkmkNLMc52B+2qiwjECOSeeVu8yjwFoGOvNv+JqET0gDZYBU7o3jBtI/YM4jR
f/oPcFib6TS3tUmRmv0hn7BzbdjuuQ059MjgFJV2T8X9KUv+9mHiOj6qNITAPu1K8W61qfQOvvLT
LI8ftU9+Y7yZGzq02zlJq1I2zzCyl1mK6gBSxKfg57xzfjhEJq0C1nBy5W8Ps7JIjaDe+f+HkhLy
A5ekvd5fky7WN2otigLZNMBjZkfiVg+gQ5K74/PQPR/rfg+noC6uZhoTsplCTueVQLNNwhwjWVxO
s8nQ981q7Ykm5dJMuE+yUUElT0HfggZup33SXIN0lCix8zrKAUF39HZjLCBZzZGsIospdgoJMXmp
6KBSkmAreMkic5r46G658KUD6TOHHc/umbar549XNzIveA2P+V/ulVSqI7cZmyMtHmK4lIo74nPZ
9X7OilUwIot12368yZcGzr/zBEfsohE+s4W+52ldgOHD/E5B8bsWutcXOZCixBooCCPbodb2l6Ok
vj1dQHEmwI6fd4hIX7JOTb9pc02qMm1C/mu7Vmu1++HLpDehmc1+aN1+spyRlwdnEyVgBy46uNM1
/8y86r9uZ0uLkZ6nvjkoTtrH5SjzN9ZMPMW+VH8EHfK4RW0Lm5DEzENnLkwKG5Bj6QbcLm79SE6m
e0DeHU8Qh7/5baAftNxx2dvfV6PzLmuWZRWubfnWXAZDwpvkwc+X/7b+m0lSDExcaFb3hNsmaLFG
Ec1w+KtP/pjYc/pY3jBBlndsvEChK85ODrL7G+PGBNshDihMJtGEYBV5Pws+s4ZOZky4ppIMLw+7
MullMsmDPb/tVlfBFwnhNBqMdL1tTacAefOsWHuyzfpZPOClihN+vex5QT322oimCGdji+Kye/Nx
Mlmr1pTdM0/H7ztStQVAVtzDbwe1HNubFzgadffNa8zTmUE0xm4uxPZpou5Wc/oIDuLhuSOqOug8
RhXcecERRBOuKZDKGWoZvY97vfAw+w1gKiWOBuS71CbY+cXEDeInzO86PJiB2Bm9oblQM9l6+fk7
pq/rZ06Azm5GoJIrdU72CgXk1m/xYp94/eBCPnALBmDfzGx0DE9CcfrVBXhCSk5xkkfMKz1w0iF2
WOxbiWPqy29tgoEB4tJXb8hKK9yjWGtAR/qZtrDmH7rDhBT0kBTuXKjQOp49FJXczcpCrUCTlUNW
2GOdyx4a2ev7nBUxnbRRGEX2OSSagcPrpsIjjzJOlhPdNm6MA0hQfhvaNkNLifwlNdegUck7YE4p
dqZ8v5V3GpCH+poYngrGGyt5SZv9zSx+YHMzmm+YBkrzoyuRzVwybdGp6wOJEd/5iKhr1HvxKF+D
+8J0l0ASQ68Gh3dovBdo9kL7tBhJ+XH3fnpsI1kFDBKlS0fYEE1GiSbAL9XSwFmwOkdlirP6ylJE
9aTUCUXgdGxKFFughX+r89fX0p1JSsS77/OleEeRkOSgvyTfYm0gCnCKBpfC/4kwzZ7zSYIrhL0R
heUsEvu8KMDoHUhBSH1CODrp/RnYpV0DIFMU7Su+SwxAfIUrkp7PP+NqGN+TgtXLKBMVQzLSiSFr
Ha5Ecr58uy0ac2JrPr/W0iRT92Zn0uMLZ/JnfIwHEareSlEl1tj5UpyahJJVNd5v2jxU0FZckcn8
IUMFUpKlARnSLenc1TK+ASWTBR23HGJ4xKGSgkhZ8eY9E+eEFUiwecb+COe84YmOReMrXzpP8EwC
9lF7xgUjaxbZ0GYHKJjLkv5MJ4h9iPpimkqsuO9nkFFBJA6CWrgxHNbw332H00Bso6yJHFvGzH1w
m3OCfFzWEgpdIFJHvd0kZJ4W2tskiIdlwcWNOErLpPkBaODT3ha7CGNYquSmcXMkHballyFkmgQm
/lS0N88XjJCGp/cCAUPiqL87oY3fFBKnCUjp9ZP/phMFQH6u1ZLc749RyJVV/5oil6W8Ct5yK0RB
Cylr5OC1yBQ0R5HJpnviUXWCUp0OXhjfF/BF3bFKJ2pvT4pVZzt0biTdKMCWiUQMgZTifWZAVpjE
Lx2TFkcBeT7iG1KWC1LPnzrEbi9R3Q43Yp+Ld6AyNkcHz0Cz8oVzy8gyUr0YAW/s11Z3meBuFhBL
ymrlOJp9EssqLK7W4WJEWyoKeMx12hClPluIfH0MxkfoDd1gxkDPGzFP9M45m0GWBOu2Xnn8rcjA
IJAMq0ka6xYeUVTae8go4sWI1O+xxU+KF/suN+ldMCFgxzW1hIERBS/k6AjUnxdSHwi1iNWSqt9c
W7ut1QXwNLe/8+XSlyOWzlh4znZ+0QAGyDBi+D1QPS5RLGUhfPvVi9bukjLGSMxomAKHSGXVtSKx
LbvIWptgGeO9nLnmzaW3HurHk5NOxq4q8MmXXnFm8IVzWdFcn+BT0ML0EKL0Zd5R7VyQBwpyzflN
iCpN2G+XJefriMa5mV7h6v66VChb853LMmCMSSE8ww05tZ8nmQJ3y+Myd7nrN1ltWd11aQ2FnMiW
S5Fh0+dMTT9F/LCuQM8vXI/RTK16vmJyjD6/8GMeLBXiXfGJmaRIytY7YgS8VcqHWa54OwBVXtKX
TnVdevkA3a/HTCljsnVsMDtDcsxUb4KNhWA3xuzxuPZZ4riPLACkc9taoBP5RvF6WyTvCnQpcrK6
NB8Y85z074KUWOyHm2Aoal+2ZIMr11M+WbJt8owjq9J6K399fAXTQOKdy9QRzhNE2EsCLzB/e3x1
1Ae/RxjJuB5PIkd3RbiJbbAUX+tDpAdvPvSwp32zJKbDxGbC114gYzQfuHWc4cRjTgLL66OtOqAN
u2b/ZF23g5KKfjEbngPkQ+6wIRdjYK7xcz5rDaE9qXZWmLOG28IQZAQPPs3kqv3CTTtWeLNh1C+G
z6coi3dJNcIBYXhJzkmhYzqQXbdisEElyQMubcCUFO32YXSwDJSYoUnR7rJFxdKGB9GnPQ7vYun8
zphmm1VlovE5pA62bCdIBXPh7lF19s82oHdOkIFh1glpfVSOj1s=
`pragma protect end_protected
