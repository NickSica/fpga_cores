`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
iQbEix3JHZTwa1vhipHlmwS1/G9xw/soq5c1aH9r1Ikmd5PFC6vG8hcczrO5Gm238/UZKbDRHhQl
8vxxX1eWXA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NYO2r/VW0Uk9iILO9avt3Skw+TFdXKrXeDrkjkY6MrmMZXqmt1ljuTdXla3Px6GiDC5iNRfSB1LJ
jlz9x6ZyMo5VxrDlXmNLima4xlcLjwQ5Ldngl558uz/vr1FbORoJ+gk4f03PWwyf42EKOYFnCVfd
LJfFRdBml66XWTkIRRs=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hXM/negBdYIePK99VNL4dA9qZWSDCbIcZGIF+wzwJF2GeTdZiC6Sv8N9/cF1YoJ4PmeE+1cpGoYE
hr+rxDAb1wjgZvfDyEG1QWzKRSG5E+oNC6Bj2Xk8erPPxuHL0sXJnNFmZt3mRdMMjzJ/oBGkUF0h
iYE6DHIS9BMznThGr4tm6wOQ24nLfv2CkGw5FtsfpBEceglyVNwc5KmDZpqUutO1UmcXWgUVf6aG
3t7duiHDJKzCaRYGI47UkrEGgYTLtr4N4clyKbc4ZaAFsMfafXuq7UodHyHPGa7sQYA60+7yMSq7
lZ6oowJsQLQdpXSegbc7gK8ezWVXMGToMCUX4g==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
IZkumnZp/JsuGCxK7A5f04eL3wOhVC/HIkiq9ThWDUN6/jAV9gkhdECfPCdAYxhe0IfGI1mwNrRJ
CATeVriO+TbtGJF8trisSNtrtJxyu7w+ARrQ3i7xJ5OugSeDn5jrGtPVCeIVbs8Otz0RthJD/ia+
zMRiRhN8wPr8+wtwChbS7LbmoKzd361OLqaC8TX6Ab1GBUHFOMfYyAPJdl/jXbS9u43VHuRY6Yc6
WqrfDJE3842973TEArl3DaaLzZwM28WBp6JNk4Z1zR+7/fPjneoZl3Dvksdx4ThM0a5s9BNPAH9V
WF7gF4b9Me6TfP8DfbNOy0URIYx+xbfpe++9uQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
eaRvVH2iXg+bRFhfU/Zdu0OhZxAtLuP0NVIWmdEUooi3G/jC4AtcmpPrp7p/DrHH2FZwIvu+AbK3
sY3ybtP3ICKGUwlnIt7XryFabcZX+wxEJ33rwyvMH3qSJUvv0NnXC8IHlKKyRjDylY/oANDzbz6D
+mWDv16FdHx/0RgRk2HTfCPx8qBZ+fT4hbE6exCfOH2KzbFjubsbEmNkNU+HUDcusYXP2EoAnNGO
lFufKr3GhljOMYxxaVeKpXEcKWjQB5Uu1M3JdONHHSUP3iVPekneDcajTRMfHD9FJggiLA6mAgel
cdhHqUxScYsWsL7cenQphjXngVDIxqnSMZgGGg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
heQDXwsWtguDyBBqy+N/Xr88McxL4tQSR2XBCb/lxs8IKaambMExKMCiF+uYl01VHmTIU2W66UkM
7t9z8H1Gdw289KkEy+LLNQNFvy4xiQp3che0cCrsbm5/JjwMeuGavzmF6wwMkz5sW4oMgRBAsxzn
RRGXDS1r2TiNXhNi68I=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WZqwWujfHGXV7wBEePMjGLVWUeV/ygCmf158CXpAhJC77z2vuuagSDsOpGgtqyakG2cswti5bhBy
iGqPgNkEY7Q4T3NMe5WssA5nf18Sw3LU1MCehsK5WrHeKiMOyz9QpdgScXEE86/e3qniqvFlM2/c
HpI+I2e/HN1QOgChXb7HzAEEqCCdY9VD1a+p15IoOmU/8Gs718QdaPMJOt3XdTu5pAmq/PWuICaZ
VFSPDj57xVELte/pDBIXo8hgI5sad9ci34UyXovDzhRyUKzLY0u+gqRalObdZFD1Ph6hGQiLfmwO
JTvUCIjoFwTzhh0dCXYGcwc8O9kaaOIiiwpgyg==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
B4GVIi6TGeAAKF2mV42cg9jGmUkeJ9TkEGN3HtEus1MF1Zmt7Nh1Y005XEEzr57ufgLlM872beae
bxX2U/dQHyW4OCP8KBTn49Kmkdu8j6t5b8W5HRsXXHYSGPOo9IxUSHBdhwxHpNWauRDmTFNl2lia
Ton0toY2wVDxIcyINRYIpxD8YGHOnHSHPMsgAGtuP7kRvUnSvNzqqhzVcNm3oeIMTawuhFgBXD+f
0S45sDt4HAERXJfO2RXmlDCCLpg7FQxibRHwoppbdhT48SpFRar2SU9FLaP1Rhu4f8UN/BXG8JDH
IE70hcE1uVmlqXL3h64Aaql7Kf0Mt19/bANOBQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34816)
`pragma protect data_block
8fgGNC4HfskTXIPOSZDcR0DhA1/xPSvMbOj8bNtDga5EG2aiXwF0zA3myzj76F47tsOdfWPcBFo0
QtYa6OKK1uX1RioPu9JRVsKPF7UlZZKIRlmxxbP2sHx0y8EImZIH1tF81+kzbp4ORjPAY5deeDbM
0BlLdr5s4pj2sKlD0/LU4iLyptBr7HRbQzcYEhvwZMWcaE/d9yt0lPaxTyu646QGaBJyaqyUB+gN
a8mrC5EcJm7CSCXth6vQ7PMFeipHPThKCUwdkApKWOSaxZinh3jtlZixdRCsf+qQOSL8fEoYVqRW
+r3bjcmT/yPYB5JNJGa72LB0579U1yeQAT6QR0bTG6yDbkB1NLOxrZPUHDeoBHK7O/v4k40EzLi1
K45ZLFJRBjhnG/pR6YX9jW+dnQcy4al0Lt8VUCu6Aehjw3ebsOMMgvFFf8qLU4Bg4HnMAoun2BWR
ow0EuR0C8xykzj1KJ+slvvvM2uTA4CiKhNcATbIXp3xt1/OMtbOOcbhjWVqjg5VcgMBX43rj+crT
jea5uqLPQeYHL7SzUYnzfqvBMIfwdYS1Xu0+UO3iJ9BSmnoaHCb0PC6C6/AMA79JgX0wTImOY/Si
DIpr4fLUhAKxSs1klfZr0sMIhtFbXt3KacUzzDxF7IAm7xFAH8NL1BkzJkAk5mmvH1WrrBG37dyX
lWeqALVNRvvLF4aBSuEPlXjAGLc0j7FM0dSBMGrHvfHabV2+jhdGmw8LyzAaZnLTui/CO6eMLRjQ
tP8jAIHUKyVwBZD0IjQJkgjq+LzwwUFUKkcXRLCydEbJ587/MCF+wCKVh3/2TwQUVJ38bmMWlwd/
f5eOUKrWcpxyxqloxoEho9ALqNgGiA6srR1agf3uM24eX2Hxhi1tggala9V6mzj4whzz673BNvTK
/wRx4C05ngZuGS7Y3g4rfH2IQwToLgj3S72yplSAgtrC6Xvnmyv3ax5nAVMTud3u1pbzWBao60uR
F5cUVAxjhOmXZhl53xuArpf7Uq/WXVP9F4MljgIvFnLUu/Lz+ex7xnplEcHKv/Cnl8SQZLQtULyS
GN3oRvjxIMgVGEHyL8bNOnxsacRnSr/5NUFQoOU+9q7NMhEYnsUyR5A4QSQtwcVNKeWW6TzVEJDx
Td+d6YzkTskJNf0D21kJD/KxftbyLCDHqba/9ddyFatN5co1jj13EUnjAgzbfgOQamRmKJZ6GPRp
iDW/AxHMeQAIHjRkYN0Vyfnp3ohvedKGY6ZUguKdHKwbOrQCP4yjLFBXroGrOjwZ4QRjZOuprIsb
RFTd0+DtSLx7ss5WvH5h3VJJSTBI33Y5CJE4A7n8OHJ5fpeNVmd3wjnWM6blardnTa8ynbh/Zgrd
8T7qQH399buCbIPQ49+EI9pJLjv+DWKY4gS7Te/NLnINmjhFVF+7mi6IkOJbBS9s6ifbsOR6Vgsw
ikPZersvV0LncRrFNONjFvERR7jtyrV741zdxu+rCwC6J9iDKM8LATur07hGoF5apEGVMKd8JyUe
qtZObpJsQ7bCIDrumX31VO8pPrNoQdUaqWoTPdqcol7anDEy6H8FirZt/Ky8SYF4Bg+PPUKdupbM
5fMBHnEFWLCwEhJSlmim1FgDrshxo9pE208+Fqm5bS1fMHgz1QObNxXwEig/rW2kXuE31OwpZzDY
l6AQiuEWFOyBt3Kh3e0XA9TuwccZOW4D8cunlbP5VTRCm+ESOQX0t+zmIBOJcS1fTT4P5+R8hDrF
fzgpOMmLcf2jHBsr7iigdLnNTf9pYUOnOquRQEo/qvr/rmfXpx57BkzY/E8D9dFIB0Dojk74R0KD
Dwp6QBHths+2/sN0WouA7gbvGcK7aXj3bLKGIvPOvxrlaGbiy0BA6x9T3rdYhbsLaJYXUq3q27Nc
qwQmFbsXCobj9fyObWDHNcC/k++zvniZNuWpUbRjSHQ1rs1IsW2yS2GvMrk0I0rX4SkVIWNPX0CU
ObOLi7NoC0qPyf7insjCPh9J9Bd9Q3uXpNTBFvsH0LjKSAAdwe+JaxBY+cMKr+OGO0m+YuOouMos
3vkPBZNQ8qDHhKB5+wPCRxhKQpgAgperPlmgBXSsEK2H8/RZ3irJocmWD4L8GiPn19dIG9pYEfWT
0fNtZfPcfWCsiMC1myKGNd1nGcx3IpHoLa6gxfMEuqWxXwVO0PH/z93/oQpjdun1fatvR/qhVQB2
h2M8I6wPVfz8wg8zFGyKHlYyRSz/3wRB+D8/yX3TevFyYriIlI75FhhcJXElpEkTMivIQmD1LIii
IVNbehAadAqSd8z0X/OBGfVk71VGQqi/3SUwvqTtYxEE3pCUku2BolSq2TUUn1TPMKeVjMo/EpI5
hmnXoyXDxbuoXPLidEL6dTLJyUmu9XX+4feAKPy3gB5GeEXdYfdi1MsLsskYPtA3z5BoTikeoHSc
lIt9O/uOqqswG+yEohscdRMjmkLUvs40HYtuuA8GJGyejVrPT+NENmjmbX+ulGPFaBE6vPmg6Ns8
+mubNdn3RDv0IRQgCW2L3keZIcwZ02DYxnMzTiyEvjDK2Xqklh/jxj/siQHCvUn7S6cD5hlsBYW+
JYEi4CC8wMDohYBBMr5tBsmR+8evnQsH2CfaVANJB6UArYszo0xddPxqlEbYCbrYnL7m4y7KPpXA
1kskp44AS/Fl6T3N8Fh/l1CGWgil1wLObYVx+uy61pVMSA9m/Dg2/BZRazNIXWXNIOIh2yVRK/gj
1xir6ehDGxCVFec61+NvDplVrNC1S+FHL/cMT3hJ9JE1IrKMhDT/Q3Egxk/pw3u0OOVZXZBRPzN3
37DA4sy8baIXiaAeWGxwYMaldRYr2uoY0cNWpt14IJODYvvMc90++yvEKDdJ96NrCIKhLUumI2IB
Gd8JLEp13NY/AvFgX0uHdVlaMdwJxvgW3bDm0e31i+yIflQQVBZuf/7gN0H5ZsPv8cjkPJFMaZpb
FC1aszVGFf/8wtYegllqlGUHwHhDwQFQyyUsUxZAJoFZZL020OY1YhovfvJPL1sEwPQ9nzEGV2bJ
UrU4Ui9NbUyGHx/O9jn8cUDn1S6cYEbPsiCr45Fko2eDv0+2AFYj+JdthTLhC+XaCgI7js8R3Xlo
jlEOhm+9grhtUyJCCspDpp9sRLUSSPFGDezg3WRhQFNIWrqGl9TBuu9qtM4gZPyp2km36fD9FOSs
xjuy7HY2nZwkE/B9zCU0jgkg2TCzVNfJhEVrh5eJf7H4s4q7U3tQKeJvPHKIKvLicDNHFwFpQ0tV
cDpA5UX5XCoIMcu/ha+EYm+4/rKcUGyI5Al6gRe0hHmFPSlUKlM6Swiz17IAhRo5qIcrBVohcO42
rer7yWAh2/4RJnQg/YgXqs4FPcoEOpOvI7jFLxiQaCNx7nUI8TF9XGHbKsSHJ38PYTogLYhIx+t6
DHr4NIAqybK7U+2DPU2woWQMv+3Hq9Yi+anxKkFzuC8+hoIfVnvsL7YHjQWX0gQzooS4TSZP616w
D0Oa9Hy7PREQWcSUGrxnc7laaPs6wALNN69yIyBBMEypTT72B1bHI/ox0TKiWNPX91BB96j0POt0
sOqqhKyvKjuuCAY/fesZz8HQ92b+bFbHVpOYvjtZk5Cv4Pbx4MhpblkFu5/jsUnh1dNAunYp8D5j
jpYPWQLr7Y5K180aLAfMxL6eQAH9jjdbTQnsc4/5252UnQo8qMAiI+shW3AZb/TJfXOvSWepR6RH
uUrmhnK391L2XYwEkKIcxXgNGbk3oe4n2nePgoRmO00j/zacX6AQ55FQmX8FBpoqXEo5ZwXpZey9
C4M1Mb+bfVtZp7ucntKILyuaCAloy7E99oxGWa3/BhFg8J9hHvQ73VIi5f97JTy9sd+g6y178fFo
gCS4jRbWB5Qe6FpVGb8pOVsFhbkWRMihfrYYKyedGQ7EyzDqAJYo9FZ8weIX1uoNVgJjn0t7oJGn
me6FOe0LwRJRtEDp1S2t3Dz4QW98kylXB1OMGPLGg6R6enHiGb4qVD/zs7O36tTDcvK9rZ/nXJWe
4MJgB6+B0hAiHVnVy+Z7NAIi5Yir4wrTgCfYRJqxBKL04dsfus19MPgRphzlXm+8C3tMsWnaMvUS
Nh06YhHuUY2yZx09gePNwKfZb8rlBphvmOSA2nHY24QmPsNuLewa/AvEQpMifVT8DYbihEAA540y
pYlcPLtfMbTlxAi2hpGQH/2if+FjT8ikQK8ST5tXqLX47fIyL1/nyZbn6vyHRtc6lJ1oL0YtyhXZ
DL03sAy8/tSzkcW4scA+EfGS1uGHmj8cSJafaT5BqRn1KtNOhSI9g8Pk9Erx6LH2x5t3ldkq+XS7
cvAqc9HUUetVEmVlB3aYlbs49wccHbKnyRlKkvoPdl+OpyqJ3xSLqGVPWj8/yiPPoLlpEM/MRVal
OHQguRX77KoK8xLnH16x3d/ss8jZRVidRujp4U4wIdryT1Gp66kv0vEq0U1E5rOsp1LHY81SrQUn
WSvtvOqwsi8ibMlK6EHsvXn6eLILMZ8s6Y2pSzrav1izipkBCFar8Du1gfd/qvlG/qU/FUT1Hdif
Qij1PgMg38k0TuNo8ggQhPJtCkzcp/Ap6YfoOVUprPHpwv3USdKjGYDsxeVVZEk5X7BNKNXdC3SI
KOtV/u8cj83iL2ivCw6gJnsf5JU74SvLGMKtZIzgoxA/eWRVSAES84zLox4pP3AfA5KdfwM5Uc+a
MF7UI/gqjFDR3jmTbsXvnEkxn88L17nSDpV/xN2QFMdjl9lHWEuULdtEikcVjEWYJAAKR7UhdJYf
rLs5oPK1kMcbp2gvu2Vi1ceDfPmhnq7md7JdlzefS/T+rpvP7odceNygpjAr/FvZDUmrRAALhOe7
gcU0avY/eSJgcdulSv70gjPyEZF71wNkK2UrmrXohhQR/OrqKl1MRmeisNjArCrqSHcd0b1CHC3O
JTZOqtp1fn1KjnDoUafDqkXtHNlBe1qoXFkMvNui0y2LdPOS5yvYNDRNTEEWYYSA9iddMBbZvRm7
PTslOiOCRHXftvi3ZYcNzz3rEdZdDnKy4kNF2nN1G2hJxL+MONHdbaYQQkI/4BnAT9u7/Yr6eFt0
RNSm0bGwtHAQ/butCDT2ABiVd6lr7gN5Bhtt4clmcFe3wF2IMFY339rXQzaghmR9Kq0r7/zVVYZf
tcqx4F4ocuTaKavCdOwVHJ9TVwQv9e6GH+UlKueRiAoyCDTq85PlesGM8rdQ7CzNXIU7H4WBJUEu
8YuVbctcbMcBM8h8YDEwvAhLZO0bjmqo6CxPo6psSNEQFiFqqAB1jnB/G7PeUQ0H/p6bah5lG3N3
pKEvJYwPpFaiNZDodygu8XxMwMTogcNk9ksJ+xmnRrV3AC9e0zQMh8EZ4pwfLxk2MCpcrV2Ihw2w
We13gCQcOJqRZE+gKCBAcxpVyScazCO/VllhcWX2uct89N3f1VfIU528mR796EwjChSwpK6J7hCw
Fpnx3xF+Z0RyZX1rgXvK2OLlULLx3itjttRgAUriu/7fH6HctayzSEn8Vr7E9owT8MLgeYiCmuaH
OM9kwXFwwfjSC9QL3z8YWEGz7pqyogf7PA/zAcZMeHHfG4qEygJvNzBNws+n3k/35axo+Hqhm2lB
m7S6IGlvxE8KimxcM8+apSrViOPlbbMzTEuqohMZs4MTXlj5Lg1oV5pfp+3sLOy4G71009ZXyZrU
QPoFv3f3vykDfLX0S5r8O1pLA2eB0cUizGsZ66DRKz8KwvAzblj+jx4VLvSVwLQ8WIp9bf5PLVv1
c3GltbVrqjZwPA4UUQ40Bast6H33DfX2vNlrPCzliQSSfYoHpkxvNdkWpk8XP2LNSAj9mKBAP3aJ
J9BYZbZ7g5dn5FEJglGaSSNK5vp5BpqFvnQIwlwYutrpvgjanCxR5TZ63FnNRId6qOSmeTXgDm3g
N+BFArHjlOra2OppliU7TEAL1ELFWoFaQp8HRTimv7EHLNLIS5E4fX0eivf2w3WiYzfOz40+6zxA
+kkza65WG5gBW8ZHAxv46zF+nFneBmWSG5Ktz3/v+YbM+E4nuEOJza4gmC+HITtyYJ0H8ha0Xlg5
tmVKpL/sWkwEp8h71zBVpi2sSJKfuqMUmVXPlPdVCMt1K65957Ty3LehLd+GJs/VQeGu015fgj/W
z6swDtPAQ1M5IY02HJoLB3uBnt7w2tzZ7wHmHkNMBg4DEKApcIH9CZwf0r7oXglDrZLK0sp7vnCl
cJCPtUHZnflOHTevD9JYnR4IKRORGFIh9qSGRVH1B9yZrxqevamWY4biDbZRfgbPSyMR4G/z8i0o
A91BDIHP/0/Yg7F/Z9W5eBegbUglNk2rs1EsVM8mJhFJbaiWZt44nbNQhzPzIxL9JeRI7Lk1dhs2
0yCun4Yzt4+W7chWjBy1j91xif92/AjP0Rt9T11z98tEl9mbiXvFYD3882YIFF59tn7ASE93K93n
madyi56hmeMvmQ0gDSlFhP0pPl1xg6H6Ecr5rHdPjjd6aEqSH5O4KLiKGs934u7jGA60n/9RIKv4
ZWZ4HRehe8h6I3QLdcyDDRWLN/czZCUiintrKDlOwAURJg4gn3J7M5SsJAR6rkKRvRQekJJUoTW+
PoSmPT6WCFNgWzW/qoO/GQWFeNQMN80bTHx18dmlVcxwnuQ96dSz/+YhffsnWqBJBdEsZ9PDdTHD
4i4+pJdVcA6qs6IW9+eHASEedh3AHBdwduhcHdZxlYcKdHcEWVtzrFq0B4qTFZu8oNq53aWePAIe
EXZc470f8h7Myc/czTc+dJhrPKjGndqqt+bgjR4jY/oQcwY8ZeRIL7NlR+BWUIpNrIGtdz0jGedj
S/K1iNAgsHvN5YLU10aIHIUpNMVG57HvTyyCVWo7CfPLcrium1r+wOBGy9MidMeWusTDyPAouGzj
njazL3mYpPw4GJ72FvgsV/CQB7OwShdlihEDhCHarW+TvZ7B0XeI7LWTFYKk1dVREPwl3bEvReRM
Qd1zdcKqc7zrglkf/5ETt8syJQkMvh1aoNWOxs2Ub6GbWDqy+ZICDlxNyJ0s7LYI19OEUd2n41ZJ
dJZlTW2aJDYBFaVT0q7ffb4Jztvo6ysm4wBbifbQRK3PWjtae67sS6J3lZMpMR7/UNwxe8+yyXYV
91q4w0HR4k2BnY+OAYBeJllAdWJTX8bfT38YWmGv460QxGbGJvovwTz1c/Skspw3l5n2hISgNI/P
aILYUrpLYYRor5txiWaj+Zwn4SPw6wtGgGs3MwfRkebkGFWXvWhX43SWBVy75pzvgFdKOdl72V+1
Wy0yQZq4u7vOCaW6Q9nfYuDgUaQeWc4D9GjOFQI4t0tphzUiW7tTdXL+1imHdCzc35SIPV8Wc9YO
7+b0fkppmfNASjDOhhjgA5wHRx6LEEHzEy/4yEM7KGTndjWUX5APGcSiTHnBl3Wpnf3N9ag8PTlb
/k6sn4XhyaU0GZkwu+j2F2qglTr3qzE+MwNSKlYbz6aEbrtYoPPCzq84Wyl+L/VpYpdzU89Udtd0
HxFdzVoTa21unrxRJNDus5iRWZE1/TzyqHPDQ3oGK1nbhDNNdUN6HoA8JEDxdbIZy2pXtQbWVpZM
bCG3T0CPEd+O/EA2Ye3g532GcY2S7ZDaaHJsQMYNXDABbDNCDjJmK4JdrqFgX1pT4aifvIpir18D
Pf2m7TBOlxmiYsLJH3POk/oDyFNArKokzoxTkd5/KtwBGFewonRccqDzS4sCai/RLgagz7IxttIZ
5rQddraZsXQgxZw/ejU3n3br+k70S67jg5gmesw1rAz+pSKXMDKhHvfEwbrOyLX54esyJ5wbjs6T
bOIbrFsQJD0ISuc7eggEW0FCNWlfI+ms7WnsTxJMrvvD/qZEd23dLzu+9V76ataenbEaXJKvA004
f3iTbFbQdxRablpRptRCn3VatVaJ0++9nDAebKW1Ezy6NwDaMnTB4wyyrVNCZcI5VofRmiWMgikT
XTuv/YavGicR2alsW6rM91vKW75X66UcVb8G67fO88e5BOaUYSzKzSKFm1208z4oST3x5qZ2rVdQ
c8Fu7Ar2QQlPUtWJB8tWB7Rmc9Z/0pzPmeYzS9EU6o1Mv0lwTI/Bc1lEX6d/yCrS5qaBrjTDwENK
0BnhiHAIafOglpm6qOa9hwQWQj82NPjwn64PkQXx6Ak982p9If+SnIXAP0+mEyg4L1iEa7NX6X2l
6FV6nVOPwiVmVmNfFmdMAxRpLuFvPikVpYmgRRGhRW2HfeJsyzMm3jp73N5kaB7MBxkRy8Tb02hg
dVh6AnhkLcR8Q5qgJegmthCnzuyO/6LU+QaGNCCZtNoXZOHrwTEuh5+EneMA92vI+2LAX12EBwia
HIDKfBS1J+MhwVudNKRdsxYpVZBsXeDt2lOduHfyZ2Qqhrw+cAEwi8M8PvtOOF3FA6ET/aqDSFiF
s9VSovf02yl3wjUVDcLPlHiYrrMUa5puwCH9Je9PwcbEezJeO3JsdSOh18qUr8cs7jkA3m1G799+
f4s10gqqcPImzhPWvzsnYBZF4PiJzLnKQqtSsOODnfcfB6Tnq/R//zw8Spg2jkyaTnVTD4evtDpf
h3KVAGfMpmw42i0GSEyixwtD6zEhTBA3AbC6jhy5VIhR8z+2hiUtiE0p7obiDIAJZDCUi6umu8q9
rfwDDzt6SaqcE8sS3GytIKAwtKQuY6XLYCofwYMivFjOze0lASOOsc91TJBpaAGdd0Rbx0bXSNcS
NzRnoAP3l27l41ARbHaYdxWDQsFBlq7m6a7bnkqfm3bprW1XCcd1GMjTw52EJ1h9ezYyCmLPJTTY
peqfh+P2zXLHyICdSlVfG1ZSDcmvaKGoU+iZUZpKzxSLMS1emUk6MPQ/oKY0p994t3oxzDlD5zBV
OhC94oNvm6q5tYkb/aU8AFwq1HCLpfBsz1p0AKkuTzalBPOyJm8RGRP0YMIQOhJBKKMWw1wMhKN4
E2O3J7mb+AE1U3P2G1fVssIxp46qVtWry4fcUjF86lSto0RfaseTcLpj9Sp20+P/PlJpIBZQtDeK
UCpKYx7UJbw+RTQ4YoneEG66kusMO45RIixbJVyyD4DiVVuPUjkkL5+NdHtWE2ty/W2aDhLD+IBk
u/SGPoIV+OBEes66Z/VUVLbTlaN0As92ZOr4ZCZQRYin1neMbpwjRDlqIi6LHOItkbD++xxWccLo
b493t7BJMmr4kKn2B2LlfwR4TJ4RlUBmCrad5oBNHv9G+GA8mYEOzkO9IFHK3HgtpPuOac7Xpsir
yCvJYIpGIVssQiLzUu+02s4zJ8ucJdqMQySQAOlxP/aAzha63LhOrSz5G2ee5NCrN9YT9H0U2C9h
Ef4EaH3zpO0Zos0gyuzTpTm9fVvO/ngRM+0Xe/eE+6n1SUQeKBx4QfH7paiiwGAj6WAIGpUcjHpf
ONQzTwF9rOho3HQYWYlbaX6y+mUNQq1aFqX3A7s5zh6uY/o5r78kyoZYtOpPoHg7KW4oIHDVnoIx
MowU+YvwMe7aVeTC1d7yhg0SV/KXz0/oI9FAdqyWoahG3+NxHUJBwM1EYSe/SVgDXN4mc12YImfi
mpIKwtNaMDplYRfI2G2VtP+xl3jlV8cRrEaW7VZN68TmvylBcI1OcLMlaVuckinuwJ4mCsdrKAL2
KMAqJOlOIxGHZJJt5ZW4sh4rpxyfJisNu0gpabWmT6iRkwU8bO4BwKbUuAzAcLuPJSQcO9enzcts
Xl2EMjtiIQ4NRADw3B1J1k5Wph1NXa0z57eUWyYRY8fHMe5OwJlxBPWJjRRFkMaKSmvCeErY8O10
+UnFa6myAVq+uMb/DChwhBAZ+UJ8igGa7ueW2r2/Whkbq23VDxwxRmm9nbZLy5AolAiNtUqaKBLE
MOVcoLCIXerRZIlprmkLFAvUdT1PKnqyf81S2uQxBhLwg+IPRVvjTf2gNx7PdCiHZZbd7j5zC7T2
MmaFi/nrNSOWhncnuGiKsgMWsmFKcxXmcMah57x23LAYhzYYR+8p7UIaPSU+OHdxEjiAnRVRriea
uuHXKcZjN9UzW6LR9m4i2XIfBsiH0ZQGUZvqkyciZwb6AjgLCEurKDenAddwjtcyXs6RJOHPh78X
seohM36Nt/Faw+6/kseLAFPzBw0miAMDG2F5dxJcQG5FiAYxvjYOzpsX4+psHbwDuiVgKkUFESQh
VnOrdd4y9dxode2L6wkL7uYOqysgAWmZB1pkGxlyLbhWu8L4+q81aw0PE9vilXn4aVluHfUZZM/b
G09oP5h/yKH/LCQ2XanAK82qo2u4ulA8qwmg8qNwZZuP5DQzAWFrh4nv38kfZjzoFIqHgqYmcbtu
2tDOw4eer3Ygypzv9r+lZZApoOV55M+NQdlRBz/ajeT5ZAkDfQaJDnzHUdwQX4rIHrCa3Hixzti2
LIfIq5fseVPGYhoqo80p8Qa1RBdyjVnsRd65UmKJ84SSK3dSJTteb8M8O24xnoLL3ByxidhnAppG
vYrk/JNKeA9RIXo8AEMrtZ5X7T5/9CdIIk6y7jfnFVzqrFVRUoUCl2JmvueMm8s6ZNO85z7OKjdn
bJj5Cdq7rRx1LihGFJNXICM7EW/Di6zG02Gy3UbkZzcaKzpHfhsFfHUL/OKBnU96I2VbTWPTIRsR
kpEtiF7mGi1uAIiO+jZoQcGbNf2IF1CS6Co8TQsV/F64i1nPouV3QmUcCFvY/9Dt7pBGCCvn9a7d
M8KZR/KuqScQmtzHwCAMg/VcJLM/geQWKwQTR9o3yEyWvyxAed4obh113Cyn33rPsGkXc56ZKTVO
qh/Wdvs4p3702xWHip45moRpGH1488x9cQsbia0uYvU0I19Geatv4zqDQ1p6/UwsbN0PF4KAKs0N
qeH44eZ4IEl8bM4o/pYnKyDT7xOCPuWGBmTB5bmjg1Dh30E+5PTVnBGhB5/AML1fuZgP8l8YOb9N
rm/W+XuJq5X5UXUOQt1NkeNv1Pua5kGOQr5DicDcPCkYUh/ls30smvz7L9ShUY2k/KilIisSJepx
uuxQIvbqoXLjGRacyusL/8Bjbubx3N6PLzPRDQ++bhhFtiQObXOWIna+Lt9C9sJDrmYplEPlkpe2
slz61/An3yI8HKhkhbtDO2Uw5fQmLrD0nnDaxFR/jPdNK14XjDDOuP6Bj8ej18AIqfjLGGaCMf93
lprIb+ZMX0qxU+71fY1UCRXOsf5OZfJpeMvGJGIytJgt2rmsEuTt6VxSQpZQXjaSbzLfTKFG5KQS
UNXyf9Gst0TDk33yV0nJHOiFR8y7eNLPuZ0ujz0d0XmiJDl+IkzJqMHc7eucRBg3VgqAChMwpTZs
Wvscey1q6tmCFUX2Dvlt9FUZB4jAq1Vfrv4Dh7rb1m4+6hEEA5RmMB41u0Ssh1bX47H/0M3R7nvF
NBeNIA0OsDAehoEUU0SkwU8Scgxlcz07jTS/nSXk5ja15B82vRkmKHuUhDaRlv6VsbsBJ4DfFf6U
Rt21gnGj1CUz8SYzr+ErOlRS/dNhh24oV5YnpCGe7Vj2MkuCLxSwIV2yP5q71UP67/98c2xXU8zC
FW5vCa1Rb3PBeDJrKMpGsbArvVwx3QuidapqDhlGJVDASaeQPXeUhmRW/zkPTGKFF2CZASog3Fm3
/mfIir7NmQD2oGjb/TKcRWJO1Oi8oodYxhdNo9/vM3qEDiRC+et+xgfxx7kOdlyM/Wzn8u/w+8Yd
IAzFaknMt/BCUBQoSFgeGdtLBUbQJr4B5X3aAyEzHMBtZTL4ZovC5jAhN8auOpm67djRFBs86uRt
3oe3fDV0jhhz//kWbLnTg9NdDZEBsqehc2ZtzYGY+86AyFqW5KRv2BgGKZtetCfurBRYKleJWNJr
KdeR33sj/pxunBa9jILy4CfI8/ZWZDcyXeylDDOa/rRU0XCdfg7DIq7Gif/rKkndVl+mzLpNj1eV
pZePfsoYFJYgx/JFEPFJW1oA3n2gxSbTGvy4WhjRfJiHh4Ag661NtPyGyd5ZmL7DbmGV8D5FsVXg
WDDDrQ9dFtED4IAR1LneeCBPQ1i2MmOA+qF2+aywXWOKJQGWpwyoZtuJGGE0H/IliddHYYhmxYkN
ycR6ytU8FisXBHw0s/UM+N9Qs4NqFw5C12nmSZuhtGs9gAH2Y/XtM1e3/GyhqXm4nCQjWPbgFc63
/8lE6JPYeyqlZcRf7tPdCAHKYC/9nqkT1f8+mI4YpFN4I+R2jnT8MCBI5uhV4EQB78NWpOiT8k+t
yUiN6vEiOIQ62ndNueEI18cEr/5InY1k3CGpEr8j4/HhC514ZsV50EmgPWN8YHEsR/fhHJgrKPDJ
/hvT6kxqKjDS9iqF8FSrKGiu8w7SqqHkrP9RV5M3UnmTfTckMkQwzVFHsqK/gUFfJRM3wj4tnn4N
U2wX2qUuySUGqeJ2BWrjiodMk2m5Pw2JuJh6tvnbxeIhFslKZEZUfq+/zmzu/LihgZNq6ZnzQpbY
w7x3+2i51h+aPl3A+eDPmkIon4k3B9/1uQKPqIBhPcY2rXW/2EpvvtjrknaQZuhIFpBZS/3L8a6v
z5Xriz9PlNfGdxOTlL37tqtFhI/UcVYAN8kNH2GB4eGAroclBDqERCM98Q/VdFx6V4vzjb9DVDdL
cTnbt9Ly4xS37SRSeM/9OXamJ7ZsCceLGC54c5FT3EJ98zJ88fzaqbeOAMtUYwnSJSrd4e+MQtzC
MttTscV4Cg49sUjh9x9oOTMfYV1WE6rBc02H/Ah+WPfGuGcQ+pNqzGC/ZfXz5wD5DXPZnhSEP5kR
2adZ+ogLTzHB9sFBdB3P6S1/UW/evVApS5Z4HFMT0V/9gipf3aHaEb7cq/VXulNDzsK2ORanJ5tt
nLPd4Ef2Wo/PQ5nIjBZCs4f/2S5+JM2a1x8oNu6uo6DXFc6hvWq0Q+DAR498Sg1lgnvmu6JziXNK
0f8oZ92qpSFuXwR8K3VfDfzVWjLroD37M2FAGGktaPkJIkd7J+Oxldj9i0KGJxORwurljr4AaYMu
mO8RySkDPEpcvcJm9mKJrHfyzq26Nza/a1CJV30jdBX8N0chLNGZj906gJ2/mQO1R8qQZZFeuHn0
pllveCVlVkr0JoNc+anM6w2koSdqv//nyBUnZ9PlQNOSVFBxhUnF3g8WR4OcOf6YbP15GWHZvvC3
CK3o2X1sk1qdvkMjXLXfShaN73TNsz915nSCkInaW8b/gAPGbyErC4Lze8pHLHZttegFrme93vrF
GF1cPrHqHBQ70KTZLJ6QvLlH3VhwMW+TdhFRpJdw9SIzlkGuM9LlIzTxIm+ce8r8feDP/guUAW7R
s7O965FLrZWD0C4OSNMedD6wy4XTfSHvkJQjfHkSeHkpAdCYbHabymaZoYWV/8SzJcx+Ee0eCIKQ
3AaIUVlhvLMPs1KavkLS3VM+Akka0SsfoDgt6/TjNfLEZjGAjP+O08+lAIiAjUMu0t99Ht8ahYps
53NwpM3+96Baj9FXJo3ascZY+G5pTZlzPR4VQjp5hIKFGLUOHBSDxVftnCQmp9jkDkgESO98zDno
3Nk8KMy39ruvjzSiJ6yKGAG42Zi0PxpxC5YM/kt3C7ow5IiyaEPs/f1gTv3Bxkd473orC5+HIf95
xNr2jqJpv+jtWMUo7mXDciZyaWW+71tSXVDqp9xZH7ronOoI2axO1GmbHWTJba+7UpRJ1sYANeKr
VKoKeqqfFSMmEWk9pbetwhXmAh33AvrRHbfI+TfHmJSJdxmjg2+fnH/fGehtBdw4TErUBFjW38u5
AeKrjaPAlXGUKzStlfQvDNWNNf/JRxJmVncrSNjvkH4DBTeuiUzAoA8kdmDTemreBfOLfD/ehXcJ
bgYVYbM/jQchtQsbwkYT/bkFN9Ctx+sUIS5mEsdqTrby7yj43dEmKtWCh6FzPnEp46dH8Wt0WoOo
dTOIyAQlk2Z0TOC4dp4JhUcrDqIQZBnCeaZYZrTdzN+1w26Zkr5wJgP5h+yzADCp0z3DaWDkUlZH
O/juUw+PmvSbR3g4ONa2M3YFKOXA8OJ/ix+voUmepXjZL2SG/zfp1yt2zqqiwpPA7dFqIcCCD7C8
8PNCvVacqBZ7Eyt3FNZViZ7y30+Suc8vI5iC2+M7vTQbo4VcBQf3eheOTpf0yJAILXoCfol7t9B8
nYyISyFj7SDHd3DDheTk9bnpM/UNeVdYcFVns1RJNakI+bvgPqufsh2SXmkMuR6cfYhWwH20W61f
Y5GB9HJ92CmcHykdWnQjMKOguIdxG58qkZKezH9shRY/LqJEB8dTa8TSyM/xW7h2FLxkVi7dg43F
z0Ma2+tjDfoA7S0a1eh72XJI84WnET48KoVDfJvzClxMPaihG7+E2UbpzpnaTcno78FoHlr6E0vc
wrgP2B/vAQZMJoSBd5ZwxYGidSmQFsDbkVEhThMUnd36tx9BMu1T7X/tcvSrO3IbRnopWHrDyjhA
UBeyidOLmpSZMFqoWi/+QdbfSWK5AVLHPYJDDdKpzkJFv6JdyqdehBm3ZR0uj6rpnWFfX9MGC3t9
fCcCOm2ll4NVWrOuINmW4Tos9lNLaDNZS8C6Av9IwpvZN59S0S7ul6Ya/wwd1EEbhe0z1bX/2qa6
6n3cpjqvXtMEWrv4L22i1yn9aSMEwnz4W3pPbycbamK1DkqlWUQdk+kfMBCuevJnV14V1AMh2cKS
xmQJ5safzr3MDJHDiOzYQacxlSyyAVTqQnZQc9oEj6cjR5Eq1YEq+BXwCDmQQh3crt8XZJpq+vJQ
VeBiqo0KCbUWlJbiwocvznKBzbHP84XwTn3y2QtpDTs44Vqa0nmvcvTLCywsGgz4n9WebehxmKJ/
YYDw/33aP38FAzubawBBX1qCPc9nHeqXUl8PuwldUwJTFVtAh0kIE8heuI8aMxOT4W1hCR/ecSfV
rzJ2R8k6JvfqkogXOYwrS55MkNJZA38IMIhD62rgiFLpaghmS1KxjoFKUh/xzfbVsRSNpYCFPNmw
V+hx0+VA92vdDlgKv4cw/rrv91uggi46941z4QAu3v+qpWRam7Gb1xfYxyxHPSRh6pfMpqu4vkid
q1wIvhoLCrwgu8c/sAyUmPdlSTsCfflyqr9Gg9pFC5InHClKnUCotJ8CWIbznbFptUlQPpDOnpj0
H+83UyPbrkaT/n6c8hciUyJa8TMR0u60Uur6C7R3/fU5ywwqAoP4SGeRlEkJ0eI6DOy06qD4MiZ2
4XUk+YMaEC1SXidwrtO+0cDb79UjTHTyOpqUTJWlGimgvZ7QkVYEDzRsRc10eRgkybX04EnXi9Kw
anHEDW1MzqWndkQdfM/kgBZXlzlWvPNjfjoKcHTWobslzzpbuu7ce1UfD4RCW/JXz96NKt/BuHO6
u5wkxRKwh+oYq3i3R4qGhb/nDyxSsgY0EXDN6jmO4fbJf7jMLoSwq4orNXvtMTrTYoJM0rihOnIy
098p436qMvsvHOpokYeL+jDyX0ui0IBMD+aIC0fcHM5aETSA8SBdBp5j0XOPUynjo4gCwKQxVtBG
B5W+Rg5eNT2FCT8IW+bqGw9GFcYviFJjtbXxHCBC0PJUifNqmTD9sewI+3OK1Y3JYSd4MlCbdLwq
0Y9w4InTGu63LyJBsnGNdAoczNDSzn9Kdy7P0ovabf9acu0pIqDjioKVcw/l3OwUYVn0f0mFGSQ8
plmbhPC3NRFhatvpygZHUH2oxJZMwCKSY8AAAAvAIdeoKMuI13Voav0k5uryKhUHMWBfcZLF1tc0
7EfMdQ+5XL4FFZ+suzq9w4xTAcgICWviBABoL/Wq4Xk6eWc56QlL9bZT4E+xajlIQGODNj1QZQMK
PEwuSMXSmvBm28y+dX9XmxDtYQAYDxeeffKtiFsFyQD5ZSmOumAh0FFHKXW+IgCI2wkWqahkRjcb
LIlggFYVUDdBndUXqRuZlhGH0rZpNAPd6Z55P9oTMkqg+yy6uSDoDmT7CjWHwBsoiI8HYc1CSTEa
31k3VzseyQCrds65J0irgdkA1LuiskAVn8smBFGDAkOVdwKY80HWBkk+cM7smheIRhV046yZQ397
gJUJF7zK5SFc9WGu/lCl4cjBUyk7f4M46/3Hg+NmrKDsSEhO9YJbOFPfUcJhOYkPTKK1gSUTU1Xr
qQEIcNzHinHNtQG67vqfuWii1Ss1YxDgcsvyLO19wTLAm4hMLXLLTpAMgV1K59nf/atXUTnslMV8
RxwMh5HdSkwM5havUwiv0cd19D9cTvGrkxKCZ2PIcRglNHucsriSMnyEDiO7dhfOFR8Gdkpyz1+Z
sJ9H/xZpmlt0t6uFCjJ1jTAmpA3Nb8g3ryEvu9XQNei+kr04h57FxELR8aXuDVdQxLkIXVB7Gh2X
Jw/B0CaZmsMSUC4gXaMCbh9hg8t5yQO0oDbbw2UndFTvirEO6zy0jNp/e43iexxS1lWvKJ2aLq2A
XtOiw8G3JZOy7qy3rr4F7/Be4MfDIk0g/8Nd3FZOLsqEGuMcar3ZPskl90ONH0QbjaP/d3MapQ6e
NGOoV5Y0LRrB7k50oKR9OpNUW/lpqGpkdS6xb5TRYQVFDVpdE4CM+gn3Ltn+nIIe64w0YkBCTo8Q
0MlI/X3dNmAaCT4m6qUumBCymZMVzhmlzCCjvhs0w451QOJ/BS9lRXNx8UI+xwlol5SDS2+eftVX
EhOj6unUT2ioaQgN2WLhgUtl+vEjlUURYkNnH/OVrN/x8GNA+S15mK61ysfrXOKOpRKANkH4oAYR
2lfC3GeT9GMlIhCgDALiUnZyjl1chU3NqKEPvgT/sgNFEUE5YLyKs5+lUXf519VPVqLxjKSIEUV9
rWP21hq6vj9nLbvWwtHWOzahVw4DuB04x6CpjwTSw3HnOWN2exj81bv5/iQXbrvOMZePuNi0DpUZ
ID7PwDwW7YM78ZAqy8l/QChL2H1tLSL1E1mJ11GMa2wjzjXLcPx+XLZSsKlJQOf/atLA6LsZzhxG
3UeC1KLf3QjWG0ypdfQiW4Nj8s7BR2IqISPt0lpRR7g+kgbhxEDIJK1PGxmcZYQuxOyizHxHv/th
iePE3cjS3Tob2wGrNCjRt4k0aJg/625HhOj1zTzvNPwpiT3ZBOeUwNa6fgLoq6SGymP+NURAvr2V
xzy2ijfAR98S7ohU4ltF2WpY9AWlm4bst4nyVXiH64rK6/ZNA29hQd+u4Xu+YucXkWHTyyLz+s0C
WS7DUe0CFlvuqqe6zPOj3XUibt9q5gFMPqnnT8RT5aSqoGtvJw+2knvUjRZTVDZ8pKv3+4MnrKZu
Oul8qvh+LIqphNvDjtKkGkPohVvmSu5qR1S1kNkTokh+JoyiqL4Yqi747lQ6J74xhp+9NiRx381P
CFtyWoL+T0MnQ4SdiAI7Q8ylwWFKyxcx12y0m+JaGEPoRSoWYvk7RHMwbqoxeauaHcjCXa+kenUI
jtpCCCd8DmGj94tDFbnvVxT7GXPwFy7MX/nP1s5Rln/tVv1+TcYt4ZNLEG9fYWI/5gVo10E7Z9ge
WcQCE78uF3EMNi1K40BUteWjpi71UubFg5tj6IoYQ+J/4x9CwXRApW/t3omUDHf+U3sau8DQDwhm
A5OYO/mVodpeVVgIv66OS2gTNrWBilvTMRCO6RlfC/T69Am6CFrftBdsdZcJ10nD2g1WEZpCnU1Q
hQRSpXVbaQ1vSWZsWVnMR21tcUSbBahwRlnF+jkKL+0YH6jgRMe24cHJRcDyhr2nfLreGIHmVYpO
Wv6VASbwh0zGZjfOqtNTS1TRGPrR3mdleB+TkXyQEptKP22vvq02t2MO4mZW81Hiu+5K5sh/X4gu
eNbVosnyKvsjUGjIP1utLLjXKrJwt2UAuJaFHMLGPEn/0JwcEqMyeYNNkNtpqD5bjRCmD14qsMW4
+42uD/g5T2aNH5rGPZ+q/F6gk0uTc5/YDO1NsslAlj7eDzg/y/iffTQDE8MZhBcFBNs2Q68UVCoF
irRHXUScavaIp/DC0L3f0UZlJYJpZlHn8d/AoOJSaoQuNxHPtkTGnwnI+hxBp06H7Iu06xXJNlId
pQolSFvls9M6RKfDEv0eeaVV9CZa6TCMPLhE0NCNJlADrMHD0+Mdu3NPHx4rHy/oODl8xOg2Tx+0
4cI38mkL0imWwxmRO2XLFcYbdl3AsqTbUNtyvzkzb4neNwo6ZVPLxyPT0hITh5vRXcm2a1285tSc
wlfSjhuFnLMHC7LEB2QNmYB5Qn76ti6h/A6jIe1v7pRXaarQc94QM79nOQEVOINP2Il1kbzCWX2j
NY8+ptJOfYoGQsQBw0sq2FyTwHw/aKWFVpEqcNBkWPCrH5kE7d3026xUuarxgvZZ6mmo3nf3oUsx
CP+jEhRhBxwvNu6PaEZmPEriSIzsaxQ7udWNa9WHodZgIM805aMpaOl28UjJYRXMRO95X3AVJfim
d4JRSic9fZosM7JCGssKDfQ45cOc4WDvsHrlfv3Sc8o9pYT0liv++Yr8P2wBDpnoqNXIoF513QtN
1f4ctGx2DruZNOoOD3sV8gFKhNjOYFLBsBBPkjzbrxdSb5j+keC3fs2DWxVQhdas6VWZJBRKCDr6
pfk0y9uPGqUzRhUomNEmreO22UpNIXgRgnzU0GXyE+IFT2GxPYWgA1XPiOS38V19tfjO3750RkTi
/1GLnwUQDfog/YfM6+kFwMBnDd7hxAqNO+Q2ag1sFR4tFRSo05aCc8VDM2AkNZ5ZCY/DQmsf5Gj9
aNHoYYWbC6OniD5QhyBPOyRdts80RsKN9yGyqY4Linpl6NrfIsDjv05jAfTZgYJL33zrnecHcWV4
CQEUrcpY/HuRjlgAkk3d2x3bvP+H9jS1m87DARB0vfm+481fHdc/3iJr9NzdH1laCN3pVx7ZCpom
kQGQzvtzlclRjflXQCK1gyBn/Og/0yDdpLnBHDr2/rph+l6GMmil426PE3bEDVc6H91M6SDukLUK
tYH9My2sKsqTo8/V4ZHEXxsWG23fpcDkkbyyKmIfBrBuHHQzSNT2cxHeTcZdepNZdN8h37mjvh1f
tv49F0meEH5hcWiJXWPsWrbnGSZ3tnqrs0pnKwtKHKj+ZVYdlNeIHzonQ0c7FFcpgCT+27ejUipK
+48wGBHC3HxTJ2fd2SZccq0TQjJ6cRe9Yr1ozeqSe3eRovDKVic/SbqzjCd43KSg4WyKuktzguJs
faXmJjI87w27SJIs68d/j2C9bVPcCvDcMMWim2AYoW2Zn8it6RQ/Eq4WX2sOMPYNxjX78e4jzQ+k
eD/ohOZeqfGFrSfP/zMZOVBgzgJYQR4pUW9ta7zDoJD8y+6kt7LvYfd39marGYCO1xok02h+IU76
X6URNPM9zxZBO2Agy7tH73EylFYHyOcQx/nNEYuGeJm/O6RZ6tZxbD4uBp2JNfbA6ri69eL5tmkd
uCB7jWDEB+LF4qRopEMNGNQYpzXucXi1f2zDhjqvHUmSRvyFatIYdJIHMNJhddsDhaJzNyVCCQnS
kdNeJOsLAFyLG80F7oPBdUgo+AxLcK+In6GUAxNe3iQyX9NZCm2R+JG6eJqwU6u4FaCfpPvwuOpX
pw9nSXzl+BbUKyykjWa2ZC80XDdkSfgU/oU/JdINeE7mmB6bu+R41tOeP8vvqeUtwC1iQMI6msoA
iU5sjrFA5sR2WGCqjokWQTXi1f9cjCrUS+EL70CdeZiZ01QReQpl8QrqVooZ+gmAUGW2jXFv0ljC
fkzYNmvhjqAXrmyvDy/FJzBmb7sUDQC8BcXQYHOZ+7+hPiPQocmzHwvPdnh4rrzhd9+Sbyzj/j2p
ub4V6Eg0UVNTePi3YSoeRYCzskYaX+oUX+lSTlA+JG9DZ20GczROZxr9EHdqOhUd+8Nj20e/3van
zfbA08xNaOzaTEN9j3YzAGK3NfEPyhDUngIUYw1HjsJrtzX/DBU4N+TiNpr2vvHEdedbQVNz6zik
fg5rgR/M76aqmqkbKNxARUDP3INtlKYox+yqFkM3ss0lN2k3xGDkppkcNEUwKum563pMRa1Dh+ZD
tH1CqAdDNq/0erNpapPqmdTn+K9H7c4h8n0rO7g0nekq4AVFC5cI/TGd0TjI6ajryzVtqauw85Lh
fXB5ZzYFNmP10rLPtmyHUVWm2sj9AsJ26XvnugX8Mi3X4/k2EvIWgSAVF8bAbvDHnrzvoC3S0B5U
tvOnQi9t8Y4BuoKf+x+me1MDuBq/hUzrAQMR2bWGYT8ry3kiLFiJf//UI1mIME1e/hPUi8VSFhkD
1R3D0wwJ7mwMlCFnrCrCBbwNkbRl/H/Z9WDaae6Xa7xCPq42DANhYhdFPOgytcTMg5XeoS1ZYgOD
1W1CZdtys2Vvmv27FBkgepaVUX76BUhqjO1QP/hmuqyE9tiEfjJ/TPS+GqwqungWABuV2JCex0tA
WbgGkcL19VaH4CzsIWYYMI1FhUEOnWUl16t3Tee9+KM7cF1MhVJLgcOEnbOYTGf37xwnTCSIwqY+
fziJOxEjyTSO8ylePoeKVvHEgQzv88x4ZGAKGfgz9JtWG+JGEVEqLKRV3gg346FKZQKfGL+bIS4n
hMKbtE7tSd2mpq4nj5qHa50Fbn5GpE3CIShD2tOvT/WqQ94od5zxmgt6a40cRLCNIK6lH5qfYCIg
wV0SC3vOONrgEXbPbeZn9YveofqO98YdNuBYxhzBZ6Qya3GmXjQiy+oq/qibXlpouscx7/yIaBBH
iLuBGmySjRhV/DCqXGBAYs+K6Snkkd+JLktOJQfvyIRW2o5XkpRnUuwQD/Iho9t3aOvAWc9nx+Ex
VQe9iYaKqTCE5ZAN9vA46fenNT4Yp2f9I9Cc4t+FylNsoyMFXH35PGtAWhsheNXOfF9fFAub7kO3
4UednKBC525OmNT/JbciLKESjXl25nbYQliAkbWpwURKlMdlLeJ3zKAeOWDC1zSV5N0zA9jMSH9X
UCQJpqOsVlfguMEZNIdm2dukXRN3grbkQLhSVZk86OgszoCzoEquecWxoY6g5rNXEr0UNUdtThXw
hiOZxc8pmyxAfbq8dIYz3MS9ZyrGY3TtBwMQEXWMtLKKyy5cjU+x1/rvzTf9HXybER9iZaQc0r0x
xukR/yE1J2cFxjwyCHFJ7BWifHWVcDMZJ0Yv3qXegSkCt7W9CdSeklwGeuGmzSxKMi+qP+n/vmg9
Xcn3mS9DB1WOYrc/vmAAE1iG3J+90BEySTiQEevA2wCPRoVUX1pbyPTzNQWJhkxMtdXrXoehZ54D
7SIO/LFLnFOcX9kTTTkru3wlrtinSdyd3ojJvEXF4CVRpdzl6Z50xVskt71qwvKaHr+ROio5nLTZ
mqXHSPjWrLUmBzwKGrA96vsFGx5/cyEW6bJ1pkSvnem14WCqomhyn5IyZAlszIUopmUukAAuN7xg
3+Ao6K3gBFQj8nqyAiuZ16g+QVuMiUoKFJvBk6ljs5o52SCX4qlII47/5Acv3n5+3wPECI6Kb72c
gdPnrTEIHB2ATKKNprWFQpygU5YP3PXMb/xI/ajdAxzovknbcvooG0toRRxQiXjywdokpR5Is/vm
9mw0bSSR46EBxGcmHVFXSOLC33iIo1SvbwzGgqOcPXpR9kdZT7bWoS2w2kmlnFlb+DR7YjY7mvaw
5xv2uARy+JBUNJZKKdNjqqpdTVYJ3kwWBxjwh4FHldHRnzlQARVMTk/127nSoRudFwSLG28e3qs3
8eaUJhohePPVB3WgX1dsUR4h9MZrBrHZVEWTpmSagSgzjDcTLG5Q7xKPs9AD8XN8FhlpjiupwhBV
8yAlGKGpFDf82u5XoGHG4LCLLlaGjLVWOm6SnRdPBEmuGCfAHpxD2xoXE9ZouPcPQyfu9SA8o0a7
0m+vQsn7QAqDcIFTLQ7znNypTWZmkJq880jHpIiZ/Pcr06J3bfZ9WgTedz0i/Ens/nCivM3zR1PZ
qjRDP0zBDD8+wnr3DajG2Amizh3YMbw6+Pr9Cl2uDl5pGE1+8WpUEwcNtWmwSAma7Dl36AoK2krd
m+sK6xd6jQjFvOdoBAkHAULrjeDCQFSS+8PZMI2qkcoZG1vBDQ7YQIo7dBYxmL1kPMGO+8oRl352
jrPUA+RJqW0K56QILPRVU6QCJVtGnAW9bod30oWQymBwQJjsUi+Ls9RMHtqGppIZ8jmL18JyJqW5
smpB23ehkM1JjMg1hU5kvU2hD0tYM+NvoBuHcI9th/JHFqmRa1kZrR7WsjAY7diNI9L93vrI1WYT
QqdyB2lPprh7sbE8ezCtSILWbRVPBOuRxa0U7mXxynkki/tdQJrRX2bTmuaTNEb09wgQKxe6uwT+
1Acx2c2pfi+3LOHvuEnAV5E2Zz8fDRF11aVASqPxURUo+p4SgRSw7EY0Ib9CBgdxp4d89ObjNRBE
vKM6XGWELDCR+tRIsFds7G/GMCqri3V2jmsTdSafFUyVM8/pFj0/fPtlNo+7/aEtW8Sr8yCrtYlH
JjQdl2yJv4T1B75hOP3YjDq9QN+xG4RF1OCrLCO6AWSetVDTXtkiIPt32jcczx1b87rxh4qz9/oG
tI5VloePRDdCn6PWKMuhfG9+ZFe+tawOVbvangoBT2vFG3ZQN7M4vYNM4gCddj/WLrYvMYoLqhg/
WcJGJbleS2n5dZEA5NCGnScZ/MqATWM3GPQFnM0rBDrZ0DmYRlNcM+DDMZqI5XEF4wpLkm/MqSMK
8EiN4BpuTQAeRy4CuQTz7FIg4Co5ZU6DVlM+IcdT8dKxx9sspVdbA1mX/ZjyOGjfVwwQMO4/QhVH
9wbAESwXogMJ557Xw26W8ZtdVsrpcFvtju85XAlVKelbSHI9FYi6oLo08GI+3HVyXIl/SyUp6LZW
MPJWdwFZ93UaBIDLvgNATuJkjiIehfdBln8s8iNlcdoGWJtZEPHrpz6cshnnPt6rozglcgGXMy10
7+dsooexSVLBKkWTFe5c2kwR8zwSLz31qtu0yYL2gnkuHMON6I1Esu71U4EzinfBEH0Kdryh5ErD
BNmjwa4DU6kg9+Qt92RePwlkHXFVwxPR7ja53lEqUFCHUrVA/S4vgsCgIEURMPOgpenNwLK7j6E9
8kw7gqDYDe7dJlijGqD2RBPMb0+eKa0SuRKVSdYNrhOFKXxorVKBCgm6f5g69gKGRyIAcG2mXjJR
HIJ2qY7G6KCSUXbaAEN3t4x7QpSnyD9BRM/WGW8f4mnXdeHfN1SgEKx2FR1ZrFc8OJho2ZGAEc6E
UAMU4qR4Ha+2XalLln5y2e5kxql53+WnCHkuOO5Cgw9XghnKDf7bhyiCcqf8ervh5uMJM34I5Muk
NPitPuZhwCmfZYRfzUF8ZwNuFxANs87amP8lOf+br3YTQeL9cdHVyVurzRjXb6FspwVlNaRsMQZO
idCivcQL/beC9T1xN3wOrMR255DHT8a+aN9wQaVWo/6ID1dbi/RZKxmH7xGveoCNVs6KyVVdjUzu
iLHucHvZqNecZwRiU/6f6WK+yjr5Zye1Gz7J2vp8e/FkjsI47eOwRUz/T6KKjBGNTN/DPHVefV64
QrzyiUgBGBONDUyXW39LK2blHo0wwKVXS0DU9nsWoX53kuACW2i/4BuxP7HdjFv84zkvQeR/ftno
Kc/Ki9Wa3ZaqZTRtqK1rPHSLXjffd5iAf9bswksqiL+38hq9dkOr2kp9SiTdBgvk181JRYj+jVEh
vlvPtmKISHSnBFJSLtCGjX+ghnPOBXAZlgAyapzA8ICM3XXBaXqGw8CZpBxTQys0iJF7ocsXFN7G
oJXm8CHjZKbYHP3XtVOjr2cu4mNDRTOh8KChr0yUmi9c8AIIc7OROujuoIC8eaUZjJT/DV/09CxI
gYsUS+wOL2zGPFgezUn+c2detXeD/YH2HogcuPccyGGjqs+C8KCZVk52LxXghYYDC2ESM3jxDWRn
MUOP4POPPyI0wRCx/zfS9XQx+p8gZS4xxKpjb+/ykR76PBzJDZhfD1pIGCWO9gWU9qkVdpLbIkKY
jvDu9o/PA3qyGQgjvs+a1xA7gTGFUa6fzDv1+3fhvdWGo8Q9rFfFvYRh+e9EnU8/DTo5Artd9SXf
xpDvgLtA9uY6BZTjTXNMyuiF3p295gN7jBAbG/H2L5E7CJw+F/sB8VMkv1c4PgMW81c3n3MGuOsZ
VKBZgXMoBmur3ump3yK21LNWG6FFaSSZ0C4sHQyJ6vq5eDvw9eV4F3P7KOtnkfGQx1xD6JBeyj8O
CbxlASnh3pHWikZRVmNt92WC5fP9mmTI7aMusb0GzHE8IHk06bqPZGmiI2s6KVXqaz7cSE2hXLoX
cgIyPZNHuptbCssAfExu3K2Rn4sRi44txye+LFlVzHJrmcPTeMx4pesPBgRVgVSs4d9kMgbx1MnX
Nc2aqdWXYIYfQ3nXvF1r4A76DWVLG+lsPIYexD9TmdNHVL2DYsrm/5qzay2WSMeCI5Bzvo24YYyu
z4TC2pU4NiwLsIATqDWeazHI+F1Pu+U89bzWrdVa1sBVUqpl2083Z89wgwgitpkCi8gS/n4thke2
GZfQ3PgMbPe8X4LJcgM2Lm4jgbp9d4zzl+K/xsaeq4MK8BPELroT5R3x9z9FkMdfVFa2F/Q0a3bc
VVD/UncBRo+d5I4wMBm3rJzlSx2bzS/Go7cBk99xu5e4A5NXjbsyxHHQZ7tBZ1bPI5R3LdZdQ5xc
JTeGB3VCbBBxlki/aYZwgEI952a5mX8w7lY021VF1kbyeuVW5D/83JlvjZlEodmhFhpPl3zPNYSa
sv3cx8nkxYVUMikElqPGLcKAbe5xfdwCGTYtdK2lEHfSeapPDiwpJ9G2BFVQMEschTnai60v2Xob
NEbgDJPx/OQiZtAqJCK3uOMf+0Z7Qx+pl8n2dbZgS7yvKrLGYTKqwBRz0H4+jgqKIII1HWW7mRBM
6zWmfIgu/JbcRhQ8yoQ0VqsXC9YUFy/XRyRtKr1b87WvVK2zeASih22cOSJYIjNdkcnIdkB8JaqN
xCOR+klpiscprx60JIYKNHT36hxZZcRkLX6RdDTEVQ0cv7NtYnDZhZe/XNK5pqigiBE68WCnzUV2
b1HHzexm0UT2wLBSVq6ICOp0itvZaxI0pbxyoXz172PQim0d9IHACMZxu0gu9Es1xD4WatUIxZ1k
VDpSNF9DDw+V7egY/Kzn0UVGS1jQnU0KvvG2GII28M/MdQQm0hkOErGSmaBeG++h0KcMbjfMsuhL
JAYoet+E1Cdd/r0HC3CvbAWyUqbO0SHXDIT6lSz8rDp7AdiNuLpsuSqpdZzMSwFpCHlOaxgJH2Dw
iZaSWx6+0Ia51Jy2C9BEnzMQAuhQ1ABi5rXGknpWw+OlXOyICFOpC0g+bvh4EXhWJOEZ8BM24BhV
4y5V9o+GkgIYG8bQLJun0rwXaRsIIwHGpJHHFcwkHs0hbnv9sJUPNYViSR+G4W7NFtcQjZaVxsDF
t5gjkKKQ3y97APd44YKRVq5rG4pwqFx2oTSgQGRhAvS6EeWAHLwG1sCD2d0/j7bCuJnWMuwy/pUd
/wo13L9l4JR1bgtrR7kTTcRnO2zVi60S/wLNuyA9JXFUf8PyNaGjk+KoLt2E6OZ62Hfq1Id9FzhQ
ZfAd6bIRr7Wqjasa908ntPTqVf6Vi9nfZoivkp/AbxtfPX+GEIYfqTD1hj2qVfxAS/D/dUQtDzEl
ZiRhRVigOlF52nBQEpSBsyIP7BpnYCrwyw+CX2vL0Kmji7EUPaIjRbjLhncT+yQgdhUwCjIN6flq
CRl78E4T4ndBn2oimn8pwdB/XG3/A1vDxSc3PfrzbPeFDbdnk8C4HkATeBi9kNORO0CHb9U5d/Nj
IYiX//bRlqhfchW8FoxUBPW7W4f0Sn2CVfBswv9uLpE611KIuwtp284SFrpvtHtAc30KcGHbOrC/
CW1HCBfewP+np/oZu9ZnaGNQYrwx8KXypFDQXwo08Z9VfqF6DSmTP5GRZBk6wz/1CVIE3nQBAc5C
wZ6tKm9i0qTlDjV2lZ1EioiRnVJmgtGDeZgo37lJ7uck4zZDRSDWB54zmEWwcKAb4Ui4Ky0Gfax1
O7Pux8FJlgJpFNVuXaHdip6CqInAFgQvoqX3I2kEMqrxnBY081awkBxJ+xbaC2p92NQx1Pcf52Rc
3iEQIQkBcjAD6TG4LDeggFtZ7u5rb201fgNGOFX60w7iuHw93AfRQqzycENCvVLrwncuaeVih6T4
hfCM3vL/wacQV/sAkUTQy09Mtt0qKFMiLBxkzLd27yYV9CRJb0klWZbEsBZo44WpKyRgFD+d+kJ6
eALUbevBIFsQyCqxBqX3hn5J965QqYesssVbUxJ8TZk4G+uz4CXyk68f3rHBR++VMb0BjM1V/YXc
CdKjvjWHm7QjwOwZqujHjpurqW1ICpQmWQH1i4QQRV477LiC3UtTb10XCvJlkw1saQdHJivKyv46
fIdwu+uHRucqQAk8sk/xtePB/9Mvt0Yx4rItIU90Csf6sllwOVNpKN+tUnDc7U8nY5duKunRfvTc
TWDgJsdcQBlyHEngId9tQYWDBC1ey7RHzfUEDQJMF3Dbbzw1YLcLICoKU3Dubw7HCEHiJoQT/oL2
2Vt0dYzIwTjlwmqzfxsHJNexU9tjyi58QPcDuX5fLn6yvea1jw9iTXarD8vq1P0VS/EQugo0oOSz
wh336m8QMkMcRRXdhIRxafUknQiRf152f9Itnm96/BMutaw8jMq7h8WwZB67LvpE4Vi8FAMMx+KT
/rt5ZxUjExS0nb8sZz+ed4I11DKI2z3y4LRBkXQruo7i/+EV9CxZATXYavH3fucavLGmsPR2QTfs
J5GWSKpsXw1GTtqHF+q1DyJLkWjB0S0HZWP9BsT0iXwsFLkLAvX5QPVWiEO21zi0uvhmfuOqHYhB
1N/1qIzQHR3nhywb+njhd2OLjP7otiAHSene+Ltv4BYbMH1ik044ln9ilDVYS1R7c0CKf3XOANA8
v0PcYcZl6U2Sldf3xYaruXX93O9xHqcdcTJB/Y1ZHO/1T8g9t3E1ipA7WawmHQb9z+E+HOg3ndj0
3hNOEvE1cxUXmpR5TnoBv9gGGVNeluIlAfd5rPC3ttU+IbqS1EJqiCfDjwBMrUX9atzi66SaguBs
4s4U1kEd2WBXGd1sG5/cAuqZbvPaGD8NRIgqi4TmNYK4HuLKZujBjskFLf01txcxwLXWPZICBC0E
hqet8em3GkuSMQkMCEahSMmFUSK3lWm5mRqX0CcNb3kErkbu3KXhWpVgAvSxluYs8jG1d1Rmwma5
yF4FyYdhVEqvh+nN73VAM5Q/ITyYAAl8TNlG6yvSf3E24Uy0LJKoAuSCFN/KsIB7gCVJJPQ42RGm
94pzHySdugGSdjhe5z+OZrzSU1GJiYD4eDiJeptgETJO7kw8GaNpQSQ/j1S2JsuRAzxVzJCOCZ00
gttMFH0nEPxkspZPDePCiNv1gtM8SNs1LfyuJV3ZUXaRygRTcp59zKCmANJGF0fBdwy7mZo5/jGv
I3zMrLWiQCGg2j/a81xqGAsNY5pWxzRuAYKyDCZTdOmKbWMREJsCL4YC1nFTrfhYmH3zXbSyvrfU
amno34z4lpniqfDpr+CGlnPclBIqyFDLNB/umU86pE/YuDHAYpZUOk8d03SVSOwV2LW+8c9R0Neu
qBrdTr7gDvoWbhspugEpL7wMhXZBxH5fqJvNLDBDgNbqJp/sQZTT28rr68DXsOKmMo0M3YYi4fCT
ktNeBuGCC8KhMIKMy5IeqKXjP1OYLnqJAOe/a8bnNiIS4huhZn1TgjpBIrh/DXv/cREfE9xi3ttK
74Whvr46SmFyz2U+2FVVwb9KZV15CMxTeg5nhSA2PJ8MvW78gSS+gie1HJVOBMRC/U7ngZnb3PL9
mXarJNcRwkSYqhLrLY67tn955DgU14BFxEPoRZ5LEcgAeaBXqqUZKHHTrQGztIh7hV5YwjQ3dedu
+XcVVQggRWsk6vZhAU2DM/tmmQAXse0DSKikEqxlAhnyEjkScL//6KfcgYAiF8o1ONoHcqImOBdH
/13dUT6s6JijO4LCGx9lsvGI2JCVND74LSU7SbZi7k277yKB1i9Ux896T/g45HrzDZ3YGC+zPOq2
SOCuA8TJglw+/bH17JK5fJM78rlRWQ9CnVVlw339V3HFKOV8PvzWauZ6nVZqC82bOStEgX8JBNqh
EqJKhngG0ddKEkv2nxeFdGosAZHTaOikAL36w4cqenWdcvuP27/36OU6/uPql6Fea0YInz1qxO16
cQYm1WKYFAFazX31TnteZ3HbdtnSCyPrir0XdEO0fbK6hsd907JwNd5mOPO6hNaiYmbfFXcq+m+u
T94MyzXJ24jyg3mzdOtesxHMFL4WCr72wpoum9CyQ8Z0nRNiL2pSSULIIuaFlYe+6TVlP6d26Ccj
p/SQVNwvkODLUKxQCT4JMXNQw7f2fWvE6FnFDOJPCYC92NRh/i92KyuPWXVyAHxRV3dY3B9Bf2Bq
4dY2hF2Xvd/4JAs2ZgqtIuUQ0v63xwRVf6Gj26i9GEpog1nj2AHcPFsFm4/ISbkOxu0fBQ2Ezz0p
sfHMhqS6AA2wGekGBXNW6Wj3mdPoVtIZE8M5Pb5a2OXFAKlcYh4Zh6MIVvkm42nug+SUhSSfT7cP
/wU9GHUuJdUkb4onnOlUSFH9yWNpAMLyDVma4AscSIcbYV+k6fs5+SAPaF7qaZpOhv5UJGjwdjOA
PnvCkVhLlBvwb3FzsUmYH6fXITgzJDgjibmgE5QawPGb3loJ79kWZUkWs+n0uLL1s0u1r1krR/Yw
2BQ0cbLcV62rnd1TuSuGPE8K+OKYr4wBF2D7tDL7dOBLSOdSTq+zrc9FVLMvAhM8OOA4n7FoLNPP
kG20df9LRiaAiZYFZ1mfKGnRj3p5iFaH9mBVNo+gZnnL0kppEe1MUPcZceunrVGsZyajnrJFVCd8
6MdWhpJ50GmetNiQHXJvvS+SCexwPc+W55QJ4JjEJauxKXhDoPs0Uf5xWPFw8OCwZWIxtdLnGyNM
f5Fhyg1YXJjCTGbMCWTmLgFgcxWUYeQrxDiOTi93nFj3jKYyxMV4lW9lp5x0eQHcJFNJhILQYQjP
mhaI7YOIBgDw2zoya+bW766YesDBzrdI7/5noxLOmbXxsF2gCQnnOwowHyRuoRRXnsUcn8CqSgtB
d4HeC6EptydIlBjkqyHhNkQBlQRxL/pbbUxaKRmFGXcjWFkA3aWeInoHyEe3ErdBPr5/mO6pMElo
IAK2CrgC7CYctY2ArYkP8+HvYUpySSPmw8P2FtyRPxL3MBhMkGxbFAd+gcFmfh4vO7GfcbIJw3eO
rNSTyBR0DOMwvKUqkCFMvSISQ/Qpkf5Px07DZatb9eWXHYACSpd7pXZICMU+Baxn7s5UnOTEXeZt
KLpTtr6m4ylgt9RGYg3Za4clh5bSMtBdQ7eyz0Zdlx8TEUzQqbcDNr6m1Vo8YCFjYApJ1OMi9wHu
DzwrgNbWmd/ac/lxyD0q1G2TlBtDmaDPGI7dA+a1op8ilIBXM0GuqxEnpqOInQ3SZBDSsxHx2haw
ybmHZ/Dsfm1lmwqqrpphprvUXufsaQKDx1fv0Pwp8vTpbWBsCGVaca5BmCJUSprvDnp93g+Mk+7P
dp1Dwcu0pdrKmuOKKqRdmgQk9raOhlVwySmNM9gXNz5qr/s21P4D3f2D2WZcaUBuPRquG5qzgwTM
lh4KKu2j1GSt0s6er/UBp7WCBKvG4ll6hIDUb+Z8LdnrlxEJf7l2BPdGDbmqmLv6qGCqbISKkH+T
GifY+ZEctDLPBLHJ/WWZ08zr5Jni6vGFcuZSxAOG/hWgbs6qbfugakEBseJVOLpBFjHIFLh3J8i+
ljyG1Wfcl+QKoYREkGPbLDhh/A3DLDnIH1QVZpngzh+c0f4m4wwEKOfGWhm27xDf7B1CLdRjQOpx
Z1j6sUTmcF+vETOCyKBLnZqcgH7Q3A3H90y/ZzbdGE9/OGh3AaQVkOVn6xUq1QyQwNu+CMbK+C1g
vzcDPI5cNyeGdilNI8k9GGgAdlhsuzNuXed879ntDjIGylv8MLC7zc4pr5xCZNoiEQqkbKoRggjF
v+d+QyRgkRzRL1lzYvHnm2oinHmP6hi8PbYx5aJI0mm92HzCUzSQpu/eJRZCJtwXazbnDmc1ptUI
fMHjgHofHEJGs3eY9lC+X43bENn3NYYzdye5ruL5WQaNFHmuIpch9qAE7V/HS6yN8laYaFHG6+Mt
snw5POpuACLWDj6F80K+EX+5KK/EF0bdJMusY2Kk18tDJLPnCOr2hFKracvrU4B0EGVJIXoxr9lS
Bf6+NToWEv4S2dVcPJSm5sXEUfOVZtBRX3KFTkxTSqf+2dDvbzfZvL8BWabOxSSlLZnCLxFT7QA2
TbOUwz3+zOu3iOCUlhaHnw9WdVRUnjo14AJPO+T0dqG72T0bSWGBp9R8JsYre4KQVhPcrMHCKYLl
1eHgubJ7jmVh6Sz2Pbusu+kMsXJdzzt5XkfTHLto+rGq/WPEDgCFzWwGCsyCIV8LRbHZx5x1n+hd
KgblYjWtUmMMyK/KSCGd++u5F4cKenQ6bUl81x7SijzvRBlZ5FMcAs3qVVQ/ptoqNmlPmFv9pfgO
pdQyS4ZAZ65g5eQ8bkEY+XxPxIngceunbcZcl3ibXLU9fsZQGDMjp6INl+DFS4W/Z7RUBv8NfAMl
qEfqmpAcPNtv9b3n9CuMZuspOFeiYPljooJ0ZAxCRPHIuBBoB4T7A/GgW/Ab/mmbk4jZ4MuNzDbk
zf3nqKlyk+Vbs/9R5xmgAhRglthAIYsmcY7sHN1k7QoV15qYA/Lan22zscNe1epvAKX9pb5M7zGi
yuyVyuHR/TB5/LHgZbn33WCfwvDYgm+lNdyirV1S7z9zNclDF2Ch7uigKVx7K5e7CmVLSzKSIWuN
3BHlJzvR7JgJJ6HebQ23Mrq3yD7A7/4kaX3pBwAglCxtgf6cuIJQ20Y/kDMc4VKTylGfgYRYyYN5
a/ar+ioZHap2MXpxtXPMsqA/Re/mfFNb1cKuRXDfzGOgCNLiE9rNFeN6EsGz5QEJvRJt75k3Pr/L
lHs2Qw5SgTSyM4NscOMPDJ8Fz7fb7X8yW+4aJdcL375MZFhi7wOAEB6rTYG2DGP+8no3wFpFrEC1
8rbkuuRqT/R9TTf6rjYyS9rhQ2pZY8t4NcTJ0MgEkNqd4unU31im3mRPCkw0d7QFz1FHwpv/qpsH
F2N/6MXqO5lzluqP4qjneYzsYAxzZE9hGSIlI/PxcfYc0U2ZZZw3Mx2HrGrbV+mp929iYVpVYfWy
fPyRbqJTIemN5/n9jpP/HLsHy5uf2IXMdnGELe4dLTdA49YTFPX2tupGtfjNzM0ejo6Njh23PEzO
tRyLoDzKvoVSz0iL/VPBqr4a0/FZr3u+WDdFSUcgOoPuBlAxpVppGoOS+Zjs/cIZ6epH7jEPlvvD
PXh55p2yKdA6boMTPYuT+hiUpyXL8X5DCvuGXzgvM4xetHZir69Wx3aFG3Xs2N6KB1GwNU1Nm0uv
tOdDhMO34slM2/QQlxafPuMwL1XJczf9HKVKx08aua/j8acPWswvZ1ch/+AROwcUOmsDhROmZFM2
SfsjseZhrNUFW6c3Wt9VGUwn4IRC5wbiTd0xrKIxlEK7Sg8pJBQz6ur798b6mcYiJFViMTqyzQUI
9dJ4NLpvtKejsV4qJIzebgHficV+kGF9kPnCmb1kV2pMO6CLN0qZeo5mVcnyKND48dRoiXBtgeOQ
xYYFuQ1MCnWyL7V6r9cpi0w6rqjHTI6KY3N9EUIiq6xWsgz+HFSoR1hQxjmbjyFQhmjim0oao3qV
+zNqjGk9LbSTHtXKBzUmpbyt2UuohuW3cfUq2WjeR3aMPgo8bjTQSbXCcu6C5fFjKXcvRfsyw50j
RaI857aI5vhcuCihdFkOn2HGaUh4BRATElTasu/xU3NMx8ArZOVs89G2cOK21xM7Y/GclEZOUABX
Fd94Fb1OMYd1ia2o50IeFnyK7VqEB3+2vSP8TAPKp408u263om9hUB3l1BMJqc6tJOYbt1+YpPe9
dGtF4oc4a0XlcRGtEwmX9Vn44Uj8R1CTgBKmT3zDWfcn40V9KSFk+kCGgcjzF4UXlxw30gpQonbK
fWD//8xYiGoVemUVyz1bYOVoz2+qqw8TDnoalcbGpx4cERrvGiNG3Eb8Si0+lXmYAf7t7H52lKvC
5JhFAXfOS8mPwsajy+CjZ6x1tnt9SHQXUvseCfeZW0K062tQdiOBORPdTYUP9OBDd3gKdgoiWbm+
7NGaCj/A3FjblZ0NQFQakUuD079XhSjagmG8hj+rL8Zj4WTlxL6SW1EtcKiRdl8uQg8SsjiB+vBU
RV4vNhlN+eHggdloV7krKYNc6XyYmb+3PekvOmOQCin7v0mzBmh51snOdQMH5AlL0TZZlmYteDEg
zFyOhRrLNlLr5jtvR/oHTgd8AbYG7iIw/3GAi4sWOaMQJvaXPS0WJYBfBWMPNJE3swZV3nsQkqE0
MvmWIjpu7CYhqQIabf/UOO8gRsZ9ZHKatYedqZzeN1+NtjAE6SBicCd9WqJWWwg0deN1s+h2G6MG
y8XY/Y/TfjI8EEOiFXNTnJCHIiNs3gQLH2fce0XpOjYNbrwkMNmfhgcZyxmGTLRNOuPSQ6z+wQKv
wel53Dp8ovIMheH1JCulrDIN3C9L8BDe8JhH5Sg5HsMd7WuNXHa7UyoNV90/+CRhLgqPncGqFiir
J+9OH1NHOZeX2rtCYjupjEvGb2E2MYXYlrR6qG7TmAXTmKuJIsydMIjEyPVH8e9TyWg86zB5G/+C
vL16w5FM5At/f3DPoeA+HTZaHqLO1nYcSUbxWI5ZCtHAop+1rfBs6nj7MhZ/VkisWpq7E+Qc37d/
LMlqmPvvNTKenkDzzlreB7fOifgA/3V7DvZkdcWKLsmVkn0kXV7xL83fay36vvPQ/KkxqUGa47E6
O35I+xIE6GRRVgmg3fkMKRUQdRyN3kSG/GmRNCEtxe4fvjcYflYXoOWEnR4sTSOT2MdWwxhXPBhn
5E8Nq+0lNqS1Ntp0pEhfAPmOQGRNETwuGpTddLLm9KmU5LloNSGQUnh70fB3F8I7X9YA2aVEWLXd
F/BrmKJN3DXBJFpI59eqPYTXH9PDsUjKekksbwhuWwW4YpI0stJhQ4dbKEpSMP4N8AvSImDGRe3D
3WiLx9465xsp9wOGk+ETzj9NB0ycVEkL2qHYgbkHp6+qZF/3c9Na0Pzv8sqocDU6FAI8Mp/w01IN
H+MG2W3rtEYkrfAJMkYiU0Pk/bP1CYiOE5/x3+mloAsgSsftpQz2RYYSk+9KNOyDHgeA8SQrV3dz
IeXUlzDMbR1C+1+6wB9lrdhXKwDerLgEioWJbwXxnTXHjc+2IfB87LAZ4kykCbMH1PkrD/MmTr8g
RtJRXn+duY+M2pYraUofxQz7XURIDeFbCE0RMXHuig/F+zxiVYHjgi7u2rG1m0OhgUVZcUOxzGe8
k1ScSgsq0HBPqRX0paKi/lui6SJ6SF8H5tfMmYAqIJxH8Cu5IHS8lq/gqjcurRPUYWtul0ATtGDS
fAyjwTSx1vawYP8DFOOXQcBNkcsKgiDVrmdvbBCp1JnrQhk72lF/cum5bRxpJk3ZLCHwPUcuYCig
PIs2ixMD4x7SaXntUGdFGsS6NDGKxEMLDaqJrKX4QFdCayVuWJhcSjgSTW6mv1k0Ebf8U7hGrB6P
gsVKNZq0oEZQlMl6p4bkBRdj298P5hmKF3a7g4bgk/CADALHuUrze5AbWgoyJ1mWWIvqR/lC2Oox
qtofObGrUfZGRb0+jejQ41dvARroT1cEU93uL4F4PTmgKfnDW4U+FaR80D/gY3ZmFfHJhliGGzzE
9kM7lPmEH3PmCWM2xkJeKQP9uxN/4lBo+1DOKjI0Tgl8W1+66yJSNwzx6Rjt8hIxP4bEsfbU6A+U
C0oFnBmmARAdpsdTo9R7F89xng22SN4C+RTaF1RwNxlX9r+pgInQf+ogXxYilpu4+11k5yqOtsNJ
5N6zfn4S2icY4f76vRPTFOy61PM7UW/t1tgdJUwvYwFe/UK7ZnXhJB9oGb1mioYeXt5C0cIVOReN
KmqLogVmN81sY1ZeXttAAjP4pJ3XKoeTnakwKBdxz14m63SitfiwUHfCPHRe1x2k1eLQAus3uUvM
DpacLuy15g2/zR5z9Y1mlpNy7UgKbxxhTSDybSJKokodwKHUqykN7VCmFDsSLuuLKt7k1EpCJSIM
9MOrc9eZNjDC2ZB50ZNS7ybue/Vo2TdRwrQbxCxiDcjOtqeZc9W5csKBKmjXYci92bSo/sJ0p5de
hAAnbZxadYOPnLk7vzeAKyJuhpcLTVOm1RE/6cGsJiOjqzXYApr0FqoPjRNC1w6tQd4YvCFe58YT
HQ8df8Aj9lXvOw9WsRoRWv72rIRDnV+9hW1NSrxy/0rOH+u1w7B29TvnUkmRPy56im9t8rH8i7H6
fvEqds1WjtUxEU1LD54JnaL5goWkpDfR8v40ZhUnrmcJGrIK7ERkNSPvL6RnA8rv8jZg6slQpvwm
liKFP7CENfaDjoWF5EQ8qdu4RU4bgPN7gHb/F3cYPZEFdDLzRMykOatAbpVNMzsbIC0Ul/yyvbVC
Zts7LwypUITpN8b0B9FubkWIDbZsr0hIChoEfDqSu/YvnH6s1UuSupCR9SLqbUEyofJBzJP/gfEf
IHURr0vsvGLgMyQDrebVJBfTZUdXSAMnsaO2RUei0fOgIhFmmfOWGJBEpNvxAuzrD1JoKs2wb+rn
5tUnK1ZuoeHf0tma1H7UeZXjh87hGIS3NXY5XbSxVMu1UgdsrLt4j5ZStD8pfweDEWJP7hAgMhf9
pNa+3S3AwmHZ2LNfqv2+EigNN1mURRxDBjiUMR6Or03G22Ahpd2zNfkLTpgW0/cJSiS0APQuQJFQ
3w8Y0DwLlw3o7hwujIaC9WwHWjwZQ92Zljq/RSsQvovV65Xcf/+NY0VNPM3+T6YOa2jxO9A0BU0L
4wMkBTDFskSoDwYrL5XNlr7zSqkFeH30TBqQwmVgsDT3ZyZ2DOvgePQIxjimrHlHDispAILzpMpP
zCJRtjxWZrNpE93YrYKG3ZDHb6qIxB2F4GcTEKeI+uD+fj803MoZXvN4+SryyFBxkBx3uz+zI2/O
AgFFW6lT393c4fPTosJvGusPgDKsBZLOtJgoJ6yY6Ytr/X5FefTClvw7sPWokg2mwUoRyrf27Yt/
uUm1rmd5SrdDM+aMIOhG535DLGxazIerYlFhxYEkwTTED4goYvh43q+4L9VqtpsSrHfWEF8zmRZV
YeZepIkwI8D1BFpf6k7O569/uwPbUposxSXMQGCFDUf6FbW+gvU+Hlh9BmfwVPBXiECeWhfBVNN1
58Yl1yJdJ++XWrO3/oqK9A4F4/m0yCl3sOFEFH0uANgdoYAt+zcVWgCioopJGL3RhnyHkj+dLzuT
EHnu8TgV1+Df6UBlWC7pvfEgy37zN3LtiOtSG473bAz2UiBjlcmwJp8ZMeBGKOl0eJUyfgscx11t
stTdetiXuJhx2k2y0+rcS8jiL1C4mOeGMRCMF5uiJsHC/Y8COnLLHMS4xqagflFZipNYkQhEs2qY
G6O4bdR9MFl8VvTkbd3VmsGzbT26UUacIKWtbUvRt9gBsc0nV73Wex03pmzJqGVgxeE0R6AWgQlf
xoXCSMsoOlbZVDg5lMrpbAGZ0qgtxx9sLNeev40ES+EeOnuUcIoKtZ8T6v2lFotvjENNJl3rBS/A
5GCopAVhvwSFdDE0KNSd9ah0OAdJYfQUp792J8iUjf1WNeTL1bB+w/I9S8VUZqabnoXk0xuKZnrb
7/nsvQVbbpYwsWoRbMmHm9EYVmKG8vrwADbKk88oc/vYgchGyhoibqlLOd18VCaiZ3kV22PLAR5C
QaBFhQf7rtQwvXIRpTwOuP5M2mfVsw858vpzsAHTHo/k9g1hjUEcNuydWYG8KmdmhLCPPdR4Zs0n
XzRHo0gw1Fh46sn0KUQiMax+2vjNgD7kXl1FpFcKbLCMFXCNm39897AeInnhBRXMaIbmp1F7qL5j
oH1AtgCsTHu0iJ8kz9X7vVe8EPyGCdx2/aU5PW67OsJApLUbxzfyamz+AQuZ90gjccUCqJ5p/LFl
7WO77SRbBNipqdbEaTMMAZS2yGJPaUJc4LgH/kXFp3fOKPQ98PODYPmIRBIQKbTC3e0PX5yWQhA4
fjtxWzFt8iVYJIEOM4hvuwihCNj2L6LheEH5YqRpUC3igkS4oGftycL3kZUbw6N1s7W8Y1wD3glt
VSJkvekeSBBCDdf8XkZhCmDXaTc947uWdsIl9xzvC7yWFbanqW/+VlShqqzqL1nJe+h06gv5rwEP
rT/U89gHWEiXCBmSdpeXhJFEu/ggAXCO0CJyJT7XvjCa2zxmyYGrDsRptMifRSa2cy4ifzcB4JoP
VSqjWeWtIgBceqVGQQaSTPgEgMCJtA8cj5suj9B3VJnf9Np6zvy/rQcCnJgbw8bZ72V1UGBdDOZL
sSyTEcH34lQCIYLvfBlpTK2ruiQwSE1/RbE8bPZI9mHhw/j8wCJW7EWpbRlfNlX249dDJgdEflz0
NgKctUI4u2EsunL9mdNWV+aTAp/OrMW6Prx7UJ5bBvGvf65rcUnJpnhdN6uz5alOGWb4kJyNbKe+
qh/AXih2IpiOjNLn6NANVAsfYOFmheqpt+yjSc+h6qUOWzqS7pKuATZhaAK63zwcNv+Da9jpIXi+
lu++bVaw1+1EIrfwhy5EPAVZzd3ZtWdo6uQHNwKKc2wpFC5aR5+gTo1JfR/ssilak2UKs4t9ODAn
kQkoH5NyGLyFe9D8uB4ALma6sSG9y0qu/JXwyJ7TSinmPM0Nj6p+jQSQIXUtrsPkJdPptfksMbgb
LfGz71z+Z8xgyng2nNDvj8A1kn8UB87sSkt7mLb/O7DbY8AZHuv4N6WZd0vLSWvo67mMlCfu96Kr
4yQmz/q9wnZMU8ZMRwqPMFULe9P9iSy0ZrWiMcy4QWmyqPPuN3OXkQ2pDS640lpEWjj/RGPt8Qbt
piTKsdPCeqnPyQUvvBOnZkVxWbAfBfCcfYbgCFA5Rdv+0F5sihocnqONegMq3/h5nsyaRfQ6KoHP
5MbTIBV3i7vFKh9opYHdZg9p4LyyMXJqqnPUEwhc68uyIbXEGrcDrbuGCiMuQdPzn3+BF1nPds3x
AOFrkqO7IXNfq7663lIl+4gxwi8lspcJhrSAlKf8wDgPImZBBGN1tiEFDd0QQRyzfekb3ejeMW3A
XAMNNB8sYSHW0XtC9DawGzN+ZxQ7ZyKAIh3vu+cp57vt4PxPRDzGNJ59CgcG1YtCJFmyOKpMbvlM
XJTbFYNpwtWnhTxjU1LTpZSFJoMQKSsGxRSXUip8ss6RrsgZcQf4HVLdqxI4FkKWVF3J951vazYM
nH2G40zkLeJJ9y6Wa5T+pPvC3A4n54OrPExY58cpuRlFuhIAAducoVnvmzT3SxW2zVcgjUWkfWHj
ANYLAbA0pNWjObhHseOUFhiyFDd9rlcHitQItKtvxOaQLTV34u1zHQOmePlN7IF/Jin7zQKH3JvD
sNtO8m1OC7pl+HeMTlJbhdb8ylZLZvUBVWqU//sCIEYHER05imdlNc0ImNhV05foe7jmzzpJnlax
wH6JHhiNBkk5I7iMMZTOzchkfGaFTk4/Ai7MZcLL2VSLwDNFa0VCVdUyujTRmNLL5wehJR4DuApZ
x3p92Zxl7tJwVdjHUhVqOjM4PjG2KmQpC/+yrkoOTXXmYm1tOFAhlXVH3e4f/Qk0nMdjULPd3Mi7
DTh2coVKdTyVZJQ/4VL8owjHbEry3dM6Fzhrjnf2P1DXSnh3IwFDI97G1AgQGG+3iMA1aaLMTpih
ft2eNyvHgnYySifDnhQR6wHfiER83Q+DAzOCAiR8bK8J/4HJeaLP5KqBkIOzh5u7pl2UWHR4Igvx
d0GMhJwPc219Q33i2jM784v0NZGfpmdbUUSb4pIWpEjkfT6kP+566y+3mLH+w5AMwjho+R4Vtrba
ynh+fOXMOzSaduE5frK3YnxOOEuNgIWMQaLquThfmsrzmTyJRyocz+7hpZXXwoBkceoABsUORo8C
YRqAERe9LZMHubGI5sen8NymyGOhJbwfrI4R0+idYYj30hHpCtAApy8qMzXsuYGvhpNuKHqNRzlY
VkWoEzGS5TTS5TFW/mbTobAFOn5gj9ZYz8Aq0yOE8xwvdzAc5BsXGTeXOZTXTc0HaX2ccPEtrwIQ
PQktMGCP/isy/OKRIs1wqrKpH6OLeucb/wCU6zL7M0Uatn6fuYT52z4RFaGk538zhVldqEbmBKZc
x4MGepRutBHVkC39d7FebJOj+uHd8PA89a2aMPflutRx12z4h0SPyLomoHKXGp5h8wD/wqtlRA5d
uMYO2/dpuKitUxQPOpo7Qki9Zxcy+Tf3JDkvolvMlmPbo85GmwuMRUOmFN/sA6/3QWlmKuMqpUSG
aP0S6pN/vGy5RsDEX3jYc3jyClg0GPzZUkVpLKAOyA/3lJxrZuRMzd+Ne+a/HY06AYpFNfLrTOYy
YGxOLPTTpfPKurYC3u3Sq2GXVJnlYjC4Xt29ZeCQwDFuxTMOGOgy4NovKj1seYi/sw/eSkJDear0
wzqaXPTfndAYIo6HLvnZQmIUjwk4CpKDZdGS015CCtIwysXaTlg5SJEirqoBeYvkqYeYS18TJ3bg
mrJsnWvv8sEz8s2D34ZLSI4eAptyZCua/NhtCgiBH8eOnSQrmacnF+EqsTIsYvW9B16OpD4hTa4U
huokgHboVgMQp0bn/T1h+DDUDR3LxE8WrUDr0BOoal+OJ20Uk8QPD23BCs1gSmagytXOw5rIffJb
Odmm7aXiDrK5tS1tRe5AcJWD1zg/jCBEkkitXhmKAASLTVrGeE372Nj4LWIVUQyajVsU6aEhN0CG
8twzzHqRQ0Ve5Qlg64VAq3Mo1qvRPPbO7u06sJH8JKPzJ7y6ff2VKnMILocaSoZCek95VFIzAhcB
vC23yTp0dmrysGtWoPH2Ghv0xs/LByFxcZYXDVx1QyOED2SDBjbMIlhXcbkIM7ejl6BEYusF+h7f
qleynzyGLcrCHaKCdQ10wR7+ZP0BbIQsA3bCuiR4R+pz8woF/92B2CKCWvpGXsoejgR/qZ6/2Vr/
xMi5zxkGc+omO/VfzxT+eckpo9xS8WwgcgdQVtYRjGytDyufd/Mo38ZxrvsD4pUeDjsgDbdbTNhm
ULRExEX5q3h8mFuyfs/mZ3hk0OWmLvSFOBIz7d/YzA7PvvvEJy/Vw7DeIzoGivk2oeFkQABE2tCm
ioVrfRgoIpL+8Q2e9CBHLx1hmqjbbIjWKnuJ/E2dvHvK1bj4zqMivi3yPQgqdCCra0JM5RnDPB7I
3bhDI2uISWVfinm/UvqP9P3GwSH+mSnlRNneBmEc56D6fRZ85hOU7XysWOOizUOtp1cpwXqkN4lV
62GfEYA/R+MNatuUpSIXPm2SoCnJAj7OYNOuUr6bEVhCiYrHMkt7MWzIIy1AUOQIrdGKnSZHQqj6
awF8fM27Pw4HwxtgFU34X3jrKRf4O6nKIBWVo4k2unUqQGID14xBBvc6J//Cbif438vp14AdETY2
lUXppXR5E8CrLrH1vjT2WnulFASMqcbEtBL+M5jjnejYcYV76BW9VSJ0GZuYXRvEXPlCLBn+ErFc
6YmoZBO2yvpwB0oY0AxaPHeTHXl+QgpzoTlCFxON2BJRk4fnwQGQqy4uDoDY57+iEb1pFWX73S35
NpBvGY2hVIUWTKOYVeO+XYIp1iR/k8boXjf2uEini2U8MnmGpDNk8V/1k5NyWbD6DYeq78AYj1b2
cgRv0XNzis27FGU4bH1kKIh+5GyKLRotnDeymV3vnFR88nbUz8B+Ypf1FSvADm9xq21yDzcnU3TS
Pt7RYZOfwm41nurMEhRW7Vi4VpOjNPurlLJfdjPj1pRWOB/gDBBBDQN4cw7EJ9aR4r34MOqKWwaj
0feaoTcMOyISO/CTaUfvTu4ECQbUc4JHspOPSG8zPAqCSNlGkXzRMI9wj3V4vEa3abgjZH3WT7a+
4ta8SBN9YZcE5rMJQibpep6oMsQRLkDQ/YeXhRUemtS9TrFuH5JzCVblo8z1Noh5End1/kr8puxS
Cc5Gsw430bn2FffhKGO9CeVLWg8uqxiVeIjdsr2kKQ0trlyzUZKpW/xBEEv2pwFZbXW3KPT8LFO1
8x9AFdfNuewl58AMqLsXP6rmLRZ4AZk80L2m040XNNrzTRy3+mOkrNj1ILdyFxWDRf1dpUr2Q9Ax
Wn1ajHiyEQdONBRw4NZUKEl2dYf0/DVSPa513eepBLnY5UUrMBvdexPa2rxo0eZ0km6Wtzgl/Aej
j8RfhfliVTbLs83h1vW5pOqU03MurvoHdu2MTMOS3cO61hyPrapfEp7fbzxtGvS+9WUisOq3OfX1
2lgshsp4E3s/4YDzAgSZm6Edos4UzH2UVTtENGusBua97d9m9TNPUFNuykXgFFY3HURSUEQ0K27T
XCwMXqrgRpV2nmZHHoV7iIYc5vHslZPS9JDLSHBvpMtY7BmRPvaMXBndQgDMVrpH0MZ3QszxSh+Z
V65vOGV57iv22bTbjhcrwA+aCzrOm+L1ZYEL+yN7Pm8N3SUZPeNWIc2UUpBW624oBxL68+yXG32C
iA+xThla9J9rzezMfWRJHUak384nYZOiQPQf2Vlsl0mh9krQn488arOM563RizYFmMu+mQhJKAl7
V1CJ3s03pS5ALymbcVe2vrYRM/iA7zxouepxfbuSu1r1gmVTGHhB5a60qdPjTjxgP7zPfujqIRaF
/Y0o1kSiRQ/wJe05H7sRg/+plOZcpBoIYj5QTOBDbnyisnHOuOaLTvuUPXxp1R0fRKyLT6ZHJ9tz
AkzO6+jlgqfMThfCx1EnHE1PpTrp/lAYZVju6s5QRXnPv1p94GAaa0pBX31NPpxoLy2w0ipBZZq5
DFp4/UZMtAbHPTZW+XxMgHwqyqF/ipad+BETgBOM6tKlMQhULI/ZA+6Xg9HpYdXBoVH6ySu+6XZJ
hlFRdqXThe5WVBP6CWKM9kJ6ExKIg2kLZMpnofM9LO7Vi+He/867IS2YmIu7Emz6B2URzmPa1qwb
TsFzo4BOF687xRjJpLRRFrESlxA8ZHntmetCIaNYzl6dCLKhN4Yd0dhrEujOgGxrWUiRQURBp8me
9g1o6aDBcpUWXmXU/7jNO/YzDUywbUywHEZmU2hk+JWSzua9fhTfVo4IrWZ7Ep9DQ9oD/8CWQQpp
yOs15ToaGf7n+amdIDnCYRVpHwtLzrjdSy18CjOd3sIiN0sOgJWVAAV9W0cV9Qk57hsGeBbdjIX/
Rp8vZGDPyy1ZY0ppMp8mlEBxj2z5cNozgqfs4vnxMqNfpNgoUPis0I5iA+z0NhRqFTasz2SjPPku
T3PWd7QPuzN6EZN3Y+L/9pEe8SqJcXlvSFAnU+oYO5EC9RJ+40nyZ3c4791UqqHyAIjhH9WyreSJ
CXFDC7z+v/uCGbjZ52i7AvKcrTC3bR1PQA89LeJeZv61U5dl6XNMgoaed3G55NhnfXRGzjJi0Aa6
ZFCHSTjLsa0+qbbvM2u/nSKQRVmfpCqoItHNaPtn+ic1JLWARWwvrWqyRrE8Rab68NXmn42HSL+q
buQG/SsWUZc9XcHwyWxSVyu8kGDvUHkRdYvR8ryQ8hbq9QoThoVVMzHvb9PZEnwR+f/CpKKLlp5C
Lwry3NrQragJTVzqLUkKRolrWAo+fvNGNEs6sWgWzy3hk4HV2u3AJKuM1LNjftVIJsVnL6S3hCRF
rxoDiQafddLdDe+lz9OlLUmXojmXtv1OsLabadUv1jVPSM/s+OtrehctCpLw42NpVuccXCnoVlif
ET7ZHf6llG8VB8SvCnQjXwduDS5l+y0cvqQjKKoWnsDPc6I4VHE6et0wzAOxp753guCf45gpXqTv
2iNl3JRal9kyCt0r6O/BTVzvTTwh+MtOzKTwzS5wDrsmnilz7ZCxgrcY6zYCD7S+XJLdnPhz4qa7
1sNSWydCZlUrpK1h+9ggJlFAmfl1/Q3Csd1fpDYyEzBYBH9/Of23Wf88FoDk4i7yuljyde3Wr17K
fKQRxCbWqPNcY6Ec7GVJoLF7ktpJayQuumlQFWH1LfiUWvj1u0APyID3F8mfk2HOzLTkhGgiLiIY
GR7MIT/nIlSrK9xX68fNRc76pdzWQtHB7UHIJ7xLdnq0QTcmf9i+r7M4COCfJO5ScfZhiuO+28ri
BFBcEfdkgDMUGHXlzq9iEWCoSZXkmQVZG1cxr4+3Ai58OXvwCc5iXGNYukKr59fBHs+F3kLyanlH
o0zIXFnb4NYLARZXv1VZdla6U1aBesg1oQsycPzk0bhZaMUAV8L4eIoLsK1pAS0ThmDpzMvEfs1a
AtWQBVsmvNrMXbpYhUwaIa/8nrMw3qteMm9W8fh5wNiRDQfc3P8UtN+bE5DMCtPi8AMDzWmyKtJ7
ZDobdVaU/d9dMYR7nemew0uw9RCs18o41S8cIcMwI2OMqyXAaUNwA4hQv7HKVqyc7UeUL0sp4wJB
leuaBUhcLUSFOO2arMZLyxScbGuOtZ5snDLOUS6B77O4G3srTYyKnAghpUTsFoy/vVkP0v9dBxQ2
m1g1L1W7ngEGdzV3wZ1rNvZuljnRBOdXPwog2ILW7lWSouGI841pgnx1Pl/6ZZHmxw4LD4U7vts1
i5/qqygpD9XcvbXKIW7pEhRazcxkRB3sNAQ4oX5OyucYj/mqz/Ir012JDT8KNpY8WfGzq8/wcAAg
ItwasxbXjZcBqsQCpNtgeOaeqzg0/18Sxy+udl5jdjbQDCNN2MhIhjbDOL0RvaGRjSVLPpDhenig
R7K9VmrUPREhrHhizUUNBgtnzhhNeb+hTUp5Nft141nVxYiH9HUfnP2PkCXAvbY6zOWWzw9p4cLh
QzMWlqHxMO6BbG7Ok+tqNXrS/M+I88lrWEfxUQzrygRV3eA0xFWSpkvfSCrGEVYftKZeik6Jyi6I
NGUHPE0OVVnQ2uFD/vlocn+yAsgJzIMW0xG92UcnZ281wF81TW58Jg8QnX+tqkEK21Eq5kOHmQDK
L/2gCCmMD/e8K6W0K8OQf5rQfqTvQWZrzv8NjGBHno4zdFF3mw5b23fy7uJMJP0P1rafppTVCTML
Rm92+v5w0oEJEmzRwKL8RaOQsI88/ek7qB+Y7AwnskTpI8SfPw80tsFS9Te5pLITdqAm5OjR303S
pfLokUU6ohT6/KkoBLuIRxO/csUyGyIDoWPh/iHe868PZ0XKXVQeFMzAIy10Ci+TdstnVxqLNyk+
iisiFEm7Ran8QjrRb0qoCAYOAct8bI44SJxsMslg6gD6e/LNB7ouGRTlxSpqY7itKtqEJDKdv7xj
DJCMOcqAVjJnEgnno+4SJMLdONud811wrxHkZehefNt0R4X37nGkltcD83IjmVnJIt0hOUOCHgsZ
3+DRZPEric2OvejCPFGgIgnmajWTjimMF/dZksPSIfF4uRa/2jsCytag5AwxRTR3lV7aA9J1JtvW
q+oew2BuWfF6rLq5MS6zilCS9H0qjlPTMzyCX3Ojd6TNZ53Q0nMRn8zqzVlT7yKlvhdjaVVktGPk
8EiKoE+Rpo3olqE398yogHU03MdXMuZ7olUFKGRpCAKHIUAoYgeyhdeBWDvtETw5N0/O8f3Er4ld
7iDrUgOP7W3mebsy8GAoQaVZGOhAmj7bzAFV+9UWLOW89yOHwQZBBdfGVjI1SmdQiF7ciAI/kbYp
pA0R4NkAw7jaRhJ6lZp+kxhhyF+rn7weC8ydf7qkdGeUvH6by4W+27MKgaGKSU0+nyvR2I7P0sFa
umSu+DekQtoeFi90vVCqgIv2PQZjPD6EhvOO2uXIYvw7xwe5aO4H0sxVuYuG9gR1vY1LUvKcmgir
bMSOoN5IpRLklYYFCG48dEIMAyNUWbXC3Z55aU4FfLnOsB5pb4YkjzpKbCMViVmVMb9k/kiiMg12
et7JpSFaiY0j0Ai6BAkmjQhXYt3hHYhygQes9GPGYgOSkSaYIv6z208hMDOsHVtiR8KMHZird7wk
IUYZSmOefA25bFpyUOQzbh4LeLNsIxlOEwIQKGwixarGN11BNG2ZRgA42GnXDQTB9aDz4VoYn6lu
JSYeyh9pCIJmwtLsNGYYfJTvA66ruMavOl5pCt9pKS89xavpl8gMKSjP9V8SGrz5fjjMZztncIp0
2cdPZmzWP2JtNp3Lc9Iv5sX9+E4OXGC9vLG95/PILt81tf0Awge3wG+GkxwcwJkjA3iayU7Je3TL
WA2xm4X8ixgqAqaaNtZdU77FSVg3eCGaia/02bHI2EINB4oZKaKMAGSrPDdK4+JzFXqxsYbU9Z+E
OaTDA0yq8lJ/QT7A+7w0LXEMRa6suKdOL3jgmDVLdQSUJ/3JRMrTS6If6229Wowdm4nadQN6bWkK
vN3rdN6zSiShcPal+Z7wo8wyC7pFIVqiCaas6sMx0y3jyXbf8fcCFoceu1IYdD+MBVOGWszedllW
pePL8H90CB21mMrbyx23z3xkt4MZjg1rET4IZJNH7JuMFodIcf61EWDaCSqTLlKiKbnfeGOlf7Jj
KOkbvTpBUjVitDnWPmzw6MC6vIK+XvFXBSSzqyhZcwbanUOa/rzVN5yCjfZbl0QjVmnVQLjEci7+
MwVEXiVp3l1nFtOMfREQFFAaDicw4ogSaF4VpeZ4IA8rqHCNbwIn0eNSg643ujzIrtZ+q417Dzuo
LZxhv6Tijni9hhXdCsm/QB25GurY4VxIhb4mXTUJIaBo9kGDC9ccpu4QAzh5MGRR7C6H4ERMddM7
qJEJG7cDOJs7mZx6tuweSrSqUf5AJKKK9WLIFTNX5W5oYuQfGUBYyB6LbQFRXZh9WwpH1oQqZkIq
oGPFn1LYczHmb9Dz0dwFQ8qZO20nrBuQ0Bm/Ap/KOCIsDxzrKrwJKh3XxNUA7Cau7rdqtz8HpdU/
Xe3yFzNMb3ca1H+lFjiAyRDc24vNduRhV9qzTUq283uUGi/2lh1aix8sC5YFufLBsELCaE1jYh3H
zEoa7A+/rm7+2c+om3BIsotGtXBd3Eljehrcs3K7xYjQf1RRWGU+LXjIZ7EYiKps5mlN46i1uyAp
5Kqkv/I/L80lkxhfQTuzS9vCWLf64fN01fbhDvZ41YuJZozpRbdByfJFvSHZrPZMu997yM0NSZ5N
ShmT7Jy11oNiaqglfGEA5FHom59XweXYCh38idQvk9kGEgIlvI8S7YKMli5VxSNp6HnJc9Mg/2WN
qj/X0rH6Mrs7SpO/6BliQydVYg9HT3FTNRzjbx3D/3aRyswMEPkr79bMoLxOwmaWfvU/vLP+Ofx1
OUknBQ+NWR1jivtKNlMzC9r/brP2p6m6/JokYTviHh5Je/OpInUKnOOt9fjwIfgCOC4dcJRnmBhB
fZeO/D3joYEskm61KTFVMQ+l8vFDIrq0vboCEECSlUSLTUD81y4pVO3SH9u7j6n0BhaUVxaCEHGX
0VRdQOcjtXOP2M53JpWhuGVcAIMzz7qkLyuCtFj9iP4iCwJ+B+iLSvEeQdIpftHDZc8rI5mmwnOM
owqoGY9yqBdo+CAqzLgp8WgWTWiYaq6u8lE72q3ytqLhptIldmmUfHErVJ1lko1Hed7QpvvCVEEL
lZbj03206mdVxR3iKpJfvx9u3PHW7yH/8zXjmVZk+wVrqPjlRqJB+Oxxinzyeeqoqyq6+ygjtDih
0Dq/vK38dwZBvN6pdQ6yBA89dMyqaqhlIF5LyIpEFIce1/OHANdc7mfGCDbLq4RTyEHPA5ryCnSf
gMg7GZitnNGzipiurhfXVnGAI38Fk+UX7NKUPxs9f/tZqM/3v/z5v+cbdN90IVtZJbWVsAT5AAAt
9irnGX2HT680ZAuQYTfP3DDsOAHJct9rj5Au22r9TbQhLZZ6PHKK38tQavV/ykQqXt48gCpXdDNv
QZWZe50KiV9gV/GWhkhoelfzdxqRLRqDL8OhOIh++gQ9J83VwQnpt+yTaDovTqhfVvlbvgtU+aQ1
TdIYWt37Q1RTu+zBzqH0xToOzvhzAN1cMXlqwl7V6GvJq+iUJO6lvV24Ks6Rs9d/wspyvRAKNE5o
QKTsMBxlMYDaCeyXxVn3QaxIPhF4IqDG5eIGUy8vnaulCyB5wUfqMCYGcAxmksRiUEMK9CP2bglb
5+n1goONtZM+3iJzMvGReQVUbvFwFoUT0uFzN/LkjuxkjHr322mjFxrixgFsQlDByP3nwkdGrBwR
/e24il3zugUCybTXbloQXHTo8y1Mr5ehCpKh1mthKp7deBXw8oJRkmARMv+w3rMZpimr5vCskEJ/
GFLYYvUE+nhPdYmRiVqLeBYg+hXKq/MnWsqTiRvhQubn+eEF+UkK1E730rMleg==
`pragma protect end_protected
