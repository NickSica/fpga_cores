`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11984)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5IQJj49NipZ8M+awYasSTowTJrB6A8rap+B7QTb8RJkWraL5C/GNCvNX
9rQWgF3ovgzhkoDfFcy66YWKBtReBjnZ29WczbXv5G2vbWhEaLN4Pq4Uqg7jP8laSKRalHk8IVki
NBMuUd5YX5sGKhSSAlU194MS5jN7h3eqzodCoF+fUaHc92WWuX1wfSom3x6wAneGsBqFn1OE1FQM
6HsZ3IMBC8S8P29BMvJd7tb0h/1je5mOIyb/D9qF7yxR8WmIVLQQQBqyik0osFwGgiBUgtH8KKdA
scFGDQw1fh0paBxdXTRk2eGdZHvsLJV9oFjb3yJ2M0xDLLmGuMmgeGKWy23VDBtWl8Ak6iHwKoEP
XKZGdvjutAZr6XV4Tsfz6wEd5pynrrXzDbKu5b0twS7qdboQi1vWB7wsgu2LQmmpsnru6Ci1HZLn
eXBfiZm8umsBiKTie9z8AnnZnTU2PzZDQkOKx5GCakaAq3cP9NUnThX1ORrkpmUWc+CYjLsqeFXN
xEpM80/4Lo7BHssVGmnC6+MnKL1kf29C2dwtMMY7wOhHQVDr2IvSX/XDbQBNHOooHG0QDCQMcQzk
Y6AJrYwmr4Lf9+s7mxpI4GnlaBjrhU/792gwwidA5CN1umYpAjy2AytYPwPoreGX9OPUIh7Y7Vfi
vYtfwKm5aMO8SB5Y8iedDNdiuAI7Zbbg25FmLgjsICDwd+kC1Ft8kWgxViULpWJFNgpoRIO+c7/W
bnXFy7NsAs1lRPbWEMbf88DDi/ZmvK08jacrFX6rhnEjItToxXychHhdtWWUjaJkRqSRDkC8msig
FHREirkUPXXQkUrVjDYpd2P60ivqPueeuUlkWA7eFu1u1kWXwFVnkCe7m9u1asUBUr2bV5422stz
cUKtY97H+/bssYXmhcTLR855swtC5XAgug/axGgLiCr2jPptvwLhPZZ05UT0FdwvuboK76m7VIZ/
ijnCP3CU92td8/t9B8t54uFhFgfPGtZ316C++cC31muFeCNqUbmfIWoUefp5XzH4jV8Vzpw4ivBE
DuVpDcLti4VeRakZd5FGtLSwY1WBlX9H/pACR+9eAcp7gSBYbB4GJsonFHAFPbKsPn5JUVDdlt1V
9WbPRY3EpJ0NcxnKP8tQ91xDimFLF2Bc6/GSZadLIFOCoCrhuAWpgci2S8wwB6q4EmspNeBQf2/e
PW+gUJcFgNVTbuGfm7EF4O1asY3EwqO3+xjfFp6NudLLE0WaaJnHaAius0ynuwrE9lYjWQYC6XeP
GOdS3xCSVpDIu6d4F9dAeZ8mF2sNo9DTfenjg5trvw5J+UZwq90Z8EIiJZfDx3sABcw50WdiDsH9
UlPeTJRBdukXcQjcH4Gs5gmg9TX41ekz9a5bb2wpc6cKqhN4ZOJ5WPsw6A5iAqljZU9r8EkTaLNe
ZjmSjmGhIxrX1L+8n8+VNn43PKmAq6g5GwghI0ePH0az7oHWEWP3/AawAaP2P6uNTATZq7dSyAMc
p2nD0zdPsxcACgVixQEFdHutWlaR/+1s9Sfc00h7xFUUH290HSmehkPVG9mHcpL+rkTogzM9umV2
l6yMutjSKeW+YOa0irIz8g7699z+Y7DeDMrwzCsm1KQeV7gJAY5iZnfr5XakkdFfhfZ2dcVGHg67
mgSl2fFsqe7M2ecNzxj9p2pP4WoYEsyuS6jdIz0fzvPmDNljnv7/qi74xxeYasnVmP2RpddJOJsa
74NUByKdYpN5U9c42+LFQ8vPphcReDRYr1dt70rtxvKtohG+/Dv6pOQ8tWM+ZOcfWiaW7oRl+YIf
nFfXwglae3VUfGBvI2cAQnCJcvAkDmB5q4WlGoyd2NUaONg5OWwEAZm8w+KnuryvIGcEf6FPIPcE
pD0W8CX1AHmJ4fWic6P3KP7cvPdWoO+E8O7W9eKPXPMikybf50pI0D7h12k6OWpPqeyb7ss7xFno
y1mpDyT4KoHtLeFYi2aMAhGeXkQpytrSpWTc5qIwzEnHPHlZBbkC3IHYkBZM+GIelvKEHpOIGB3t
v4VEigCbaqghJno8jZ+XHwVhW+PFbNl7Yp3qgxlb/hFPG8aDTpS4d+sar8E35QUDrgEO52Vz9NhU
yUE3usNz0Il9MCtFQDjkiFWrvaTvifnJW3DSgsU7n5fnd4W0ZxwxW8l7gSmGhnRPWbOXljtfibJL
/7DwPTGFgES+BSSzsNYfn1sWLtB9lUmHnN8rxPe16oBPZZrXSGaRkq2weW3yXr7OFf8UXk2bzABv
JUO8dhA51EI+dUpRvA2VL7H3P0NwwtcWJCTfWN1rEYqPS7uZUbRWNwhIldAwrbO5vpItL/ePQ3IH
JiJQUAdsiDw+p1pg2hUNiLJYOkcLPLOSPFiz4IVGAlWFuDSTnsKhqixnLHpEk/3WcRKmZ07g1Gu/
bzd8Cb08uVzM6/Ic9fVUj2ZuLOtLDrHYIK5hQQFVbuKxVpL26Th8vIUpjdZSctKaRNu37KW8o4NE
1PjRzLfyBF6bud2SGBj0YfCr0RXRUa2/kXQLGpRa7k7jEMqh36UVG4/qFb0XxzEkEFl7lJTEJwKb
Nn8CflTRMDMI25CBofGVvN6eWz/9w0cSlIQvB8CxPe+jluQu27B6taQ9vUyUdULh8xS0xzV+Ub6e
O28hoIct/dAe5hPX9ePYZzmmn79eaQWrQSnsdXs/lzGuKIRAWstTS7G57Oa6U7ijSJfNqxB4VJDZ
sYskKPPSTsBtdalnay7Ul3VVP8GXvoTFC8uRwxv/gyTR1wUJwd//BpCrXAHAOrujzbf8TpyLJ3KQ
burvgciBL6RgdfajKrq3fGP2rFK5accNCwknz7gXkdktZbwEpxtidBVBM2XyQgnFXlGG3AAFmFBW
B8TyPArdgZ0RGX2/jVYgBzouXZeLk1rfNrDXWvXUNqm2yx1eh7s7Z0xROnQ1fprD2kAi+YcLtMX+
HvMXOPiHebNfHOvGTTrsoQaz5+qFNulBs/1iJ7O6XbvZdmwW3BBnr8NfvEyymv0DOyln9RjViM3n
I7P4+gOcTxx/lGBgY/uddcPhaVVrX8IymEanCLxvkhqYhtSNpsKPJs+YQ3eRDEzhJboYJ5jb8Jm4
l0RqB5CyACyGuNR7QDNRU60xSi5s8G1TP/r6xGjzvcY5yqARv02ecegZTKmNDYubSHSlVl76iEAi
D8eyTYAY8HReaqUSQcIMJ66N4wf56q26tgEwvylc1Tfwcd2Lx9T+vzuf+LdY0ZAeMgzPkaAEvbSq
HFF9sdSsP+2fxgxFN/p5cIpGTdg+wYajKg1JEoD5+LRjFaA8ERfZGYeWK2a5hPhJrvmpCV3qsar8
LvN24u7mQ1QUaZcHASiH4PX1UO6PCC2KqXnBMR5DJDtNwTPmTSWigXio2Fsr6k7j39sparuchJ4w
wXCD5ECFyObvD5nuEcIQf9AOcfXVuNjvP0+nLMkV6fLVSR1rRL/wMCvr2UoEMd1ePqDpXhujemDo
wwX3FGhB+WEUmzDNSYilmTYPObaAFqrDJS/q1jkifgO9AeHWDzvvPe8XQee2aZ7Y8obrG9juVfrw
IKowfQMRBY1izsSmADurFCrjg+KfLutCqcJ150Os7SaqXLAus8eBOe2IPzudPLk+oagcPBst9Vju
WD1ul9JgTftXeT9O04Dov6iX/7nArqLwkYZYQL9LK2zDnxeRGTTSvdJ0O1JIX9Mwm4lsNsC7nV+U
Tbqy+8hD6HNF73UpQOTRRd84QwKpXYHxonzco9U6dvsOhIrIq005E6sBWAEgsWjq5gKw0ihmiWeW
w8rsrX6mmeA4ichYYOzQUb0MtzrWXdSDK3pCLkS9Z2zkIR5+929WZLKN+QFsR5NrKeHHZEpA3BOd
ZC0xUBh6xiXEyjOQMYrsmHhGMQ8NYs5ukw1p+TsCdPGUhnoV8z3Ij+nLyTZxA6+xmwj/Cqg9ueKW
RE227PZ4J7ZDWnepXO/CyrhxBGnfqZfmy0tAPtuQrzrvkvprYM+WK4PYCph/4jaGxFjMxDWQBf7I
1np25NREXS1oFslkB8fgEK/pBrECvtl4KtEpvpxhHH7gK6PMovHCKft3P3tzpUgMrJHIUUJD31xi
UxICRzofWi32LUfn6uSThZ1T/sk7S9viMxnCPU99BJSSMqVKeSWWCJ3+bFsu0VImMyyuA46uM3+U
UtGtAZG9tmDvZ5WPjtVgxxFsDDkkmxUj1reYKW36O8s5P7pKPYWo9zEQH/XwK53IOjY+Jbz0ShpA
kFT56+zv7uXXN4PderG6JWtzU65YgP++yNmVecHR2rDxkfm7ltEVYRBl98n9TciFGkoeJ+VMcoH6
Yl+qEfMFyfYOM7BPmaQej2hn0dPeAww5MH6RPjUwR0LsXFbUcKNdECAEi+Bw4lcio8DryyKAmFLf
ZVjCOoqOYtKDVubYIH60AszNgILbfljTIDG2Vvnf7GyQYdLgIBmNyLzkouN8cPRRhMzOK6sMsDOg
gm41iR2nlNZbD5tEzMycglqiE57ZR5OgopBy5Gn94HKC9a5/CxhSNdtPrvDvTLHfO0LNl93pGOf7
fnjHc3fbct4cTCEs2mOYWjvVeJ0pREDXO+Pz5Gyt5VftgWT+/Pwq0bUK/Qai996kYRCMAvBTSJ/H
ktpi3n99lPOg8d/t6+udRwXqqCg+yLViAWGL7XS6VeyBL3t/KFWHxFq6o98lZd/PyTuEmvHVZ7PH
2nZdNd8qCTJg4mGGgTtAZ41AR6xMTrhiygrCwFthzp10zTh77v4uSvaxHxGLd97sS5fYte3dVMzm
NzAnNL5MO9M7hTnZ27TFJKEeiABW4b2F6yy+LCMqM6XtdgZ3nUzDNUM3KDAKS6lG3c8AKueVE1lP
9lZ3yiKHkwiTjEIu5AXmi0ck/hUxgzq7QyQ480/p9l30KGmW139A4Ssvp1r/UaW5Mc8XB5POg4JC
kr5Z2d+TQzo9ew7yzXP+tr36wONbfRIWiyj5jD00eMVf6d/HyBZgSjh4930XqMyFxGbs02BYUSkc
3fExFrisRpjOIg8+uzDCND7fT12DxHHucNaC9FLU1ZybSdrfDvsJL6md4bYGrex16UdixCBIsUYb
7hTUaLzfG2f5OsdDRiOHUqusmGvthyECCpKod+Ju7jyuiEtnwBVbtWPh8qPPZT0Qy0CTNxr4Xj6A
vi8086+KQp61JxojxBH7JUMcJDE2db4weIpWy8o950Qf0+xSNhshToKDitoobZLQIKcecxTy517D
lPllGLfgbB6IdOZKQ6KELdxIH6TmcclZjRKxK5Ig2G9QGINsSnw4RGB5nmXKp1XdEEw00dr9Avno
nmYaFfSQ/PBPB5USe11wEB6tgKaJKc1IjxiMKsbmaLT/4CHH+51ppsxbXdnuPXsDxbQqt956yBEm
pgefbE4OHmPQf96C/Gq6Qg/WpE3CoQA8jpCE12taPwyzA4KfFzUrpNUzVkb8xBBwPBsG42epejZd
0YsJcK7m7fLriFNG5YHapogU2LRt1w2gwL/6botIGYv91QEVOAi0wt/N6HxMhPDWOCaGSOCBec8u
XdJypsnFZ21Ij36UYG719O7qR8kbF5wsebRSa4R672LKBSIYKUZG74jY98W1eXDWpGYxcs+94ERm
LkBQ36VvydgBRHZhkwhJG3djfug6llGcN11A02on3PBqPkjh+FrtCxsrkLbXfuyY4G1Z3UvhCDOY
xkgBEkvaVK+hc2KDlEgjcUJ0qTdG6J52+fqBg3refBggf79/+ZWoc1OL3Jbegcx4LBpL9OwK4Wye
KsOLUUy84yVjUWut7obwzXzMHslE/ai76nCFrdYBC4D2E0eWJWpGL1j2erKIT6JsQyNsZCirHMek
QD3j+KVsV4Ma/XlKzIULKSy3Ve6tE7/oRCQ/2c2mHplBLuvxjYesWx8gdc6nVRpgvX5ZmiU1VB6s
wnoO7GV9QWAcSLWrVjCMTIlXWpoInCvG2en4h9JzoVStVOgP33gmmnw9QmxGvGCDR2oLd34jw7LB
Y5WS7K/uzJxMJgTPULyaDiG86QD2Cz5zhUBpwbuDMXw58lpVLgkuvO/JKSmyfrT2FuxqneL/3OXR
wxL+JQvzI4EU+HpE8LbL/NTeFcXsznDAATF8+NP46kh4oN6pTthFd69aO06zD6jXLPdjFqt/DBZl
L13Wht44txy+6KSPG6WanRY6uSqhoYHAsTBG0lzx67NethskDX0ahaN3r2guN1obGpRkxN6MpmRW
BbrvN1gdkQizHAjbv9Z+AzITo5T9rEoc6M12KYs3m2J9iGdy4fjhXAWmZVJDRwZodi+9pC6Si/NO
/fEtET8Pzq1fcb0PPzbD8dksYCPUzJ/t/gkCXkOHoQHn0pkvzG9ioXQd0IpNlDB6f62BLfNwjOSP
0kWDszugwc7xzU6Hz7F3vkOFrLUotXtmB9g7xwborrUrBRwBQRkoESS0waXOsXPVMAGXBdcpZ5nA
FhjHpawnkrZcYjCnCwOixvX98S4K84DnVZC+pa1JT+sDEdvQH6G5jHexdpw73JeKsI5Xc9SlA5xf
93i8RZ0TVHwf86YL3GDsS5p9Nl7zgASaUiDglpUlbAiyhtuKKZX5D4p6UL2AeTtWQsBDF9oSMGDB
6MNGaT1HMCYTpurmtv12gOESoRclaG7r6osuAU4Z1JeyRI0EEabvY1f/Te1KiN+EVgtUT2+97lL/
EKZk2kD5/fOU6/KvqncBGX5H0Z4X3pv7WXlH7iEa3MDmozIwa9iC6+AUK2VJzKUz8jM2AJ3N6tv4
g2lwceeEY0gVtX5S5TwqVAVuVu+wngwCgrH/JUr2sNn1AUHkOFOXvHnqCzQEQvRJU09G8LuvychE
Zj5LC5N7x3LhtHMLgoh0bZLZ7TqH0lQPA6FQgH3oGaJ3A5wbg7YroM+ogt0XU4cVzwBZQ2R1sbkf
9Q4muxc0ttVVK0g25M24UvZS7zoXqa+I0CjcjY+xLz25Eyv15/amBCjWAXk4HtNxqyTTi6A9yJPU
390TWzttVn1ddZXPdzmr2lpuix5rI6hkF8a+5c2fRNjzmXbWhdEBsiTGMVxnrwhb7yJqXnXJMSR2
W/H5FnFuwcbNsHjAQCxoUx/l1Yhe0+QeZ+c7/By9uxKR7gsS+D1K1qqRp6bt3uL9MU+DkJoqZssN
8sv6d798sA3tbsajo8a7g38bSYk4TmjxZjXYyUtJehD3H7BkkzpUGrDvnkGzVhGgpy+v+/B75ZhK
kFhmAOBgO/lTYWSeyLI6lOzthKSjQyFlpCVNbleyZX2cX7cHwH8BnCYGqbWd+2792e8i/8PMRzGS
DyVPHQczIwLV3T/H/+Zzhoe6N2wy5oJkcpTwAcYHhvtV1bv303z9eU1tq7O02I8XV0yqYgc09WM8
zQ+OVtwXFCvdsAjEJfpD/Jk4znGtURm/zyJGwAsNZP0Ym3o4urrx9bJ4KmtvGbLSaesxczifhzWI
ocn3Bzq2trDuRebqiXA32C2/7kMRyeQijr6Frhn0tyEXy2T9cKfCnthIZaN88Js26pJ/CthPanhY
en9PoKCnAHX/uyRX/wILLrcL7w+APgpeQgwJfRt89d/sxljhMgDlf2ztK/OwZFw4hcHx/TJQJtyH
OYZVaW7jAGFTlRTK8oJDplmLXoT8+EXh5KfOtZ/vR+V0FxmWtNVrzVYtbE/RsXVhRWFXbXu2g8E2
oHP7CSuywf1Hrf2JfU18lHpQ4qSjbrV8Fw1RUK4PYRCQnr+u6oR0bifeWIwNv1HVqtsUCq382olI
2FxP6tRcX5KX7o7NEh6WJn/dTuvhVUGCK1oM7rFqxHIott8D6VwB3eGatZbPAPuvdGG98BCNlx50
wu1kOdNN9vNd74n3CbUOeo/jDQHlRVQFqNQ/KoD8G09tm7diSdZZX2hk8mU9NgS+VBnWmjQzkNio
7XMpXa2gBuearStf04NQJKq+w44HmUR/naEECwB2UXYlAvlW70ksESH1+1fHkAhnkqr5EbgbgPCl
iO9KREI/4DNOlrZfIPATtcJLIfkpHoZngZhBdYULiwHU74/M22yWJ0k4RuGPrNFgdRGPW0ba65Aa
OkiU6B7Tlp1x+YUHB9/Dvrl0+2VxApNeGZKIyGusuhFpY2ky97wCQGq5bmeQOqAofX1xjDXup/tH
MleSV/dkZUYTA711cENmrfMnXpnpubNJbHyPDr4L6cyJG6iUjVUPdGIMx6uV07eZSuBB2xBy7k0d
GYON4omhmSYeSFH0kBvgvs8kIIV6zXtnYZjn0oNG3sY533eXmhOh+Yx04JhIrzNwtb/NOTGaJL64
RnLlihx++hixTzKo1Al4B1rS95yqDNm391iZonJ0hW37LC8FrjSu5vkT4YF5YtthfvanaDtNuHuV
JQdTf/uEBTLqrDRJGmuhUjQMVvVEcV9nLyUFmIOtArsj3uvGAS3sMX0yutszqvpOxTtfPPuKqkHA
4HhxRCC1jBXi9tlue5uqZpFtCobegV0qgE+YXhUluLBwSXAaRgldBrVC2V0tOBENkCBQtPbXrD1R
mu3YKzmyGCbIYf01NMH2lrhkz9jrarJPIaeyVMaCxgM25PDRWGQGIwBbrX4YMGZ8z3ZOaCKamOWh
sFexxJDUEusdpSOVVBnRSnLXizsDlB+9mJZE/7j1C5WV3JdspY/Xz73IrXaKh2A9nNV3u//kirSl
IEyjKESmgE2FxRzur5PRw+3hVcdJbmAeX8dacEWGcjbFwOadkdbSdLzQ0hkRe+MnLoWBicmXmhca
T6wxDkSiX83yO5u7F6n8JrcVgJm+3aQrpE4ziXGJR7Jf+0lWtWSDMl1SXRpUzkceo+jqL1PcnuWY
jq5bcRAzHCdhZZRD40HQZchzR4z5riCdDimU8VxEmztL78V76h2Zh8TM+bzbAHOjHzCI3R25E1en
nK1EK4DNfDHM/JHasE4HcWdWdIXiN7hD8PRPblZWUo6FVQjd/YyiFYinrcH6yKmudhyvksrMQ9Rt
Nwn96MlnXeK8n/f9dA4v3U0818sZQtPZo+GeZLoCLP8EPD6Y13O0bF+pr8qlVQ5jp85PJ3M3cl/b
5Tmm5SnRL8dDu9oHRJja4FE5JvFbKUHuGeX2AtvisM/67AFsdeHh8tEW9Vz1GV2WT45oIe9DKpdO
i7NLqEzuVxlZcFRyqZSU94ZDjHIVfGv00gMYnI2h8LOH8QJD0yHdtTU/hHuERzgdqiGKMciPPLkL
JOtObl9EYHPIBxSghSST3lET7R6Y8bWFAN+nNRsisI8fUJ62cbsW6Xl0MrN50KQvdo2qORNWgVwW
DoASFsoJyhKFVPZWfKJw8vVNcI6MKl50kgKfkkuCweJO+BuXK2MZeK8St+WqaAIdGJerKrFSdUmI
FPf9r5aGY6rC1qutcPaV4I6SPGFdZEywvS2EIJmKEOqt/9KSbmBbRmadG8BtZHU+G+6jtIOKhHxm
DMAxZ9LRmjbIIjw6magkgf8Y3ZgfrQQ5gIDEXeHD0D8MGfTjl9MwJ76Fce/Hj9LW2jSwUthYOX0g
VFK+rXW2+e8ncXKwurQmWrsImjnOZZ1HgwAEHy5exXAwnftX/c64iQ3zJk1Zwscw3k+KKAwFPIau
pAAcy1DUPVuF9jIQ5xrvENknQD7uGvhUfANaj7B13n9OnnbY8pDvmcgxSIJbkRonDhp17iD6jgIc
KAO7LBC99GdGdj2Wr4wnWMTYWffBCDURWQNOLYHjspGb7FNbJVQLK3IjKEXJx7fBkKjoEahgO8lS
mBuIv9GUQRcn0r9rDahLyLMznimEjTYZURc7FLW1ypbeUpn6SBDVFGD+d4U58OfsKkiGaCWmpzmO
mraZbWmoH6nmsyzXPxMR0d6nC030LTGMs8fNEB4nRsQJEMYxUJS5Lx2+c3DDIKfXGhJfKffYsz+f
NpT74mg97J2IE82of7tPpxIlQ45T05a9bv9XSVPnNZAbwyscjG9T17V8sUttBiX9Cjav9a4Ws8Pb
PsYQUwFuS2Nh7FOrqlU+bmZhfmDc8EoH6YP7zqjWyRUqk6xfRNEO2HNjhW6wc81Hb/SmnL/DvNil
Af0yhKvns7j8jrhppmH1YO1sEFaorzUJG0dyG02Dr6zYagjPu1QrBajcRfwce/FpopK1KOwUWLhP
IoXbx8eHCzj3IaXguIdabmbuuJYS4LSI1HjAATeDAjjomAfh2dG2oeVFvCaQqoor7MWfpPm3ot7f
jyj6xkEp2m8iEmhI//eBOoHFLvQrMOcss9ulFw1EEnd31sQLBtw7yhkxP14oHkFe71Qzuu7QOG+H
JEnstaV/sdIP+3qSgZgq5W9ABO1pcE+tfR5bTevqxvzuKC7wlKZ6Y+NZh2hiX1oE4ZdhchyEkNHr
1xw3229m2U02eN3ZFSHkn/isbVyRUf3xRS6tMPhrc/uAONlrgubt5qVAYCx/uSrHWmjPLb+QCRgd
V5ckvD+0Um8gfOavX4uDp2qDb/YiR0LpQpCXB+S/uqxBVr+Ln4q28QKOjtArBX4s3XsFy9uha3PP
TyIqiGO9Twwtbcp9hQ1z+ReFbLAcvp+j/ZsPfXZH/feggEuBUzTUY40col8Jer9nxITr5lxygcM6
nq1ZaMOtpHRHVO3ODCZc9svbzrST8NGePDVAKDyrp/WTCDdg7xhtsoC8uAvB7E3JTvXVvo7fKITF
fMDnq3mvpZPPS8gjuOWyJW3lHSUbNHrlzklWzZr0hzWedXWme7ltIy/yHinEM2zI/hqUBqxNORSt
KXXxjwIaATBvpgn+GUrheGhUoVCMXi48sBOShkFQGQ4r4WBnRq4jlvO8WohXrqJUohNaqDzaokJ3
Ea+XjCM930OS6h6Ke2CejKX3mVM7Ob+QL1pIP/AWMbWseyAF5vcIu6y7y597Sf6LVQ/v9zq340yC
bTbMTnhXgh2eoCPg/Lxg3/9KItRkjfKGVERIt5cUA86Jd8IsVnEM0tc0MhEdp2eM3oPL2SnKKQOB
puzPMMaiDt166KrsNQVlUD4inNTBQ9PDGPAeq80wqKFxgMNIOsMva3eRjF88L7TfG/AHZru3TM3y
cKVZKh60LnjTCsDyepptJLjIpgbEnOm0uAzNIvZ7l9FMp6QJecDq72Gti1thRwGWazQaY7ZNzos9
Vw+UPy+C42fnVpwomVmV9UayLwsGoIQHGTC3ojNx1iQO3fG/94F/mZ7ze2hFaLWdTUOg5EtiBizq
ignqT/8cWbabmGYVvXoQQMQKiLayrXjENXy/pbvQT/fEJkMC9j24KBRq5zOl6dHNCm4dGCzCVed6
vDPNl6A1XjYwDP+8HOs7qozqf4zioksri2brQHU9Bog2L4bzZpCb4JDYg9cRnPcSgkNDNaDfr8wy
z5ax6GAif4SsEhUnfS92R32UI1zZ7frtFCuOG0zRoDreCjf6o6rlVF/xTfRydMpnrP9IXfCNUqAI
4Z3Kf4WBSsPdQEJINrgN3f1INl6MJpX94xPDgBZR78zjiMOemGZD+0Mr/9xCR2dVcvvS/CSD9M0o
q/oKj68d2Dq5XY5j17WZ138CB2krZAUfRXuOlaxK5kmhR9VuWq2zUhdm2wd8bZm8kVyGMlD0Yyn2
py0Ce3GnwVB6lvSyWWA5iJGNb2AxoxDuXre9vhxmTxbGBD8DBL5qyTGolDY0z03iB5lDW7a/0DTF
C/7hIJpKixuIbtym3Cr43bpB0b3tU4Om/z27bowezFUleKJRtZfyPYi3ehDEGzRvrcEiCDvn3yIg
B0GDE5cfH25OLvbhT1TjCslJv50wvqNuEzzWTi2MLfHbWjPTobPVy+n3DOYkv5E5+vUD4iJI8Pdf
B2on9hqQv7Sq++CYrFB9i6riKe1MYiiPWjTVmyW1blyK0Qwz9iIwgp/9LCG80qQ2Nyzj8a0RMG1l
NCkCc9SPW9YKRVJI1KJ0pEaaGcB6++8qACgutXxPVIM36w+etL5t0/c+kF2EHj7rZnCF5cB7Qf8+
n8kLr1I+GfPKTKJ7+gNJfVHibYqs7Rr6wFgct+XUW0Svr+Xg3jH1sYat+unToGa6+0W7nEAXIs3I
oifSt8uyyyOzwpI+MQw0Fu2nEOUR6w9AwoMWQoEhIDu6QD4vtYIy4pPSkH1YtQXZ6lnLONSQtYRK
YKjTI9ZfYmf4ETgQ79ymMxdkcTtTJmfI2UIdARYfVGJb8jbEpN+txY9Hyw4/rU1PYGQ2MNGp4ARS
H4kQsjisWdEHbN+WeS0tHkoKt04RxTqArqcJ834jdty7MGcjG9w7BNXYUBGrF39ZWYwJZ101JVfm
6q5PAAt3+71Jfcbv6z64QKAixREx9cy7XkV61VVLGFVnANAN/aIuwXqsqAoH2nNf7f6zUb6Tgf1r
N1JincwruGsGr6PtXP8JG0TB7N227jQ9LwjBgmdbgNGImDDjOY7Bz0x12qOs0rlkJGZkOAjkOv3z
yfs02uwkVNWyb/YiO0y2PkWn6lBCLB2FDw2GjbZ12P0OZDw4GC1t3SuxU4EyuSiF3xje0OD18DEI
LmdA0UtNd/UvVBXLNhdde/wX//mnN8SAv/WUAKamSweq4UEReu/x0XsLrqEIRTy3QFUzts99bOGX
NnVJkug52AuQ5w++jMWJQkTM4+rP4FWgNQyQi03N6/+ZyLBKhar5lewgDINqtmvk+vaEZ62wx7fk
GzIT3AdxK0n6JU7wP5taf8+dfMfcDvkjXmHaeE0fcQCSTiGXUXmbzOWNQFtf4pKGL1RJj3ytsPrV
GhoojprweR4UzyyufxIqVmBESOY4f33RqeMf7iFimdL5kqnNv9hZorw4ylKaAh1peY9D6oT0s7aO
58b5L/5dDdGFYUm09w85m7EMMYICx+14q6i+Nbgnxp4As1RwRVzxXvIR+13VLG8+Iq+qdjz3CPfA
zd1okYNMRclOiK2y8F1km6NbzCgJSWEgoeHFWwtbJDt0MD28kAeXyNkTxQXYalZMz9GSxtcq1OmM
JctoV55kYgpLqZXxQ8m/12YGw+wKKwJwl4y5j9Qi0cK6QigkJA6cb3VIgOVeS6931IA1q3bfZTff
cW+QSUzupBxvzIUkaX2GiBXH4ZT7woXmELZ/8d7PSC1glsONhM01DyVvmlp7PC73FGusleQsOi/4
e/Kg0ZZ2tIzUipj6h73Df8fNl9LXqxjh1EUVREbFU0List6hMuGJEBcogai+FS/w+7A3VmX5qPFA
T8rhbKDzLuuGeNcgbK0TxcLkoG1j3BwM1sK5oP5fsIswb2tSX5sfcfCZBmQei0bG5aBYVWAMDkdF
iy9uQMzvkNe5L+cJ8mlT3R1aTBT5v8ZVu30rccOnVLABHxN9gV82YkxerIGOxNskVIdk4FYls4Io
otUTcNgYO2vtPL+WVAefqns37vvA6iu3jBUZz4Bhkt2VgkVgMjTVhZUgum95P/VGRqiKQ+uWdWtA
igqw0KKLyFnOAY6RL7187fXFcRYHO0Ne0a7/YkXsFwD8pbJLQoHECHcjkV3L5q5ltLFP/WpvJVex
IQCk0oaQs3nKTwLP3awEOdNNWnsT6P+WSw8HPISUGXU/4QtcxqYLVBai7g0opKmyG16sTrrD8Xzl
1VOcIm8o0n2berKSQZRLtbTfe7Lb84i/+LiDWrl60Ja66Ruoko+OzCKoLEA0MHbS53RRv4MuGQnq
ksV2ukmc89sdvDcjxNkW3+iscDTz1a2pr0Wv3yJzgdqC8V0tfJ/2h8dRLM1ZgnUjV6dUk2OsG6eL
Rmpnw+701OgJKS2G/bgqqTiLbxeP9o0H/zmarO39/Ao8Pqgi0vOl43dhkAIbB6jUwvh8mw4/NFL6
1oyJqFY5raXHh8FqhiHg+bF8J8QzwbhH7tShXpmiF2RH4rLkHGrNRVk3X1aKROUy4jIDw3ild/ie
GLvot1mcqp02oJ5EOAj23KW1IbqoK+w8z/KyELGc2zLK0v4xS4/pnvts6v3zerwJso7S69RKEoZM
7fSayuuWUa4leanEjAVzv63yJ2OvhHuiNPCsmvv57XQjrrL/GQoHXYMx7AGNEjqX9JLKlH+81Ywv
fBwwInRQUozPfe51TXUcHT/cGNLF6hOR96kTWL4jf/oMPt8mR1BlLEOX7pJJV7HEjHo0Ybz4eOH8
VrN80PZwCkXfolANVVpj8bd+znpYkl7Sflo0BIcBQMt4AzpSY6vJHXzPAeNrHt3lFOED0Q+8M2Si
pi/20Az2AGHdbugqlqpIrL1XFe274rLchvVTEMa1cbdH0hck5V4naDniEFUE7Dda59Y5ywMo4Mz+
/zL4wKklPfL9gqnUkbUJ94gNOXFNGaa3Lwe2GC0HVg9nHmNOVbDD+atn7WYGf5rlZYpXjw2NLq/v
5tuG6EECawR95+hEjFD1JyAiV894bjI/XlFlDwlz84DU24HhWLXjffxOxPV6iM06Zb5w/B6eDrJm
KtkiPbSQH/7YtNOU3vTa/fu4X1lva/O+vMlTjADMMMszy5ChY/t8a5Mm0ZrCL0YYFgq5475WxR3G
MiO0xw3LJVOBfFOcCekC0i1jbsRY98s0WNHmPaYQ0mohX3aJza0EdFe+KLOMeON17fHZGvRa2UhC
Oz5ZTkS1IC1zO1WBdch3w5LPwB8C6Zt35gpHu73aGq7KzP/34a7C5TpQ1BOvt5loE2/avFI7aw2t
PwRLLurRanklfSvDwlCLXfmcrqAS/EX3Wiuu1r1oDSrGT6phSgESgxr1vLc+zaNRRPgan7V9N5p1
sUnQt1aGdwbTdRpaMIlkK0VNIGxroPNp1e7uB4C8HMPJyO8S0rfR+uj7MCN23rnFhR6qpHAa1+N2
0LOBhhLeYr899eLbjXF6vXsxCL+uT6SVwDRzK1t2JCH2gOYjN9cLqyF2BfnP7K0tbLAQTw3Zxbtc
uD6pBErH3x/f5BOQHVHUThCPyhmU9T9OO0NmqRDnGBfPjhQpxxeM9O3tQILKqqY5giBI/AuajJSJ
VowEBt0CVnvUTAaLLiSdpj5gZd+lRO5Cm1b2ytNt3YgDcQrc78PaFf/iALnHD26rVblucngU1Imy
agyOoKTgnCb96IZG185WvXmu87MZhucFAQ4n8MAwqJMwho8TaSzaipYODTmZS3iWbqKqYdFNZkUr
75VtYkAiIR3Sxoa6kc6MK3KnCnfcGFIaYsQEUTEuV55Osp7t7++BYMjoim/h9vHOoXJTspfXMI/O
7cMdx+qciv2Hw2oY940cL3NMU33ScFxRSiZIsLaNWg3DidjO7ITjrcgvlg2lVAgQ+RPqWCtdxfvw
lhKb5XTW2o6bABfDx2euG5H87DmE/wo35tnbsu+qW8TkJShcnOYVocG2MQmYHlbp8SRMvX57Q+fp
3bKlaQRssvh00RfS0IR9pG5KW1rDXlWkME9KYk8Zb0uerZWyomp5h5zXv6+tRYTQE0DpD5M0xJCJ
A70zFefVhjFwOgqXEgOwYqs66Fi6x4iO1VuHyX9+2w338w0PIzeA6FiFbkOO0/yFCXyztVbccuHo
aFTSWMt5cys39lM0aq8zxkw7edSkpRDLokRqdRNwHR0OZ6215UHfUtHcwD20/bbX8z9a+5bg3vdu
QZA2OFk/AfQqSyi9v3EA7O1ahy0FDDLMsyKHNa+8iUf3hSUPoCm+sjdbvYu2VkCGWoGl3R1uu1oI
GPDv9rXSFpcJjqeTVvtW4wsHL6EjYboeWnDA19kgA465bPEnIBzpTIjUoLj/zO4FJPQOt7LmKHXF
iTPu/c993YNkW6YZ+PlG98ajQnKqRs0tv2h/GqeO3gkuln6ymv9cpPYrwB6rMbZZWfF9/ORLh9V5
YAVc+0mwQRRZeXL+j6E05snL83YWtbEZUA7j9GkTTHr3/2ttDJ8+BZoGhAzzDO3aBn4wMK/pHh7b
ibeG0anQxcTtOl8UMaJ3BIXkX5u1BTWy630dx2+ynAydKWLvwZTx8jYfTqcfJlWLZ5SxuIj4lJKp
i7dtyuQtHQAIt9LEVHiZVQAkUGnFWcaJB9LFbHgT1a9iu5T7cjoIStvy3u6EFBH99RvrA9SOsc4z
ZDymdpMO+iwSmiZBdbc=
`pragma protect end_protected
