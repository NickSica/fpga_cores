/*********************************************************************************
 * Engineer: Nicholas Sica
 * 
 * Create Date: 06/22/2020 03:37:00 PM
 * Design Name: 
 * Module Name: i2c
 * Project Name: i2c
 * Target Devices: 
 * Tool Versions: 
 * Description: 
 * 
 * Dependencies: 
 * 
 * Revision:
 * Revision 0.01 - File Created
 * Additional Comments:
 * 
*********************************************************************************/

module i2c (
      input logic clk_i,
      input logic addr_i [6:0],
      output
     );

    // Start condition
    
    
    
    
endmodule i2c;
