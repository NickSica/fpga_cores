`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
R1WqgqFekyFBf+R1EmSjRCQxUuOx6MT9aQyodTNNebOe0CK13nDxh2Wir1luIC2E+1RiIa720P7G
30ynEHVRjA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KNMY+1Jln0fE2Hw6EJV59uwRAjQ2BHIWVdMuSpeAltv11pWP/JZCrd4z/uZcVTngSRY8jZzhCZTQ
WJ4MxCfVaXUWBZm7mY0qLw6qcMnyzincQFakqwRdOx84IckfsGjNGJ3OEjUVkf7dW/J0o6KJvGRq
A/P9gVOYmGcnWb2CkLI=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
sL7gG3oizEXkzDHancu7/45cwKfdv4EnXAdeK54QMEX/eoc5P95Q2IxqcI+tnVljSH1drXWj0Eb6
Of0W/iXPKZ8OP77HA72GpMs5rDnQtlgP3rECZlxuTJ9RMJVfJzzO19m/vMWeqMysX1t8PW29rrsf
0Tqwcs84OG2uxBTuyDEWCBSCU7Yk0aBYU4VmF2rkELqh6jo2Q/udlKIUXrwoYSdX0O9uon++5ahv
mjzu8SGK6zkA4uqzG9ghLIe8qBE6KYXQuzvdlMdTVdy8eHbCbzVTNoB6j51Qlq+S5oMMSQvxBaRz
DIAN76FuevwCbX/XKHESsvee5Sen235LJDeW6Q==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NTwqMfOwske0aroynepwGO4Lz00SLylJkTISN8LAcq5uE8ZoeT6aFHS3yIuZsI6EEE3s5mQQ8Cob
RXh00Ler2BvOA4K7lNGJUpMzGqJI7MZao2GijCVpdWL1r0vSvaacAIY9nlusgQmU63NqWs7cQx1t
7NMmVlpgPTHr3KxO5lMNWR2EuXJ0I0zOxQbbrTneEEip68PBGwJFyFdSjQNe3iwSj7O0u1NlI0nF
01F/RGHelGngznubnZikT85LEu94GTbx+WNlMlaxWaxuIaRvhH8UG7MPhsxH6x7sS5ZS9GHBkFDK
gyo/ARDW7a6331M9HUgGOcgw3trs1/Klf0nskg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
F0eZzxJQxbI/Xk9S9oAxZw5Tpi91CrcqL3BrQB2lyqn9Vl25Garq+8JIOwcSUfEju0nEdI9Cvd5l
ooe0NMs4K3iY8tnE+FiNZhFGnmyV5djhXaAeRPiaySzeXAc0nSnoahW36RgdEHyPbHBrMfq1pT3d
S/0aa8cloJNV0EZcGFq/QrhQOhscPpDi8uk4IV75ihx4K3Y6D/SPBsIijokh2lVOyPsWt72NbpFl
R1J6iXczzSEND79HNenePfXgQ1Sr+h8Z2ujGHirxn/++xFCAHxWZmhGcFFwVO7AI15b3pfNiyQF1
2SACCg7/b/5q/JpHGBLoFY5e10UGMoGkaXNq2g==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eShHfvBzKaZ/Wp/QUxGlK7/6Td59dAgzaJsrKOgtjc73r+sFOocLpKUK8YR7XmM0pkfLOBkjrXYq
jGiy10qSwBo8l2eE17VZo8T9nQ0IB2FFGgVl0zNGiZaKSzE4a7K5so8c5gtUyyVlyHWXKqYAj6Ro
NzUEnqMqJPppbTPQbvI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
VtDvfrNdg+YlmytFZV1nO9Ch/hNzGllGY3c+wOLUGxBvYhloxzDDcAB/7/ljwrwghZilvxZm/DJg
2fzdltt6rugwiyCDZPTj9bYqZhAAM0bSdp5YpZP0gTz8EvbCxUo8+Op+ufZee7A2QX4lG973f4tu
FbV42AkOjECD3RCU/zC8zhB5kCMonmYQSEe1sGWBe2+Ga49sur53s1VC1GSUOY3PQLHNqtwSq2Ra
owo+cSlmwu7mHpq7nDvHG8vWLm58VKt4pglBRfC9BYdbhmSQeWT4IcMsVz3wzwUMY4HmFkj+0Htu
JAA3fKLFH4/svF3ilwX+klAmiEhOn+ftw2QOyw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HHgo2A7au8S1PE/PLf9TgssZhqFUk1LyRHoBPoQd7KZOhYH8iTwJV9W8hjvxzC2Na0peqSJ5zF18
7DRfKJ++XfNw8OtnyxfjOhMGRjIzpk9/xlZOxoCpZPFsl6WTW8CoN0RLlh22HuIAeiFQu4jBiY8s
f/eG3F7z8aDUIS222+2y8Lc0ifWDx1YbNoJritsavlDA9L9WOwq+EXi3pvUCyXszhqfkMn1JVCVR
qUhUx37i3M4UJEKXpk5rfAol3dwNa+jlOtqwiBj8/VnhZxY2i53S+bX3OP8N1Zx5wRoa1UkpaXLd
9XQOggc4VKKTgU9CJZPlRk8FrwN41qv2G8xfRQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1568)
`pragma protect data_block
eeCl3Hcc/V4mGRBHBrnlVFoZ1nOFIg9chMU/4Qws0N/U1+2/E+VmEqKlbM0tBI9fvPVbu/hQoP98
SIVytZii6XSrvJPSRw2jeS3y7db7+MDBncyE3hoFA14HiCfaHO8XtdRvg7FBkdGIn5pp5Adqvu6p
JQpntv6dKctNmH4rgI16sAG56zgsBR4aTAKcuiElJ3GW9ZkWztxkiet9u+Dtcarnf/r0+3HTcsYM
3uN7DrkZgAcW34KGNFH1BDT8VvGnPMuR0Kui0cL/gzz3+2o+XvYlVWABQIEO7nZ593+WvEncfamR
6+GR/6H4maT3GbI7FU32ot0vpTWKTyCVporDFnoLq7ClAkiZzDr76rNjSe5PxHNAhTK3ZmsY7MtE
nn77StD2KyEMzFfey7MogkakyDO2Mb3/lh6opr3YbWVHPhE7kfqaFisLh0ApPpzRQlHLXXJsnQ7S
V1XdiHJ++i64IF8X3ys7l0P6Zi7Uc1s+bsNGlEQLuVH7WbnJ+o0R+F0Bv0pvdSQiVOFlsD1F2mGD
l50k8BNYcdi2rVcqBJ/rmuLyHP4GZ1TKJRGe8yQqvfB6hcoxjYcK0+VXkpxs+UFWjAmkHzDk9FGM
znRzS4ORx7HkkGlkC82l0POTc9et5W50LYTOroA1QpqkPHwxtkm07DtybZpuaQdER3Hjgx8ZLbDu
pbKg8V4LX9rx/yTHBdT6M/+URZlzwxB+DUoYCnz83Ut9h7raZjoMEAuevcFZuYcycpwTmsiZ4GoT
k6IEi84/AhZrNfK4MadQUiN1OnDXQcInpWyyt6M4uII7fA6EdehfVolnLdxKICHiH6EF2GVsH9yy
vKCHL4Z14SuTzwP0Tg5VWK/u9I1mnT2ScREqhWhoPe06ZogPMvW9shDCZ/pevk7kR3PS60azfsvR
UEqq2cRCx24IcCewoKIAy3U4kPc1FkZT5CfEpwnuzWdQB+8/eBmUlAoDjwTXSk7tWcZ1YAYyNlYX
Gz4oX92C3rk7n2CYVLmYdH96piVrj10O7wC4kTJOpTnx5xN6xsfyn5MyiqOw0WHvOsdu93HMGTPh
FD/NROsKMadgAqTu0Mz8FYmLYrOhegqUS+miBxrswSN6OCE32TSFfrdAqB3b8ZD4WNk7TWdAGvEN
4HXZF0bR5C4qGr6RSU3N0r4wMe9WVTKiIs5psjcwMe4Fgnuyewh62fDeh2ouWlBstsKFjx/SQlXl
WKIFBM9NHZEHl13Iip9Yo2+fRQ30zlhWKqp3OsDgkL5yuj/G3m9yzBH7eIXJkT2WSbmkYEt3d97s
8RYOGMVmT00FVNKFnaNKLWD/UBVVoCaZAG7VAy+YLVc49l7MdM4qnapoN406TUakuBQlm0qeG6ek
oJDFGZ0HQHX0zSyvn7BPc59EMD/IcH1X6YO5bu6O/tJWSzdrhAoYK98yCwTnu1HlmWYaorbjt1Vb
2Wsf3qPfgxLRtyvq38X5bRhBRN3ZXe1wZekb90npPUe6DNtb89nYrzO6IEhLfLHyKlFrwKyIdAez
jzMQkkpKB9jX1mtU94LdicTjiCUvShVvPI0QrNFAQSgKOBdjvgQLIdYnHpITqejEph1H41jGcR05
1ZMjc/tYMaAvHMtEdcmV3k8TnnLJc/jbKsDMI57ZAn+weAQsF5qdel+tnqsVV2BWqcf9jdY5pWDU
qeLH7PYntJm5iC1QjQSwoyG0KB9NOPx6wFKVi3CnKekt/he9XhIgK54RVTQiVmniMgFpecnmzsjI
fzbU6adbLfQdsWVH5ZzDUR8YeltX5h5XSQGkvmKivJa0Hh6jpEBgyej7Y817jXXIBVpNSVG/+kv1
8O30KmL1KaXWrCgHrxqwggYHK0S9XbhAHFmg48hvobnuOxiaX/bI8Npb9X6UKXQMZn0BdU8ULlEP
yLmhjyxIGItNw1/KpzeGSRhUYgVm6Q6SJPAPil3VuV1AyZbkWYA/B5snWD595pnItrCTnHM672Dt
2w5NP+r3oZBPm4KgYZ0fFf4NLYfyFxeyiLcC4fqK5sNZis3mnygRWkvYEhAzj/nfO4mkDzm0yPln
BZxtDxBw9P1lDxYmfkjezskAy09gPrzu1oV70QI=
`pragma protect end_protected
