`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 9424)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5Ja4CL4QB91YR3n8lnRKMwg+uHePEGQx5x3FV4ifQba4LJQDGUUA3eGv
x7Kj2W4qEOfRShFw72f6g3/uv6fp0IzIOAdHW7nFsG4Hmp1dDAsUrhiqZHqdcN1AoIgIx4Yb2fxe
T4JdUwuWK+SB44slQba43y7J/lLd0xcI9ZmQ4fm6NGFQ4oh6CSU5jUzSQa/57YYodwjGECqmppV1
SQ/04VqS1UCLWTuDdUWl37wrFtjFy+lPwXdMLDiZU7TLOO2MTg5j4AaxK4V5SsVBUbPm0FiLNgHG
sAae+DOi86Dbb4NCoAw4Go+0iEnI72K9+e5ajjyIDBlyjaHMEYFTqfk9QZ0QNgytR4xD49D+4HAR
orBYt8UzEgqJlSAtVfIvnzeJfkG5vvj8kfbYuOrgpHgHc3VIZmEcA0wg7+cK/VhDirx9/GUsPn0G
O53KpCFbEu+WVp21ShW+PR+JXNUqOyV2Bb7Zv8s+Ta9KvF+0eqCEeVvsxP/sh7uy362KQoeVVMIb
eTnc3yjS2bh4+vAYkk6WdaXEcsvium60CBT8a2XO0blOUb3n7i2yua2XHcePo01ghzL9hil91u+D
C6uBAP6x/67LfOxnv1jXDC91TnikxWItYVu2dEJolL76109X74PNc2jGgJsjh4doDxT4XPAslf+C
z/3ZzQmX3fIhpKvteAr9B7r5efXZYUYKpk+F5MMxdQm1Zr9CQetatHKWGijkQFAYJNiIrsfrge86
aT1Dq7Tu3MRYn/hYXW3QSNzYzRPxgqt0MRgYtn45p0QzteTkdbIhMFM7y7XMzzVyqqmORTzmcXNx
hvQPT3+JAf/sNP52RYw7QUJHSkC8HNZDtou//DV+hEbilzo/JE74TKKXTBS0PToM0TFYXSWcbBqV
0eBjUQCOh1Aarcd2b8gxJT7BJS2MBhVw7WsVP+74TFCk+vAO0gAhjNj6EFPp5xIVWVBaX1kD2yMN
ZlKtYS0PCuFE3DFK2xYf+Nn1YO1u6rj034K4w+gCbSYUDXUuInfvX9YDChWzFLLKYmw3OR6S1SRg
ZLF9mvTiFTmK2BG2+maD9VvdHmFGzPkGTVCX8ASCiBM9sod3UQ7KYunEIXIr6HaJkLXRNSbqDztk
fTUpvB4kkvZNHHNPu6fTpe5RSkWHZ4a7E/I+ZMbJLrPsDDN5P1e+efPvzgbmk3clyb+LemwhJWgD
OpuBvIgqRfB4V0qJWgwAb7zz5zvRmm9pEOoG4r3PWYeDcnW9WUxjjbU04wIHKbYk7pwbVhUqqgAz
3OvfSxmn7t66Eh8OVNHuCu9J07cmbInocinw3j7Zq6itOCjdFcyZXt0nIaJ+yU5ZlA/L72BJd4xQ
gPUJXajvI+MoFF/fHY1SUjySTmWaMxaJYEFMSaV819OICPEAEUtsqQq8M2Yx4kfm2FXrNhor5t+c
/i+hyRqTbw+EV5xIvBIyZK/HAnqGAhk7LgYOJ3PEEGAkpvFqkdvzM3yTl+W9AC+GEt3c5jfVKcSK
o9XywPibqsA/wMJWvpGQ6+vdMMoIPcp6CoTDHN+NmhQiQu/gbFPeWw0mrNbNdyBgESSF4hF7V7EY
20ViagAa4xfJ5IA7Qqmdv3p8E3CWM0qhoQR8jJ7hHj2kLjEiQlF6Qvq5NrrKiLKlLnhpYG2JRqjJ
EaLM4mZ7rdlglDEox9EyxN9ixiOC5SAqd0bk9X7q+MR/Ofq2OOmzvQnSDHPn34iS9tBhNZKEVmGI
kwKlbBEvRjRT2RMlgYyFXIWAdeCOD5xMrf6J7+AQKpislhfUKDpmHlCimI0M5q18a/yOQE85g1rU
0N5AKoI/D3De/efPlkt9KahaFGsbHxrcAw7qZRPQOU1fvtL8AOfW4x8G3yn/4JhHF7Cb0roZuPbh
ODpQLb7t0YKbJiQBXnSzzDazYzJ3wBivbRHwiFfVJ83mURYKHTRuOgNN3DGLwWcdLAqqFSFKxX9s
PPFINCM4RUFQvC4/0yaZyq0iFkW7ZaF6/evcN0S+HMvyD31GHHRMurEPHJt9v5Bn0P8QYTir/nqC
8zQ1EMMGCbTzFfAgoqXHwG3kaSl17Sp+UKATlpB+SzSE/yL4vfEFZLX+Jp2R0MkrzU8JmsLz23Fr
n8SeWUzSEPwwUSQotdtKnho5cfzCKsrtLTJMHJWh1WNK9RKOiFfYNG80TtZWsaVZI6MTwZA3RLn5
4O4bwzVSidHJW21xOuVx/DTQYuov8PWzqgaSxLuQ1sNs1RU74Q6njvtPIjER5N71brXuH0s8grhQ
0NlLSYMV/DljGkRFF8lg9Rc8LImXZgT/wz8NGcprqIkF6cniq2lLrZlbtw4KiZkkpn/AJ3GfmRGN
ftrwiCnRFqq9hyeVtCJLAYWBWq//ACj4OnueG7CuQsTNzvsMkgMl7W9Ntzec74USKnrGJe3952fV
g5nMlGDtMU+4s8C2y9s30575pcnQHH7uKiYxgratAFc2wRDs94ae0+sxXcwNYCS+WhvIM7rTGcWp
/uXsfVUomYZUGMIo6HNbiyiBip0v8FzEF+dgVKVwzrOSGw2r3d+rLVj6QIbGdPp2Rm+6XyUflNEL
4DYJHWEDh7/TAqV/vfKDMSThOOLN3UTj562+gJoIBew8VPiqqpS2qVXerT1ezNEPSvOVAvS283vW
/HDzWbLdZ4FhXWobHKHPFMqEP100NQsyjtpG6w3M0x0JIDBbaPnhcLn4Xh3xDPpCjtnDBK/Kfzs6
O62Acmm0xfDl0etBe+kR39yJz9YTsVdfjpeyPdoWIdRGZab7kk8xKPqIpm8tjDjZq0HLUZTfyaRN
Zlz/k6cvim4mQ8YNpBBoK0KnA14BFj4BWuEbHkT37cyE5fwj9I6cWlfyFI7Wk5XaLy9zg0r9aPj8
WZLFl9h0ph2twIzc0Eh04vEINJtiSuJiLsxW5MTGG5Il1Ff7lTSHclkC5uUE7HbBgpkPaeJ5nitr
01N9ffuhPKI7W7JI+gTdRvNQ44l0dmyiqBAILS0NDZwRuzpC76QGwJ/Z8Pg3XIbXIND+fjXq244Y
8A59CaIm1zT9ff//DXOQW6mxo5Nm5Ui36zBZepo0FGLBln0cYQye2ji3uBoX3AGKPxiYQVrYX6Tg
g9f5KO+mHLx/bYGkRoT+pXEQDsm+l0HBTbkwTBx358xs2vkX2/nK2hdc2ZXevFQUrDrR0bmDPTOo
4x5iGWE6gjXjjDSGe7lryMkHufBJWrAj1bsLXw48HMNJuL94NLIp+yxw4IFTgI56NqiZWHxqrpby
pM2xpUFUb53C2zIHmzvJUOtJ3SewzKV+zp6UequiDLojXBE0EfJd/aJtVDK3taIhOSlhs3meHQYE
DAJsiILUoF9zlV3Or04LRNR6fNrvNo/u8uvXbTE8DME3viSxoyIPZ3tTVrOePMAz+0wisxYqwSI4
FBO0Z7pgRIMC1VCFw7XYjvKxGOCGjB+ugosf+ujmU+IhglmtUYygKa73+RksAjAzW4WNm5gbNLpb
YUEWh/MahvvT/iWkP/5yXq/Wu7mX4KJu8d7tzrZE9y4N1ty4XdwxXAYHSMvmS1Y7pc0mRHQNBxYe
aWfntTOoRZLKxvTdST2KaSwe4e9Sex2s6tsc+nBL0vuG5cOGUaF13kMSWBV1xCkpqZJYH2p9MLZA
M/1HIELOHcyMS1xCubBbmXfiJ9FAlbCVx/EquYWfEJaOEZC3Wjwj2Fr4tYV3yiQx2k8dXFgS2A9J
qGEZgRkaQagiRIWLjg6T5/VgbUosQ3X3NMW09d74+VLiYSFNI9bxNy0XGxQcMl2XUhtq2SMC7oel
FKiU3ey7amaWKvDYfc7dYZbLx95YghyVholjUv8ZrdHXJAxKbFPVdr0L5wA4hEVzAuoXbNDz51hG
/rwhPLYMAZ6FAfPlbtj5LpjK8/6aXKIUGhSbW4dwLNOCORGCaOz+hzC4osC/oUPNPUAtsResE4wq
HWhhPNcDSQ6FLS6qaStmep2pylAagaUy7wV4UAb9M8Ok0uPsfiwyZlZV7uuCghxBQV9KR6lArME2
YcQUL328PVTcIZdvQ89dEwzzRsFH9629x3XykhQr7Al+w3yjZfy2kbau1TiJ54eiMyoKCxxSiSD/
a1l++CDUa7/z6OC37TRQ5NSRWLJQc8MV/Kc/t8ZEuW7bV/PEIMCnPEfm0RfUskLi9Tk8ThmhAagp
56xXmC6X0I8E/a5MsH8xLsLnfpALYyGjC0Qf2+fmGenlxvOK532SHolRTATWlOm/4JC5dpDCqm/6
swIcMWQlqe8yftcYGb59UM9gKcAds/Mudo2NaLQ6ap49JKUNlmgdWZqR3RdC8Y3L1lRSewz9H+ii
xHfz3lXaCm5qXi0v7u2QXbmOF7gMe/eB7tsUNXMq25GIVxmJRiiNutqwW4asK73S+ypwDOpEpSRU
A1tU/tBPyGc1gJ+oGsdQK7egLvnh/TQO9fC1K2Se+ggR5UQf3h6ET78rLfuIVb7MeenG1VoNtGIC
FKUZwhbIHX5fj6NnVJwbIM2NXvNyZoBN9EmFhignHmH3E8ijgknURuVO7cfWDKi3R971MMaWonoo
WIpLlnLp6SfQg/nxki4TRi/a6w9eAVF128elcY38yNOV/Iox3/ww4mOnnBcfzeZUbon+Zn2fR5pe
0I6kPN1tKnzrsCSjviGAd9yXpvcDnek8lZHhHPgGUtvDfoIFIhq+F+N6Dj1DY2xz15MQbrvfb9FW
6Q1ox+ZOROaoQeg8uUiJLM8PMPTO1srucgw11ATFHUs1vPyL0amSrfUg8bomsmm+Fayp6xliWK4D
zLWom+ZWPblSdg+mUtQtrzp80VfhoxFw1jVVUk70+ZbVdDaFB5fwfrl9VyD89G1r50oZf8Pu36yj
hiytGELCYzVN+J39nQokWegUIyXgYiT9kcp8EmC3x8t7B28Yn2iefwDvQPN9exW+m49ecsVe4xip
z4T54/TFi8z0Tjk4glaoFFT5/dzAMpFUHk2Z6CgrvgR77OqKgD2aZp511lEJBxalogyqoYMS9SZE
GMugeg9pwzRAYS351Mfke0K2Bz3I2srPTJ8xwG2Gy3qOvK79VWVj9bkaFAkp2L3iDTRkr/WcvZ+b
WKnJCSU1xnHQUWgxlzD1zB58Tj9E0mkZSmn8TmahFj/p3A0GQXxeCnRFXZjRMM3RKUc3NQCMABM5
h58hpAcs8LTNwfmJnlFQZVmq8imJ8ssfcdJ2qVXMQHg+PNAUpnN14j1u201cT5Fvpij/a00/D9sK
MvoOzknLvXFUkWw6kGncBSdnyVEEGCUEFOKzN3PK775yWvSOVQXdTTwuFhwSKBiQmBwCxM387TAu
i7Sd+YQtXteHGGA08z9Um1yuN2S4cL2CmA+XqP0y2OqoyHEE/9iDZgHozaCCEUhn/07DnmXXaYOw
KkrXa+6j/nykecuh6TrN8G2KQcXHo3X9d0pCeA+rWpJ64P2QryJAgEpYapLVa0eLB+u5opaBokAC
kRRkVTafErH6baCSRA/PynjXUBFfzlB/af9WB/kBBAAYGcT8ZRtCysWbMxS0elfdNnhk9Oqalcgj
oF9fB0gKg6r8M38CEF7i6dxeG0AnkceBcF+48C0KZpytFDSONvxvsJSbAGw4IDrcTqXjYuXyMKfg
BoDbmD/iNeT74whs5o2F5TEKh1/o3w+19FOwugJdKC3LWxtPuQ71SHzQzE3UwOrDZWuOJqWWmPy2
9/YkpFm1yKh0za0WX61qCsMmzgUf7aG9fmtYPXwP/HfDgYJvUZoJTEyU2DMWGBqEyMvGspgyivdI
LJWkC03lDqcOiKJYnRHCuwk2TyYY0bz+Njh3XYtUih265RohLJ6DbjhFl4BcCzSzQfa7eJKqOhQU
5/Mm+IPv7YWeFJrhHCVS3u3Gb+TncUPHpXsfWXh3hFWb3Zkwegvb74MswUwpF8Fn5qjEnetp26mi
boYvNH2jVN5+HzWYOi7+ywJ3fZbGriZhPndbROayrDBC/kWz4oEbkrG2E+xNTTY/ArrY9hicrMMY
aEqTjtUrxEqA6rpvNFajRGhbwz58V+yCEnvvwf97FlXN9w+vw7nAv5F4O7EVv8IHBfQZw3r9gNtU
vT4lmihnhkmVorKG/a8rirL+TI53yJR5AaXhcL2JltpTFBio87hXOvE/cVscoLNcbLahVSS/54Sf
D9jQhSFjUZjHuQ/4YFpFRPGGtdXQzO2BxGPxTNDYNu44xdh/4yAoMyQqJGICPl4vqRciLMMqcoRR
FDkyqXIgUGsfN4e0w/TSkf1E3v9DdU9bvXV1i00llYEjXUHgvN0f3q0WlyRrMwmh/6+lrOItL2Ir
ubGgS10r/lqD9D36LI402KQG79W7f+c/873KmPd3SN7eJfRzrCwpUblu7t/8cHC0szCgZwc5Hn08
ZyKRFOpqW/4u6Ig2a2pvTZAENBkkKS8Q7NnukVxxVGSn8IDLyu/psmXRv8QU+BGBqeeCLmQ6c8P9
9QhUc3rpQsPbcRaSEpK3k6YnBsqNtQxA2Krixt5MReay8/sjwWE4iekhskdKt/VeSTyll7GXbR+B
yqhfrxQO6jbAPW6rfUQ+X2tWczAEnWr3MWh/jjI6lZGA1cBYugFbr08wALhFCPYTtn+zVVa9FsKC
4jzw7mOU7Q89RgZ5n3cpwpaORmA1iPa48h9nlYAZkYpGFjofwbm2l0czvmP74Q0qLvywn3PTc8MX
jLh4lPuL0cMGcLD0YGplIwTwpDKh/THJoL+bR1J9bZdsIiHKP5fi7SwPMqWGgTa0YOS2E6BXYYNp
OPmqGBDyivZ3EzimX8/NyAc44yda+f/79w3nktYQzaVvNv2QVGDaUih5Y5JncytFgv4zARsRD38M
feh7kY3t2uwtBnKWKIuJCuabu2YAMoJ29kpIaR96jJwSkR0ge+d8FsttAQ7CLSyK7c7e10/xbfEn
8t9hwsqbli1MkPreqBrIAm8hrIqrw8UnY73xKFRc1IOmmjqlTPM5cLYLLJ8y4uAOw1amHf5S+bM0
0MKmHlrAFHVAb0ARkUL0dzZPdhT/x1J2my2nucigpvxtFJPlj/XysFAS66mY1wTuCEZz/E4hdXwt
nYJasKHNtlUbRq0eVLRV+DHBSn7pbVGfMLpJwTR0YXCeky3Fq2UXU4SDoci+GsG6cg7s2gVp7G4W
QHEOyehnz9pBXm2GX+Hs2QVkhLjQBX9VUl6Rgap/wAhacx3qa+hNComcU2goT/lHQfCBITbkbxab
zqwTsJnPU8GT/TSRz286uc8Ff3xZsjl7w0hNTez9SNzHmVN9AAW2NhX/TnpyT/S9w5uxAorTRy8l
4cwgZcaDrrVebEtcJmkNHMsmfaYyWM35JO8JmL8qTSGe7Xrr9MhIn/wJCqEBtA8i1UizfQwYFMr6
n0wNlicLugwCmppmEnx3O4Fr/j7K5XtbCI15o+CyWMdjrzSzc4kqLIeLs3Kvidd9vjalaG3mSBNu
N5+k/NkZzuZZCgsvFWYoKM6Ps/cQUmUUlT34ZHrLXVuzxsGQnX0NnB5tnFt/rA3mFOapjSK8MYcO
fY/3h1tQo8sp6SQGKpyE8rnjdOLzcgb3OHfsVKPVtQG6EjZMSfutRPwlyKwAQECNnNamShsvBu84
7ryGz5aj43mqKO2lAE3du8Ll8rJavjTrqdFKRcqXLCmXKi7v7f8wVjjOSpYhWuCRYrTXP/Hkn9gN
lawvwpUN0GpMp6KN3PPCLfiBdc/yfxfO8DqJqXHx06hAHU3aLullpZ4fCAavwvj4vI80bFvOOSMh
tOZS1a8ZzvtnQsphFyR9tg0TKIMuFB8NAOKZrpwBuKMlhkJCDBZfM6iI8KBH2TwVG3BRDvClHb5F
ANTcbbQhkqcOPT9ZwunNSFL6FFi/snooItopB1ENMRQa4PvruYex6jeLty1I+SdwJy0dZxK0dY35
+oust30XGYWuc+Ao5x7HE/LPq7y66HNRplqFrEYH1Nu7U6BdKyavDYwpK+cypgrg8qn5cDPQWaF9
6xuSmLqJh/eIEBmGoKedsqsj+qV9Cp9Ygid4+qJ/TL/rywweh/ZYANdaXbxE9IG3g7m+vF+ylVR0
DljnjDDg9vRt6JUFFkgz+2IklmBp8k/BeH/gBMp2ESw3ASaBZRpbUjHrt9s2+fyPBFFhRQEUE/J0
SHC/M/7UdBBk/pgrGvxn/T6XUnSMRNrJLsWzqo1s+SFz5d9ty6AnPMq763Tz6BMA6CvbJHXA7qL7
ycBUlf7Lyc9AumznThovpeQgNEloKFBuU25t5a6jha6QKmHfFml1JbLZNuGuZstYncHBV0rNhCI9
pHa35OlNb8yzmgSERcOEO6IssJi6Ep8164U/skvkqRN+RsJlIKjLoIsSR/Z60CdQgQtti7YE/PHA
FVOmzJWBJBhkjnHM20thhj99k2+YBiwCEjOb/t8lq6VFLNU0rcxwwmixcxPwvj7+4Rcce7w2y6zG
6UdeRDigJihW0N/zI7CFdKU8BdTckSYdNCdgMgTjiewMKWy6dOpYo4vTQ0ga4Icp1tU75HjAU3La
4TU5BmnzFrdE3HT+zsQ9nuLz/MzJAQBghUzECpevjzbaaqGjLaazYov5KZXFT+2Hu6VZvF+grCy4
3NVDS5T0iyvqGmJwQRl5hYNccv9LzIhG11dkeVbD16ln17e/xt2ebWGrS7zq8We8zz0zvgu9F66h
nwAA4jUvJ8U/YFEYgk2Pxmapn2KmlI+r2XT7F++YHmqD3kBJcY2jMUC0WeK1qZR8wdnQfPJac+5U
nypQ7nq7lQ+zVX7W/W3AbmpQxeBIPiFP1ZKa2HXKu5g2ZEqTZVmzQx9RyDjEPDweXB1BnliCaN/B
eSCXnVeCCT7cHHn/GSoYGh6Ho+zHvsxBlRtUWtFyGEi23GMwjhmwmY0V3cH2iK//b+5EPgUaf1IM
HtlLAIYGlVCPwAXSwZCrSV7CMZmkFlQ//cEjuCAO8Jhd63vGq0EziKoXI+iOyt5y0qCbe2wtj6/8
79zK7Mfn+5I4JD8z382AXRHvUJ4AXihoYef3T96Rvww3weAQEis5F5IAFnRVtDj/wSFAPZE3FeR4
Ld+pWACMNeJNC0wE7aT0dbIPUPbKBO2LapubVGhkBLKPCYn8sZyuAfiTlbJ0WPZjnKq87TSndYbe
OSRhsjjVntQBGkv/JYKgNdaT+IU17ldFW28OhONOusa3JWi2H21J1Hti+yqnCqiey8apmQvW83Ki
SQmauynTwcpGddXVnBM9cQsNjVLhZs900u6Ks8TxUf8teZvHO1VtthlmShI0pRslgG42BxJdU+0W
v7vcWnd5Vxkeb6Wz8HfVWEA3/46ahs8uvNXL4kmyUr8w1qOxWotuiASO+UBuH3CKdPz2tl1lxSgq
ooLO8tVweSCU6eztWhE6eE9GUPC1fl0pudsilqgfZmyWV05Zh2zSckjQYL2mfDYfiovubzhgaF3S
MCsoN5QneexXmsqBWszJo0D2IOtzohb/Q9d9/m3EVJu40G+NKAHPbZxuFaYFgTCwCOoVkrSyAhBy
qHoCr0f/5fQSl3ajZM7IrSDxrzD4ZUc6bTZ4MbOg9Kp+GzzVqZSkL9UOKBW1CfvoEXP3J5ZlKuz4
zT4e0sQ/E1X2Ly49dVS1s5Euvh6opNiusbJlML2dYcjOfqXMHLNq+90+7oCzm/J4GTq1yMkvihZJ
+FMFO4aFkV3R+kp5ld4VOaRnXhjdGW67j5LZlmmXzGwDsrqcs5/lFrTk2yGqskvGu8HJciFzV/jQ
uTmYpAOgPdQE237Th1qJDdCc5FPDqmNb2HTgpR/QiNECKp53tlTmOYJznCyhalAwVkCStCn2jvxe
PZ/LQL8FZAB13qvpwjKnovKvL+ogrlgzZsQ8VhbVVVpXSDzUgga/zdEHJNDm6356QQxgErG+Y4wk
2eWgcIjKqmsmdhKmJZAID+ScoWrAQ8tAdCx7PnvjUsmV88IZwzVLuTJdybkAb5g87WKq+fgiO4z+
ufWXB+BJw/EeYovN9KINiYf0TrOrCly83k85s82Bod6ROAfat/QHwJL2RxecbMYeJfnOWXCh1Q+H
ljshpPXr8W+/cBkfws6H+JYVfuCRttBNi7hq6+Z+2bDJ/rB4p5WhRbALIHlFbPRzwmcZIdVhsEG5
Z6zt34UByHGSd7KcebUUkpmUG2lCJEyoT1Grrf5CMuycr4ZU0dI5jl5ZrswwtQlDmUokikNTfeEl
fk5wFu//VsT+RSI0o0JbE5rLQowMdvDwxyqysy44CzE26eKL2Szyox8Tzy/zNQ0RN4rjmse+r/p2
VFo9v0WEXEaPchws39heytVq2kJfwMzA6ouN1WfCo36p0rRLB0nbe6jw2RjsoQMGQCAC7Pov6N1Z
FJjRgWdtHFJfLz7f4spqXyiJJpKAcGmnrqzCskLY/S2HJ3OvSp3ZbKBZIuuERqW1R80cPvWI+wWF
csT205zgJOJWpVdtElHk0ioHBB+26MFE/p0QzCimIh5q5gaLgJAo88+maDXqgK8/V0YmK4qNCAzg
SEUMQ9UGYt8VKZUyZKNeB/3p1vqpFzmZK+EVxohwI5gyWs1CDON+cSaiSSTzee0FH3vE0vzux9T/
QWUaL9hO+xfOmFm+jlg9/+YTfOLm8zJEkHlKMtjmEzdkCORcG/ZzctKE2wT+loaurSq/EBmBNe1N
LkIyGJvKYfugju44QvA2YPRorkbr1zmVZx/DS0t3I+i90Dsg+91L+maMeOcxe7XHoLvKORtcEJb0
vyf0CbbEvvoiQxw0vp99XkJAA15kDhoZtkLAbrsbQeXsFG5QE3u4otpoSIXDC10KMl+uANHU+T+G
HL8gJweOaCurGlnMitp+GLtUzia0yA7P+TBoq3rsSGWMgKT8l8UEB2ApVhmrQQb1jf5BGixkG40M
RPsr+syZLo0oeG17nVWuxuk7rNzzk8kIBSmS/sbIn7zPECozb5KV4+cet+LQn6eEdBcHfGX2Pfdj
tEf0ytaNmd0BeZ3CpO2NQYuN2ZkQWV25z3w0ayayHIYnQC4j1YWhJOjEwGOBbQ8qjU9IFJhbz7nw
KDbEBqdZGs9GQjG1iM7d+fAC05orBo5u6BT5RCfOHLSI8PDzmoxJKOd0pdIafpApcKVP59h3s/DM
aGbqj1iyUQ+F4wTPAXb1y43GV9Lzz6DAsXYm+L9T2KvqxlXfQ1elU++t1RAG4TP3yBIheI6qz+qS
8CCClqVzuR8fRKcjLdya/rW9TKFs5cr4/FgVv9mlTCtpGk2nTxq+UhkKH90W3WDjWpB0YneduFeP
QL7Pg9Bm4h0AaNisAU4RmWXFWsXdSZU56AHv/0C2FaAFmRxZqk3D6T2UP2lHNP8wsIJK0pE4w7T7
3olP5Jc/8l2yYjJB7LDOHWN9yVKvkNSKhTxL+nRqk/fCsq1rr8UiG5OofnbWl5yjBgya8wh5Uf68
GCPgpoQ/hVe77W4auYFUnW5UOVHSbB+sOR3JBu+bsjqbuu4qQ1PiQ1AxiT1UpOrMy18NxOAKo0bk
QXXXZeimqQZf+9+m+GlcUihuKH9KWAd5lOXLlEKeTXTIkt8lb8p8zrIaL7pvge2ygN5xZzjni77M
Ao7cTLCOSPDcvMFpNMzrsDXdUDpajNtb6U5+STdt/7bpwGYNrIPSk7zgY6fitjQQTJ7ozfNy3Xzu
lrat4lajTXRfUpAuKLsmrhf3SdpEUUbwn37uUEygmd/XWPbHqjj/4ZuqhgGoS58e7acqRzN42Lim
53PpCEUdVYEHC9Wp7SkIl3ik9Bh0oM+2i0GYcrFEPMuBFbUb3DBmFW8kPJmpiRYIKb87pFVOe04h
PGe/dje3s7HWq98vCw9KRf6ZX1fA4wOA+HEK/04VOuqHEwp0LD2KZrvN5AAOKu7maJ1LXDc4JM58
RFyCrJu8g98+qaE+Ie5C/9p/LF8/QaiDGKFbYcBqylbS4WrW43joYt4e5raWgUHfS90lHHAXjkl/
6B6HomxrSdKobkB5vNOT+tE5yUuKroUogSfnozKreu4vGX3U3YWn4odJ8AQ4DMzXkZs2YEqUJIpk
qO9isF7qge7jzLBXZibGozu0lY0H20BbsCRhIRqMNd7sXgygycnbPmTDaMCu2uCYuEpXVpmS6WC6
Z28Abw5X0yxGsNzaizEp6PZgjLZCIt5zSY2Y3o0ELLlPeXZQEbyL/FXrN7qx2X94FPH4WLsPLgYC
1oR4isVzXqVWykGobKqwi3q9bjYV/0E1MEdPuuz7iiZ4hNPoU0vEF9eISGtj+utT1G4NZ6pfq8qc
iKixRlNn6205lelfhIp8r27UWulyyKNFmBE9y+cXqYB3WmIQVQu5dzhQpNXNKR2TGoNcRZenlRON
x6RbBvbgou+ziejaZQNHght2/HMMLbxgwqBX4x+C8xvTlZjAwhgt4gnZtA3P4kPYaf6eh4dUSHGN
knuMSaLi9k8kJWL6K151Qa5gTdgmkStq6Vjs0YbEbM0GiGcdrqoFhmMq60hlBWwIfiq6Ducn3GpK
pfMNKuvr7I2PMi+Nck6zqFJrgepLVbgRPnpGw1CqJXG8MT3dO8+N9kL8foom+CQaiwV6RW3eK6dv
lZTxxISEfy7zK8pk9CcA6ZTBsg==
`pragma protect end_protected
