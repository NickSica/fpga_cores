`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
V82h/mp8FbHcv3//3zVZ5VW10Mue/LSt5dvjsUkiSGtG5WaH8H9Fv7j37k+xy+3/pQvfXcpqBF/k
iaz4/vETUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n4WSOWV3uUjyMD/l4IGcKD1bHONRRplCKgax9lu4YRYlORLHEpckVBvOD9geZHtnlLIjTLNUcuHS
rc4oO2K5x66eEf5+m+hNzaPYWCrVKWQI7/tyX0imMAsD4JQXzU2CP3ATsQoldRyYOQZmggmbIMiB
stLQ3uoRuVc4t0kXI7U=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zgo3FUzRcS1G0FRTCr4C/JBs44dp3dv5CUvkYU2vM2fDyGtu9ekJcjDXnFGi3Qx2X0BV1gEyWxsJ
xqQkFlu/f/1mutspkUjOMtKZNCgPGDHkGfwBEPN/xT22fOBwQJUR+Oj5KSeDWe2U4t5UJ4XXcGMb
ZV9syPFreDWYOTWkkl85cAKcf/WXC6oz+tOUowqV4nSLA1PaSrK4ohf8oaOGNVX+4Ji/w6ViTIJJ
OqmPJQ151npm7Kbt4RW80tp1OmABkNI+o6h4rwtTS1IHzM6bJ1Krrp0V+2aEmmqoZkuKINjX5Pw3
P4Vi6iUmJI0uMpdsCPr3MEC8HH4v95WCnjh0Qg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A45QQ9IEoKpoNXpmniz3AuFZmGAAZIhtA2hP4/pi+Iwurx8nPI4ZkKpYXPnn4DfH42bSsec35aiS
Ve+A8f1Q00bmFgtclspinRe4YgFesk40ftn1mzy6g6sLCNXhUm/IIjCSNk+ie6jVQS7STfOdio+z
cvSm8QQePoJjzlJz/jkNhsD110PhDAevJWb+C5fforY6kT0k7ZmJmE7btahod6wU3o7t2HM6+XGU
DDNZ5E+RLS+IiJYVCOwsdqQFDuRaWwS0k8Mk4UuDiVWtU0+QLFZ/8UGJhy2ZDSYlL/8TrrsWcD/1
Vku2N+fkWCj38RSMWEEe5TmUHSSzP7uBI6QwVQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b+wEsHDGMmVXUM545W/2toIjDItLsHFsIOyFDid8Fv6KhzBePVZlc9t2c1LfdAa6UEpdqcx5kgIr
+oVEglJG3R/fb6dRp2mvlu6+x0AYh7FK0My5t84q7uKZ6EPBxHnDds9FLGQdMDUFv8E10WtGrG31
lkto5q+L5WLAzYgiD3//MgdbP+aqLc/75XWIRhw/PfRn4OqyBU7xSBeoK9TDxBwOscUv0cQ+dauJ
dUQ0W2ZCXwF6cP5c47k76Ikfu69J0/IO+FTLKMkjAB7Wzsyqbpl6RMVdJ/iYscNROh1xxo2k+52w
4l9VnVKN7wTWZdW75B3V/MsNTrKb2I6dBdveDg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyn/owx08GdB/M0CwlYM5XwpK1DLRGgNdNGvCa53fvz5ftb1LM2R7yhWTTXlm8iqXlg1S70wvPmw
WVO2ZNZ0csmDdQcX4HNMiokrI2gpR08Dk8n3nzdOhqyFyh79/eVJzQItyKMQmJZNCvFfww0mtX5K
FbNe2x6ria5jEBEBp3U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J8WwILioFJtk4e6vNsFHYZhWTjvAMbsqHcnvhYKYzsY6fpaoYuWnjTNNNxS6JYZj7bKOFgPjdnBA
rKaGPLghV6UU9fx6UcBVLjNOj95AU3CZPEjWGC/GqjGRPxOkhGtDka91PZuOBRTBqJT8F+5qIgQR
vO7WJHaKezpaUm2zbeC7+ShM5p4Wm9L4dzJ1OuUGZNm39p9FbORAZNzAWa35wpfJ6PPOgATFMi7Z
sN0Hg00oxMFCKSg1bxvN3p4iC3rVT+wV6yuzOecq97B7Fu+tfvP+shqnUhodTpF0WYfGWHeK9ocM
Mg7nt62XJybi4Tm5rgYGMIIM0i67934etK5Aig==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AF8EDKLpUnsf5U27caIfzjHsL1dKCT4FvrlOxjBwD3ZJ9vsXwbWO+EJTOJOFymKnoSSFnuslr7C8
ZCAbkJJLJrLXJwfvC9hiPRksxuYzuxWrtwsjJd+5KWtue3gL5kHClD8Tbo/V+Dnr3gvKzMRNdFRz
i+4p8dC6/32xR0/NITJMYT1uOYu0oBFDHGLR02Wn4PqghcTR3gQMVeL0RsDhJibeNnf4Q0NsKqCF
7OscDpis6r9ZAFao+mdpLGI93rreTlZvJBUPh2RcpqOjL/8IUv0iM922KOCZ6j1LtvD0igXehvHa
5hOx0DDcMjOoejqJiwIqLij0FB13lDBsu+fjWw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 87328)
`pragma protect data_block
BMP9G5RAk03qFRu5UmzfhEl7ZrPdoJV4zXjowSW95Du0rYzUwgDEcAAWWrJkGr8xUSoALX535mtu
Z4wah2p5r+DkafTouvOtf2CqOUCZEPD6lKpfdkkVRyUhL8kXrCpzRqWnWgEOCQvJKre6qIjIOyK8
gsdAK6b0x8mtSkXmGDuXExv2Nf1FUyY5gcwNPZPqvsMQbM4VgaI0WhxM9BdRxVzpGYlueUtIo/ew
+/v3pRJIbR+CCCdLwNoxNOvTwc7QWkNTDAhBU/Uox7kAREWMU/tKNHnsaxsJ2Ri3oxJ/ygKc3a/o
MyyH2s44CB+QwgzXjPlL7c7MSf++gT6ETDJBuA4pyNnxzLlf7QAaQ6sJa0d8955OlrBm1bQsa4Lh
kgBjAuefHFMQv56DqpMABsLRM3l754hrYBZmziUG+m34Wc2XKi/BxvjY/seeuD3fDguHk3P5xm8T
3CpauvYviidzehiGdEwJ2hbhZEuzXN0r4N5q6RF7z2QroQUNIfLPepZkiWdifMftnmGEXX8iYxU9
RBg5oaqXuBCe16iJBlufMNHqHhYzp9WCghD7DqqF2BMeDfT+KNiOxKEyQCAnytmahSRJlpfEdrPJ
t/joyKGMtW8jtZIr4xP4gZcOyfr7joIkxGFbl8BgAZFeTCVFaI337rcidDwBa9S42aZcAxtc5+x2
L9o1995VsNNGKY0kdqVtrEWMTswBbn3XobiZOMjLzw4WdxiVTkKSwcrM2QKebUxfxQb8Zr5Rps+c
szLNWJ5Dntm9N8nimDE2LIDf/DdIh+GfJQ2+UthTmjdtR+70DHruboNgOK53EqGGjcyhPtERul3d
70wpjoPt+eG7zgHqedx0EjsY2lF9Voo59jNnlKWYPd5jpSjqZRuOusrmlX6gDMrcZRyJ6CUNTAfW
vsEtEltUfO7t1a1mQA9sNXdnrFa4QSYzA1xygWpye3rumWjgl3V+CqNhbV0lSQpr4ovoA4MM9UhV
6gIBQS+ngzXaYuU4iRCiY5CcPeJP010TJTRgE5d+ZY82a1cCuQIrbIboFgs/oDtOUhxzrxfPzU8J
JL7djyd8Ojzuj3wSn8t5Hpgt8tXik6Swq9IOAYFVojTZ0Zam3bZmJ9pl1nK44pv+M95bwUnr1E4n
dIxOXS1xdJjzJPojEI9r+cyRRfSoGfdgsEo8FGoro0+6l1qvXZH48w8YiS+TkLhVDuY2hSibJm4Z
xx6BtNhz2sFLFfJBzj9KGST40dr/JNyX1hhy3nItBWuumptH9CG9xWxTkF+2idYz3vTu5WLNQs8o
x9bXwDitxK5DbBik8FA7JV2FXLJqu2MFEmql7fLmqJvzoHj8lZedMcDgRd4U/3a7D41W5sSuXKV4
9z3p/ouQMU5I8zpToBhkKNvlgeYhSPXXXTh0jOOuZZZWy/ZcJFLNENY4IRHqT7Z++SDGdI1vp9RS
eQLYTSA2xT+COOkq9UzicV8/mxkGx+MUFPL854awlYYpmYE84QpDRzPEstqocAQR4QswQcnl9UzJ
elSVUaBilt95/kZUI4D9UEwYZbaFs++T2dOTZJlcLEPATBNkCx1wJTgHehIXS3y+pe3smXT1+D69
RI4noj0LZuMx1saurEJKJsbMfjArwi9KiVxBkrB3IQ1HGeeVSJpJeDVkMJ+HPPTrZt4yR3kHbBGg
0xj3rHFEwUBkxeYzAQG0r1Mbv7ha7UFOcOgYB5R/E4W8IyqesXOdOi0fwUaYHQ6/ZzOtkrN9GBky
2xTsCAA05nPQS/3jIY5bY5WRRwZtxxkcNZC5YyJTxG/ry71eo6mdfNw3XWbj3M92bH1/T+gysuhM
Y5a6XYDhf1atJUrVd4yKBj0qhr9C7NIpaIpeoZq9qKmzsV4Ki9/hbbvJ6FbpuQNqqX3PTfWPjgHH
xpv+UKd4Oc9cagGnO1eV/9EldmCDijJGW/zPJmb/Ly6UDkirxKHlvEvzpCAfkDIVk0U3EDopjtWe
sHr9j85RFhiczPC5X1UWTDqqD9v7iAHDEriqyh2MxVWPAGU2ZNySPLxkFsF3+S+uBgOB6QyRpToJ
aERqpkh5rqsALBJtQih0BF7dYwNpOLFc+aXNxf8POp0RRJ7RTFPPSLs3IHV4O7D5ANnmNB2oSpwt
1J8KcKb0yJcXmdOwsMvvBuFyU8WejcqlOweeNlJXKHwgs3pjq+7sZDlDREodVaKSH/PQ4gB6/LR3
jyKoj4P4G6sdfcwX7jBa+WSq5AgE2q2mgvI9LDqoXnjdihlGdFPeM4V354q8m7wXHSpJQx3XwuJx
P71JZXRR21kvmQQVGZLsisdymuP6xYKh4gxn+ClOZXL74mkESK/3qcK0ZUsymj8AXlkeLYVQheUz
v2xZcA91PeNmf2nYZA7PzXsSuc2NnKS8rcUZMwmaoyVQerkAfDwREuzUS/e0jN9AC7W4/CDiljRE
AyMbjtRjiV7Bhe15opalLYQ9ZOVlWpO2IoO9xRWLH8rMwVe0wvWQvIt1ly3udemcNSvF85/QSrSu
cXpbW1zUIgoNwcwNnc66qqFJOODxyIDTQydUFVianT30KvCu4agEim2fnJtyYTk+/JBtiw0Pdw90
Zeh1O+96t6eZX95YaXsrZtaUwwwiXNGlX1CQzwaeGfFNTLTg4y2FoFuHKMHYfhD9Qiw7Abkm5zfC
m9yNQti6R712pl397hnwF9n3AxLZtXclSKK8FCsRnIo06AL4u60pk4khJjOb1003Ipe8A+n7RWc3
bpCudiDGAdWLUoeMTkKCKkoJ/i+hfWirt3po8xm96xlKV+UQK8kIsmk1QOaS2LYlJHT4rHxvIVA8
QqirXydiua0F6NQm8iB74ZC0TRr7JYC9r2gL9QAc4DVaNZw77eCtUlqVpI6NSyWtr5yfQwh1CMdm
gJTrvJQA2xG4+cBUjnOe1opMAq59elsLwkYnBoBlvq/LceTAMyChN5HqtJvNbTbD7GcpRTf+//xV
aNILIBN0K5l+HKOFZfZ4tn+GPPwfCuHivXOlal4+X2U28nhUU5VCL1uNbNN11rDie0BnftJJhJix
BvRvV+n7Qqt15TGgqIbQDZmmsoli9GlKTqqO4bSFpxbYAorQQtBbvAWK8X6pLwAAnPQTQT7xaBx7
cfLk55JR+qyx/QS4Yt632b9TsleH/xV26+IiG8XamgJiOy+aUENljhdnylTW5s2yoec9InBEmS6a
OVYgZm2G8cYk+vI9Ek0rLG+CiutWTGXESWHimzVG1EtMYkeTV/9MAOTqaRWUjgy615wDzUGckqW3
cyfRjOy3VxBVejLAuGx1iTX6BHqyrAmKoF7M+RpnZ6lNmkkSTOV/U9r1dtycQhKwKIG3F0vyLq0F
P6YOyPp+Do2v//9VRTKvsU7vVNNPT2KxZTxi4q0SKrRZNQoVGS4AiTlC+LpOPLVQ7MXaQPrtla0g
gUE+M+KdCna1ah1CYEFWaXASirhgVJxfWgLTFbJJ1flcH7UTLynLYSPtek/ihthulvm0zR3TTjUi
rAY8ONoIJXM/VQqF6mbB0Qa4p0AVkv3aUdsTP8PS4jaLV5aJfTvgBMgpiwUw8YSwR8bSj8CKBJeJ
yr1cOzur2/QVrPgXdY+sPzGmI6xBzafxOGPfRA1+MTTycuIvnYxXea9xuR0yeXvatLM6+bev/d/P
pt7eTKd3pVXfn784VSHOuta2HIDvE1XkOGNszehqr24H5saV6U60bPasp1FKBlYzsu3XpEWkeNMB
JD/EFNwz7A2dM0GEs/FiAzdXaCa+TN2XA3qjT9SdKc5xlgtwIRHlWNCC59o/yvv2aNBmOMFz70v6
GqRJR1t7ZqE9JBFZdMQUGFiC8I4bV+zLCAzOolzysPu4B64O0L4lAO2XthtpoBb/v4wgbGd4NGBE
4wOjpHcrvGLePMVkMY9SVqYZ69eKxXDxIWAmnoo2u0KI3umA2U1d8H8NOUV2PNcwxP7ldezw9RGK
xavkBboRLyi3azSFLm+USsyAglaMCpkp/ikwXUgRsAeEE/Dpq4uf2XvItVELR27pioVumKukoHl7
uy4HFN2EdhHpZQq4vjCfPQ82fVao1q3hkIaRbAj5Nz8U6wW5ufEBE2i4dqCEUGgjSl+7WAEpZ0XK
Smhr9rJvXQZqvOv7ygrrkalW2GJKZZrPhExiNH7j5crKIT9t0IW4kiElZ08wgD89jtD5zULzOu2I
YixMcgeX3tXaeK86i1rhK3taYQNZynylgvH0BUW5TKyb6QqmWcMbfqXRWu3ND/R2aaWJBxFy66/U
1PHWvlYki5eUhi7tr1jXdc664f1sD1iZuZZTooFoUxduroA7No4rQ6FTNadFkOFw3MODfm6fiCPP
wFSFaOVn6YQ6h+eOPG0lTT4hRWg+C4FCSzhx/gnPTV9DB0aGM566/eZxt+b98oKjZ8Q3fWYOvMps
QzUQQ3msWJZAUSM6aBGlOkMDj9jKqYlUcIftvaZ5iHmJGsPlZsTGWHAUrtI+4QirLGOkIIP7/7gK
Txim4wuBjoJZKF5tGC3Vw193+ouAjsYgCFUPphKk64YZfrrmCClSylhrtLWRK4nWstKkniFhFsc1
nBu1zy/eu4VJX1lZoKm2D5pP0KYMPJmgW8qmtr/+VVMB7PeZS6NNOKMHGtyDIdk++SLMIgBgKM9v
W7F6IzeU43mTAIDQpXe9xntCkQc0V/fu0NRdIxLtGtqTgnjX1RqFBN87fkGRyNFzK8tgo6AuyXEu
3wVarHK4c1aHo16fhwpJkN0Xg/Ypbb3WxC7hoVdaqGQrXhAlWVNjQ1mrW2UoPau8yEuuqXHQ1krx
DBdOzPwS0l/hUWR3cpRfJPmYi3YsUITv8oBvKf5S7r0PiCU7qs9B+mrRR2fVofi/rffgFHcsVdos
52AW/SX8H5zofvy+/n+YkQc8jiReL6CcBZNos6ZVmkJNJfWTub6Rh5maPWOEAwytQXu/ur3gLguu
Rg16+bJGi/xnedJapnU+Dwf8TGQ6b/+zz4UXbORVDCRbkswB50tpb7nx7LdS2zuvZPOWhw7NBQTa
XZYGzDKy5xP08A0W/mwaEZ5BUxBddkMyv8DGS5eZ7Hb7O7K/MirJI+J9DHkCBB9ZeXB+dcLig2wz
ucBeFHyM8tCQAGQU55vwaNTf68d/juR/tJcwCJqArBxj5M8rltkSuGWCQvrlOygWydd58L8Gr/cN
Zi6lAPmy8yoghm+ReIw3ZUaA/eS+n04QIKU3RDy8rDLsDuXn2B2Aa/GkL8YYlSjNjqCX1mgAWEkA
LFgb+GXcsaN7PFli4x/7gOu02/4NlQgUHrq/X1Ua885fEUdukZqLKfUORFxptyBlydnWMJpoLNpj
4cr+ThkIHIVVxH2hzhWs8tDBKMOjiTcshkd2//6lOLtfcncvpgOkTpT5hUPxqmf0evHyZe/O/6Q/
v86N3UnDHsL0YHiVsDSNGhZF04sSuCFSi3EeC7NjXHfoeJaPJWBNkks2b0KIw8f1kJGGAcawju+k
ysL92PzoILwYOougpyFVg1pRVJnrb9OENWT18+rYpZ9TqXyA8V8mnmrnkGtV8qAxyZk7iSvTZxVd
yynLy9+k2JtmQFvKbQmIPRaR8J7oYQpGxvULmbRdreuAe+52Jdj+320hZoW3fL5a39VHaXCfRe4Q
TQjLk7pA8aT1O1spO2BAof7ZMbohjwgPkRF3h8o9FQaIDeiQkIZrSjBex1hih9aN4x4mnjAW7XE7
waA135mZ41jRYznwVpDxDMcjOxDQ/VmaZ2W1QyNtUfiFvU7za+TKexTRa/SdJP/RTNVSahsY63LX
gDQ8LqMsfjbPwyeFZq36OuG98MPUOOg8WMb3yL2mCet/YnjQp1lar0yBxr5D5Ab+Y/U71x1+RG3c
hfbAI9xhUB5VgaTphWlHgNdN4QNSMvl9pYjqlYhi9ebjzeeXbWYrojV4vWPUHQi6ezMsMKmdkSL4
B7pnIG4Inef+00JqY5Vx8qRWX3TiFjALnvy8bDE4fH5coWQrmNoa9E01ohkdTIc9Je10XUemvpWU
bszK5Ai9huWTBFODAOhFFForaXb58CT90AGKVLRuPt6glxDjIUWZH2AmcvgDuM3JksYVSEpt4P5C
BqmFRjPvni1Q32oHoObghQrxNWt0/EX5Oel9iEjIT/xuJoHRaiqaAXVY0o+8WCBDrh12114RQDy5
lybJzFxyELnDrDyEV3e1p4vTK1sin/q9SVsT19aOWoWxYvopQRO5hBtcYB1ctklfVo5S5KcIwM0t
MHQdXMRhcgU5twjoJUTkkgDw96bSBrDzCr69BBwv3ve+Pnvr7QS5Q7xhINhTFJyNhYtOcXqLxsKM
Xym+aUf6wVIBS2zGVX9DHkQHWVsbpPi8TCCTIhryTGavryqXKQjpOOKyNi/0zeDerngY/NEzLUh6
QMKIiIIA4AgtHbw5i79QDnif46Vrsvyz5r/MNJt+I6GI/HIjpES9w99VkOJEGv0Rq5/oQnpBICaR
tVAo2e7rxq84oApDW/zub/Rb1qAfDH010W1BcJ6AsDlOzuRgd/R5TlwWFx2SG43rK+sre8UMw/DB
3nHVIZWp1ri1ueToDUs3+ijLQ2LnZtjx7Do5wAMiUk7bNTWQlhZT4vTLvn2N8D32pvTRdwRnH4qN
TgC2krZVylc9fQg2mvLwVZEtCpLXekmeLZ4oxt+GfkCC2tOXnZgecZ4sTAqC/7DBKt+9nhMtr6u5
eVwl7cOCw/gLEHt3//t8LaJdMQSSYIhjOG88xgPE1alzoT2h5PhBR+q6MTRBkTa1lGiWR0K+urQY
zq35DIbyXMPB+01HItmDYkY/FsjXXfjW0+y95Boy5lCFRJvS8WWVSlJHUYUcfaeFnbs8RLW3L0r4
YQfn90XPchtiZnBs5ygI0XaO+p+SymHktT7X8ySvYzhO7bQhdYWLO89Eo8kRkzIAVmhk1sotP0/c
7mIlAGdQqglIfQngOqp61XkdJH3Ytiy1jjQYnD9eW35AGRRHssjOIo5nn2Xg01BGULryjeSLi2gT
/Hw6MAlgl9srIVfrkYBxCM9i/kglDZVWDu1YoiJTPLXYeDPETpaD6wMSMHLq83xQMED27+gS1pq2
UWObKO83v/W5btucLAxxYhh+H9AGwsSibeFFaIR0lB2TAELYKG9Lv+iu5osLtK0GbGMz4x6FkqTu
co56WRpBlCkRWuLbqSqsQk0eWB3jlxNtAv9z+jFiyv/sPZ6Eecy2YEjMLhMyOS4sGvnICXvlgKDB
WVjwbPaoOAVUA4mLjI0s1oOaNtAHGCbX16rlQu/PZb4G5XbKxkL22h6S36PWFKgHrcXxaQmvSi3x
Kd2yrIDS+p7kRDCBD8525NI+EoW38kMAby1QxPiJ6+IPxH28oVp5Hx1IrdlDb+Y5RHsuedXEwBW1
Dj1uk4VbbcCMfaTbcVy3Fzhupnj+MAmPExVmqhb0qwXJ1BgQNCCStOeurmTkEAa7UOBrMwMUsZHc
fPr07KXYYDP63i2j8jbZcHhNcCU1A5gJSRembt8KENQCM/d/nXPXSU3ngfw+ln1G68KW8W5CRZde
qexsficDPfHyOExrgSaLMaBLI56biUBK/fYV0ha7KNaEWZVoGE4lRWvM9joNyHHvlsc9YrO6h/js
1gYOQV5NEOZR04tUqjKGj2vUoLLJRfNujWb+J9z4BJkV+C88ze8eYZuko3Fm1xUB3fou6AtCNRIR
+NP8y1X/JD+tH78083P57CcAOwDlXSeVAI8e88oyWpjGPVtZd49BTP1+WZMJspe6n7YCFuDo+yEc
xr/imgFLULYBMB1V5lsg35NoMn2XhHsyyQmLzQPJgITPJ+QwYrq17nPr3MzYcSQCursrZOAgmpfN
gTxopp2SwMTM/kXwMQxUpXB62pJoyMuALTOxXaWHltKDKsKWaHpofW5JECj8wg64/G0DF/zLCFg5
J4kbOw/sM48EfegfaBfg41gvLj0fmmoj1WJ9SqRHBECQpQSrCNXl9XKtWbQ6MOgFKXAgP3sW1IBr
YIQlrdrmcsiRzCGXvpHq5Wdl6faiGSUU3otrwWt55Ws72VwvO+jXwGLTG8JQGpHSQ5OH/5Fv4yHf
GMwX3T6fTO0quhVMnGJEWip9Q4qSx4KcTRBBLrZjPFRfcPLaniU81Eri5xeDfn0Y3FmMKmqrHoI4
5QdZHjqDdE1Eq4O7lTe/8tUnHs0ZmpMW2g1JfrrGweyvr9SChZN31AlB5u2jFiwHPlaoRbXMFgo/
9vttanvrxOSMQojHLShVGo/frI7uVuy12beafKw4LeiikFXgKcWFlOuevzS96HaBYL27wsJN+GNL
F1/Z8UOwwnxu+b0hgMfhtfE4u8bK0u3qkdG06qOXQSN+nluR8z9Q8Ct0rO91x0lHt1gXqVf708qQ
L7Zn5ziU0MXysXCWHdffJ8glf8z0oguqdBgwyWJJXOyYKBYzHCpMEgMfZtc06SLxjjg5b3CyHUJI
m1RwezB54Q8bCXIJ/P6dsgfw/q5lgC06Xc8jcqfRXD3NGWoeQTyYn9Xy2+eTIpq2f4Jx704YOJN0
yVQNFbjsIWm+hYetQIY//PzK5K/Ytfqoy1o2elE6YUslOGzZZLqnnYo4Qcup6E5rdBquFJxyuNEy
NVJ7XtdWvfVFZeKOqX555CahH6Ri0RKq7BeVqSJkxUnkDo+5dgapX7TTv7gxvAzQrTe6ARzqp2dr
a+iDKhtYmAVmd7/IVDN2fB+8mT0dCdwZGTyzNJ+W25o/Mi9t70HcKkCxkwSHnpD/3yTaWxJGlrDS
NKNaDuI9KiGcuE4I07gRMeZGBBFI6YKo+GOBivbZg73OAWOQw2p14Eyl/GOj31ON2ai+lySpxNmH
JxVaBLST24kedi6iaTeehaCBhfbjfpkkzBgkmpRooW5SmsLG/o30KeOxTEqPrxw6XQGx9i8cGkSx
np+uWIlfqZ7Pz428ZtUmQvqp2zQds58hY9ARv30Y7h1nqHa0i5uFkQDcMPA7Kat3E1is39cZDglT
9U0NzIs/r8zn08+hRxxugCYL33d9lKzemicIu5tSLfcaX4xAmcFE8qYsNHY8/g20pDHTxiZhzgZo
/CO7364dN6PNsceFfGNxfaCoXTWBeLvh2e/3AjvSv5Eo9DewDV0ALLwFlFXWfvCezw8g2aJVfBod
Ux8gTG8MZRKO64gd2l43n0MqE3f1qIL/oeXIy3Fkf/tBi1uWvEth/v6tWIkXVgKcuCEXRTiY+fqy
3jnmhm44Qc70GwLCHqxgmgj4aisOg5nAN1HKlAeAZAj117tAHluF+DKFxA9Qf85vMs8GT6F3Hoqs
2NJD4pwPRo2Ah4woz5pnrA/iIJVrTGYoJc3hB5K9n9kaUkemYHRqZgSxZ2EpNXx4BiLUq8AY4ILd
Mp5Yd6yOW2pafT9PcZ/wP5h4h1RkqmIxYADkSDm8oojI2lkOsbjkH0EuNn9Mz/B1QOTk37T46em6
vccknIuUShGapTc590EwfIL1AOwx3L2iHEG72voXfXSKqdxW14PF3dds7eDpgDZf2dGR16G736qs
xBXlcOC7IWkY/ngIYLCvTg9pRuldSqc5MPsymplMP93vtpb1DjfR+gMRyzQNDazF8NRn4NoQIqBv
2enM6OGycB/QIse60OnG+5jkaD/zf/CcHubxJcMckcPppEGqTNTNOCMtMlNw7IbJQRlHaIF7mzcu
BOnufVDALkn20bLhrOCX7a+dthigfxVVjgbHVC72stLFi4iYPeK4VSFH3HfLm++0d4l7PHDd6jKC
R47TUcx89E9Lc3rw02HovWG8X45HlaKQH5LIyZmVSkbEnXnNYyLc5qu5gJAzqg+m2mzV3D7gHLtS
fqIO71YYJPbrdX0SsnbmkPyGL//p4m3t5PAjZVetCPVD117ZAGQOMc/eZ61lsE8Hr+4nun3MlSdw
ZIZxjlFgyGRRcsnfwCPcVJ8p/4rASLh9ASzDFM8xPAV3ZB+os59E3oBs0x8xUcXk+s8ya82X2MaX
hX6A8g4LbkXkg6FUUe/4jCOWppCNnvDtwHB73V/eDsH1VKIH5DS4ydbQgbY8M0BMmZ5/bRUbgT0k
lkK8xDweLpd6eAHxBoi2F3ou23tr/WS0BodeEIL/qguNbuzlj9sOy4MK2x/u7n30qAuO/zWdyNZJ
4sBupyfsU/+QDERhl8Mc8N4XQEb8LV2u1pdRegSVqgR11sANL31ofz56uUrO9zduopl7b9+ulZmx
IyxMEKKRv08IkrDJQ6nrV9qLFauPtYe4B7TwhoMhDU8twt98YrDJQ/m5gA8EtPVbq4hYLKNYCdI8
mG9W9fXtkT9z0fhmeI0hzgIcMjut9djTC2LdBptbN6ncJm6xtwV4Zow47uXR88t/JEbGRuf0Q8Ui
k2uP0XifjITLPW0TG31kK+olenG27Nonezq45ioEWr2WR2zvocPpum0W+kqGHRJPx+Q4LqmpQqp4
HwrZiwilnjin/qoFnipoFgSe21xXDKFtM5bVAN6uWHiWHgIzjCdSVk059QNBxouFszqyGeSDroIF
xV5svHv66uxMuGUPL/RnvA2F/yd0Eo87qvCDt5brk169lyr8c9JBkjMY5kWIfE3KFV+gFmC9n5s7
mAeDUOYUD1S/7NDlpzz/6sMkD/KAtWHCgBCg2jpp/2pSkC8ncv4alMbqwdrIGgB99YGPR5HQ1GFQ
b3x0UDFMfusqFPKRE66YB8Zs2Pz1J/I36KQQa49KjaPsZ4GFIN8dgpQuIqOYFnmfjZqe30RpJBj9
A2iE+vNvwjUaQpi6mGLHnsufpg7iKzCVkodNqOcoROBy27wTuIXFteGHaDBdUNFXIZhfihQLHTMg
0eaCmg8GzvI5B4AdfrkGwg1hviijBSJkSo5dBN6aRhV+IN1v568wyBDfLmCOjf6mKGaqcPkNDuyo
SLvseEmiJKqq9oydLlw+/gBUrI4ywVkQzsiNWqvvMXLP1A2lXlq/9uHpqI4cePaV8n9RdV2PFnbC
j1+8OEyxRVCi+V7d0FUY43qdDrtF9QPqrDZHrbsRWsNHCJTjQNu+HqOS2u1mRyAzSVaIw+2q8azC
zPe7N/QYYxKr02UXOU5Q94400E3et+vwf9YhZJwxGtGSBl6mzOydZ7kYYl8PQKQDwdNQVATq8Sv/
4nVWwV5tpX8rkLnXBKrn/TCcI4MXpToz4EnY89FSsjGwjWpyRAbNdTuQm/gTAUc5i/a9KQU+fem/
83bWbXEcw3l921nO+IimAPkTC7HtkjwXxjbuGIlktPfrhePPTslDpWW6/ufrrYyf2HuCokngvtRW
IADYE2YzjdFPrgy9anOj85ERROq+WlfxSnaIt4awD986jCJywQL98cghalw5ynu/s68iurarl5VS
nUjnQZtR1zi3/bObHu0DqY58tmo+KottsRF9yvmw3o5ObIQFwz57oTmp7Cw8UtZui9ooQ4HIG2Ar
10fmvwT55+MdJvPVr09FEIQfNRskvmYOjPzpV4ND24pzE0YeUxb5CSMNM3H9mL99Zlf7zNbBCMws
oyl0lsKTCa/fMcMKSMz4hGBdaeuqg7Nh9SJJWWBivlIrQZwNoXoj8UjgN5gBB2wTaFc3ZHb6VBMj
Lq/TZrL8sXAluxuD2MXaaS2xOuOKsoFk9mTw8CEcYNV+T285V2FS5r+MeYmy959M+RmfeE6+KsEg
J8ZDA5bRfX+5vCpFzpQXWWddH7ggXh5gZRkC9NFicWi+mT2RROm91ewBusoH6b381+Ap5Uqi0sPY
AFd5AsjAbcXLPlHf02xilv6pdgsmRgjyGCinGeGsfTVf89hRJD2M/62V4YP1p4Ja2zXxKNRLp4pv
JoCFkkJDU/fLamUy7ylwa66cUDVG83mfNGGu6M2ojldCKU4j7jmte9+h3pPmrD9o1AU3P7Kqwcfz
TwrOTlb034eLRM8AdF7LRrGAdvCe0wD7TtItpWSCor00cioS5ezLgGIETtK1G1IpJwk+3UiDa7GT
OYOgCZUwh/OdMRjF3xJTkidbObvcO8eCwmM39obPorluRZwpuAqj2PA+98K5tkruzA8W/H9n7ZYW
u6GTtVWpNR7WIUB5o+vYFD+SktPyy/q5U4AM8l2fRa46uedN4p/jjQSUcJ6MwTsuUn/QRyftfVoU
QFyMigVxaLr5Om0NxNET1j4IeWLvbuSRNjDp55SqJPUE4oBnwmKgho9AR2WkE8l8UMplZKa5LsZx
Bh8e07ATqOEyqsdkGHUmLnWqao5xsg6tuo6KYqBQ0oht/8ty+iUxMIvK+VL9V3JC4/w11Idde/op
5W8XbwNJbphjXmiOkBAh5tMUK3ZZyt5MaBP8jRURkM8jwkC8WSzHA4nxjjrlBTC/iEglWPTpJBmO
N8NyidH7VGT4MUnIIDTZCTiYSkWCNVIrLBVDW6Hp3ReeoOfJXwLhs+xjykprIRSd/ucvS6+EBvDI
TRdek3qerrqz83cEgBHp8at/veUgk9JIB5o2xPtWBmaKWQq8o09M1ZUhzTKAF2jJ5wmtaBNv/JZ7
igo3b2mDLm3wdEkvlyP7wujxDJAQjbn3MtE7+LLAutw8ZRdv5IwoUMtIs4OH21GmaLt+PCrIKeuh
tqBnHimZbnXirCPLWFqL0KM9KF+XZbzLh+1FPMjjjCCma0MnMQNlvTsFcLBz9AsKiRvAAz/EEgCl
GlyRjgAxwqTwBqcExZXtp3YW3qj/f/WZUgiPhNWp3bb+1KjpYyJCCii8U1Ma/Wdio3NzE30q6x87
UCsdawnTwme0jcQYjoDV8cFPSBjTXZIXXKgW2Ah66hFcMNa1/EZMlIBuS/izudxQs+uaKUPqOM03
frJo7Qm4eDil8XwG1bJ9wX625a9mMexlPCQN3xv0hiP4KN+dM/6JPy62LxHQSBsBQXlYbbDpzmUE
OAiSzkRREuUe0OB42ei3aiTddoYF4sZTAUc0MLwYxtQhaCRYr7jPFDDn7E8gwOK6RFwAIwlb0tE4
FVNr/84oBA++TbbyB6oB2xZAXR/yEZivkKp4uoYU9FBu+NBePsuPEEnVlPt7aC56nO9K7ht9bWDq
qr4Xkh5OR4CpJwQ6j9YWZh+U9VCWOIAqajmVEPnIjecwr0HXyNrPXckAqKY11fsE0DFpF6fsBl2R
C7XdNZxtbE0G4kCxm9P62Pgla2JcEIANg1ypLNIprdjyoqLRVszjh11yqK/gWgr74wJOM8OKwxgo
SOnKfx28G0mKMB8lFqRzKoBLLR8/JvXs8imhE1BT+/q8dWSuYBZF4stx0Y8mX2UNZ9rxymCKv8uN
Lw7bnAskqWXZnuiT8Qa1fgey1P+BQtuTk8zJAOqZY2RCr7kfoyt/C1cj/JA5sry/lpjtPppbExK8
xJwhL7rMDAASRT3Krb6Gvjy2dMq6azf5bk7Sf+Nu1+kX3xltT0PtpsFiEzCof0WbjCIyQ52ZuPTD
QuZOQRddWrUMQcUMhfx9tXSwrPrZOzsc7VYXorAoQGZ6P3lSJCiIlRv6XwsVBa182JI5vkn0qyfR
I9u9IvxJsHjMEdZDbGnMhwkKYxF6VOywZtoPL9EJCiEjomgST4JMHJLlbrs16GEkgvPEcaIRwpnw
SqyO1lIxDA1Qgepdz81ndYERC+Uvr3mW85qKAnNn8nUdyhTefB4OFkwQGadRN4vUnbgm5R2PH4Je
uF9Sjnlv49SYXmTCblJVFygdElCa1xZYZE8x7SbDTPvwQi9iqyDnUrWfoXWn0E36JJIdghBzMFVa
9FUpzMw7FTJM9z1qWw0w9uwDQhCgQpwdUjWU5ME4/dTfCGn6/SKjZk4dWkc8WJBocozlrJ1lQhoZ
Rp7FKIFqPwBXhaXjzQEn+vU2Hr0kdrJBRqbYosfDrQWdxR3OLwMO9eICU0Qv4dxealevxYFa+/Q7
DzT58vrGGxc77n3FGk5V1AtxsV659XYoyGPZ+VAoecc+LSGzipivJfeAykQi+ohKaK87g9AWevpO
hHY2cojY7k6AqDE9lcrpm53S6aBWEIUvZiAhx7H6zlNQ4tUDfIFy9ZNCPSp4z76ZA1CTuiQOjFp3
NxKLrEfetDQh8QaSPHewDr5z95G0EsBFhW0b8KaRFIHrrxfCz72yt3VCVumReZMRJjZ5qrEe5iei
e8Bs70z9aPHHTg7eNa8fblEWvBjLYj7uO+ZYQyW6MCgUQOx6SmClRDbjT1RBYBa2Klq9Rvv6fZnx
WNDzoKjlMP6LDZMu7QyuWXE3LsaAzAjfQX1rdTFi1Uz3NcjCJKAps2GxzbKPylhGVsxgJFCLnllJ
ftkA/yySZogAeVLoQfu89zmq/cr0WXda/xBxa8VJ2/NUO1nF4ukmtyBh+PUujPAYK6Abzja7XmFO
hLRvztZxh2NaBdagLQyrUCcP+ycETk7XojppveGrT9M9ihHbPxM26k4e6lc/ssVRP+itohw6Ze0Q
iW2WD3EwCWvrgX/80qQwqVK+bQ6E3TsNhnZ9J4W+lsTic0/eDMMglIZ4buEDy8Ozd6vxuM2rga+4
2LsIIvQt0SCNhIQvbf0m00QknbR6yzs2twgT9SKsrpFfCwYizEp2EBS7kaQevrZLzM0vTE754zCd
bOcKGaF68ED0QuoewOMgm50rDJrgsK/nRR7Y8dt1dfxNds/yR3sP+jUu6NiGVenyMoiCEdZgWNBq
rA1k0EVhWw5bh1npjXPoox6DieHq51uAL42XqICsFy8a3IUn3bt5D0MWZYFr9n2ABUcQiI12r4pG
qaLbogSeoGoQIIQ4t2bScNIE/HSxdJeJJWLQvkyfI6b7ZnnXDUiadTP8fTohrUbiJ7aq6mwKpi1W
QLWvIE4XbsrqI7nAqA/DpWcLfd1lFEe0N4yYw4QLXs4KNGq1Fn8/GlpLlPY2wVP3FELwqgTs/mvy
mD2Z7cXLSnuTwLVaeGhWSYmdtEfRDqRpc0PVcgCXLI14zH0PrOS154xQrEGO35ZedwiA+h/wVQPc
upoyIMBWdUfkjH/hg5Lu54v6neYyabif9MFQj4Bjl//3fYrKdH4dY3KW3Izn2Z94eAWC0dOlk7TR
W4xkDxk/q/DdCqEWYwQQqSFQGwMsyLsbRZ6ECBSDHzaDUJKR5Jh9c+yODr54VRqKF6JKGhFZXX4u
UzKEKR3N3kyRcxeRBB7AvtlM7wJVSKXCO7aXaiqSDfLS+bocr5fcUZThpEI49319FzRcYGuoZlfo
73iD8z1tws/kL5VzG4twYgZ75gndExuQkjLDGedUtu2JdVgr+ClOylg38ZmD15c3Jz6M/fWueL+J
++OHCM70sipshh0S3ouAj/ZZdkcMhbCctVKruHJpcn7OaXBPqqCdSTyV4RWeNE0EZg1XAHs3oKJZ
FPCMCU3pRS+hZZi9N7gCZN2A13YKUYdKfla934iXpkMiI+ETX/bWHUYgSAEh9zfeGj0/w6gCRA2e
ZlzNPqUvgOGAXAC3iIODbrkRyy7MvFUwxmwGIkc80kjS2ttV7aOvaIFLn4EKVDGlaoF0O+D3XiVc
XTZzsuYnUM+dPFGrIcZAMWgJ9CRp4UNq9GU3DVoWSEgEYYlrufjs7fhEJTwnEGqex5dvZvT/Ftmc
XNB1ciKcjO8u1YcRirN5cZqdgXKpAtRbIMLzfcoM9SjJtTZ/zO3Owh6hShpngXGlppnv4Mqt/VuJ
evzR2t4w9UpOn1eMIB/kBvyYlIIFZdd24oa4KyeU68p+IDI+pzSqDVaRbdRcGuoM92Vjd2ItXfV6
yjx4HVY1l+ShFe7luim7t42dv1xK/td234PMiq149b+c3BzwYyuD5ZgCOAJnXBgjZNRMt/bQve9T
0kM4sKP6UCN1jaLpS1Oc769ZDGFqcmELix/Zc03iUQPaffV5ccbaRuZJKwP/AbmIEuWjLTkV4ihB
+k01RiGrwVegoSfiC/9e3633Bnsemhx+RqnmCRg/OsDZ9NOIR+YMGipb+C/KxDbxAO5PsNK1Inqj
gsFQBHQA1TpwDRhSGGlSuxkkAxoi6HClsMIebJqkIbdRmzyWChQAkeWtXWbj6aI8cGSpfEig6/K2
rtme1ucviBqJmg5/8DW+l6tQG3kB560FrGwTgxskwr+1Y/ZTw0gzWii1Yto3B3c+95QfNCMm/Pd8
DE8Vo5k8LziGZdnGRKTHTShiZr98WeUrHFDuWKx/8n6M+V6R9D8kga2dRleb33eU5B69kRBUGtui
Kcvay3fiQ19xqySnTiPE9lqjKvEL78oL08TAe5paJYGj2USY3rR7idsCIdfdCrkuzf5nmC7XYTP7
ZKKHabmBNuoBbGQvh1JJBa9mrekHGo9Ikkc36n4Ha8uSYUCfBSS4GEbRR9kRbXRX4hWIq+9lxgX6
3YHnJ+fSsJBIaQ9gkWiUu7FH3Tjxc2IEtjhFVxYyo6wnPkNu2KADbsB3eYlHa59FPvxjackeqQ27
wMm5SSZTdoQ2SSwdzBb5loQdZqIo5PSw+Nqqb1AZEFWs/kDFtV/77Nzw4tkPX8IH7/Rh/AKlje4j
PePWQ9anSVDXBnTniIijgofXVuUklymblGW11lv9vbHfswh3xUr2KpQlKisGGeYRZn+bkDO+/Fh8
4ytnXJSyXtZueEIYq65bL5b0FEY1YLwPsyoInaBauL3GMQQV3e4NTUvgA4ErfLQp4OyoaMqTTxAI
G6QHvvcZ7o020K/36ebw8JGk+sb5+mKeIFlKPGPj6Fe+1BjBFgaEEgeN7nh9soc9g/+bPTccLXVB
VoMCTBPqqAD1CXHwcfGLqrFt4K44ThBvj83gw//t1wSqqLDYdEpCp3bwWEbazXY3u+YssIlutTd3
M25hhHi3W56+IBGxCjqoqgegRIyAqgP+1zCRjc2jTnsMiOA+DMkhly1WCkZGQt+w5boOsetDObbs
b8r8PEbUcfJErurS/9MY/woUIQrt6Xm7xFQgMwiOiV+CNRXwclgj2GwCW0YAlmMfsz77LlQJ1UvR
X7JAZFl1Yy0P6oZHLyMkEqgwTFzuSq/F+vVy1E83sV8T177/8uM7W07YoH/TwQGGVmcqQ4ex0f+d
dO/j0Cd0JxiewwoH8MZx8msfGP57MmgiNQkgyOMCSIA9AJeLtwgyfPrpEKez0dK2XSV9QD8dQ+N/
mr5i3HaPOFl6lky4WD1mlp2S5EGmc/0+APDbjzk9Ce00iHFdcWrvPNsT6eOnuUZ+/QBInXi87/b1
J2riyFZ/qi7Csxfm0ZuV7nLfQqf4CtukXapPk9vcGEKJnW/vP3/JuT7j+jR2CLT/tX0OZULMO0of
XTsvAUUKTydr/Rb44AodmpYc1AjVZORi35T1ktInND5+67wjIrS2v7voT3ym7J/5v+iQ/4gqamxm
Y/ntPl+/CfDpX/Sg6jG6yC5+EQgKTEvUU0u9n+xcSU3RJ4/d560HPXAVtNR5JOaReu9u3cWDClHW
NC9pRHx+JJJ6SHl1Svx+LXOAEEu06hFWD2rdxVbn/viulYwpKYle80zVdETwVBU2UGRLPaFBBBFL
Nqqb2xuQBIex8etqLPMQW1AMHtRLT5alTkplzsTD+ApeKJioLDQ+wIJXsUu21iqSt2FcYoGVWNw5
BGfaqj4PMY6srJq0df7jNSmihK8AW7aBjrsFBDMbFgKWQ9yN7uA17aBgbNmXHB/x0PbWtZeHICZW
pMbt8RnVZo/KmRkvB5uaQoP4ZdnYalprFSgjYhH2EgFH0ylKyz47OvbzDQ2/KxNgDZiyAt4sJHEF
hx7rwleMveNgOeHf6+B9fVk5/JjwqB7Ej6I7aM1pNOxTYyEwnVVPfBPJFEu0DiaVhKDCqyzd7U3b
SH3ofWvDtV9pnyXgfFCFrtKBIjTeE1ww4d+vsVPPHdVaqxTKkUxZnpcu8b++nXey/4nvSS1w56fa
lP9UlulwCkhmlp+9LstDdbo05WL2FdMkFbBVmtQvZBAaVWxC9wGZ8WaIkzYYYNLQmlLSPbyy6e+f
glsF8sHfRD7yNiRHMoq0o9/40yK0wxRvetT+2e1uSX9et10s2anyq9sUhBXl4zuOQHPHRshCGVkH
DfTLHtRQq9h4QbOKO2Fi2TFg0RAKm5RrJ7TFE6zMH58mYp+OiZxjHVJlew7Qhf44CHwwjCa6L2Yl
XYRdutxKkLin13aofrXmlqJyE8u5N0fbDQsweYft2PvJm1CdUMJEH8RXG8sc5YrpkzdhmLu07mYC
Qcfq65/PocOW/QZ8xLNq39hNcExKICI5ODbrEQGzElo1niJVF9ge6v+E1/t2f7RHu9S2zdvnQsTi
BzuUc1cLHwd3gehZQ7ZPTdP0rsGe4e+vr8plxCdLeV7+rJA8c4Y6eQVxdpQkQWdq3hPqGg1n3iR6
e1bf+v9geKZ2o86I5zzo3xWEy8o6i8uc7W/TuXdsI3oN8e6U1DOEMZN275M1mzYIqqPcaba9rpD8
ETAIxzJHv9yCNAP2NRZoJMDvj+P8hyX2lVlTLl5yeqHoIDtL9ZnDnfhTnbLbv5afvrW/m8WRk5Rq
XOBQ5k5fBxrxaAGF5am8Kq38Ul4WBshJUVTv5FtJXPJRPnd/tm4Xm0R6Yqot+EPNsK38K9JKUG0v
p+MvseFiBNcR8LUKvbsMvYwZq9HhAUNYOWSdZFPmuZBh4GMojUwR0GIrewRdi2K53dJehh25L4Dz
j10gfmIaKK090Xu1v/pJktAuHOp5OCvk8c+9JOkqmCg+T6ivmAsnrQNbz8x2WzvOLAhBkeG3SIaO
nRQZNMj5Qe+24W8+XlJKsQnzWVN7OoWI09tB8NAQCXGQc+PfKyS3eE/GqQ/J2NeIzWdGuljjtYSS
Mrx7LjKfv0Eu4lu5ObIUyeSUp9p8275ZvHCjVq2/fOmAEOk7SbW20NGvtCCVBhiVl8H7gA7rnc92
Dbd1Djc175bFoZ+D7Uv2xNsdOSotpzEC9ZK0Q5dqvlBCrCHg6DmbjWULxUVlYFlbm/MnfcHx8dOo
e4O7ZLA1wQ0Iv8tT7Z9BXDVFKhRYUCOqQYPFXMZKsI5wdNMLkQ5NxPzY9RgJozhfSt9A8w7lPC5I
B8awwRhEo8lBKNVNx/U76255KO4zBKhgjrsvZwEj14hQGN0ANjPr7Q6w0doo+hrSZ+0AdUChCVjZ
rRN4RxvH5l2IPlgC9yteTRYheAM4WEzxAWM1O6VaHnG5hYw9QhWTmsJBvJehWx++w9jk+BFbV58j
FPCqajoprVJvPEsa5rSMRGrmAKEggtYq/BAy7y5ki7403hWK+rR8twYjanq6Oe0Req0Ao2OJcJm/
+bvnGWHRfcyrlQMnziV9Gj5nF9LyEfwC9oNEu5NqgQf5ZuLvSvtlaOFdf4Q+vpTuX1vtUB6QdrGC
wVoq6GpxCrB7tQ6UVC5IrftJ0r/XirLLm99jaPLs1B+NU/Tzkv7ulpmqQ5OicVVJiNE+OxbeKk/m
24p5p1gB1bVucbofPxLulI6sZbu7QgA/mTpkEktKIFDja+oQLIxRKx5RqSjrebKb12RqYgIY8IJf
djJkN4UtCez/gDxyHpuAm85c+V0MS5cAy7pAwlN89QNnxLsIt3LWSAtlyYW7/TsF3V3kNK2WN0YQ
tZkGokMUGFUWWTbdVQDpO9pbhKx/UJGbyf/9EBSKkaLT9l6KK7ZgcOm2M9VyX7FtmQJqvNBhsUoX
l7MNvZmzYmlbAIj5O8Suj5Ze8ABh7dQzWwGH16dIt6cCMgfLX5a/3HX3Mtq3cu1jTCBjEkMxHJUX
Ps1vPeTvGWv9eFLVawKLYignN7/fmrQIIBCJegRDwqECPxgUEkPGHELwBWuCdzOwC8FWcm6HREW4
nJCTIx5dXuAX4e3csd6CIRWvzmzYY+kXjSv8VG+tjhROSb5bHS833lqsefpA4c610m30Lpz32aKY
W/YsqOTOliV0uegnRFyINDxUclKj2NorJF7rUnEEbg+VF3t/KcFZDOlg3Y4+QRyy//SXdFjBAMlV
TTGAJR37FkNTIsGCTTp43dbfU9+PFrclko8yFIagaA7dWY4UerWoTi2lKiN1rYmQF1+lwrZpAYsS
kGKwvqmxmng2S7xTrv/j5P5hy7ZRweS4HckVwUBZQ+Lr4Gvbv/D0RHXnlT/US2SNkzoM8wayngG0
v56daFGIGhycT7VEEJlmACVk+ZK8T8yvmL2+l7nJ0TjzVsh8AFdUW+mursbZ+ZRug5VfPg7X3inz
Ks9RdUiCsJTavRBusfjsTstWN9kH4Yj5m7NNljSsVCm5SM7Ovy/G9kg3lAntkeNAfK3vnJp/TKqa
7vAaXBv9kmYv/XIY6QO1B9jJo6+sIEigfDxce/e1VIdxXjVZ+GCIiWhaTk22m0G/ilb60pHNb3UD
mtC/dMvfW+W96fjPDf/0mc7Pt9PSMtyqKVlHxCu2CwrFaWJijapXj7D4WR7bO1d8T6C/+tMEf8gT
9loEmNu/fyM7LgLBPcVpRJpJx4Db3VyqCs7hpH0gJvbaNsEhL+/MqZcmBBumBq/L1svo97Us3IXT
W7/GAuzNqGrh/yqgQp3Rbv3PM0npHC1xaf2Yo5wXY/tSIyT2TZ61Omq5NH8sYWzAhw67WvjXE4xr
/PL01Pz/AZHTl6/LyoD05cMpKUvhZqltVfH7migLcxJC1cVD6Ybz0l5A6VE/wQB+3cS1uWidX26m
c7+n0ngbH74O8Oc4VzHK60HkzNXyqLn1qDfj7ocZp72N3i7fubWUZXbq1kVzviJKoUJlN2P7fLhQ
Tme4V/n/d9X1ACYeS9hmLNIKfURsHnAzhlecEm4PHU8AOZrOxLD8kSemWuqc3zQF4SUlLJA7/5pk
zDIgPWWtBSbxNDV3/LE2goLY0L9vScnsSuly9sebjFcDq7Kgkdym81WkKuL9mTGXowGJZd2CRyru
In7vUt6h0SQvQLTx/e3vb+QejEmkxxf5aeB1VNvb5y47sEFQXmjoWj1fyYv9oPk9BKHuBSkcUcnR
Mf3/m4jfbSUiABzCHaYZ9pOavUiRSeDmwItQdWhaCDdL92mXN0ThMCsFVLRXYhVPZKF6HHLa0e3i
ssZFXyuc7B2J1dfHCeGxfKzaNW/293bM1U1kcGVOdYdCpwcpWva5BwEv4WfIBXys766dLgNE76nM
Sp/o/NJqzAuUubzMyrKuiJryTdeNZomUf95ZkYiFNm/xbP4gKfKIuq4VpE8Q2x3hVMq2C2c1LnHG
pFfyZao1x3fHrdneTfck0JcnBa5ZY9X+1Aj4g6Gv9xx4BIMhc3eqDseNDcZN0NtPKCUISYjKTV7C
tUuBSj+256rCj9ZdgrBD+Cg2eq1sZKtEmh2wNq5feNjsEX1AvdUAyjLQhFsMFvkvHPE5i60J91vG
eRuvAnNZaYOWwzWa3+ieWp2iiIvJf6l9G7/HhLVMf8HpDxLP+0B1Sg/SeCv3P8Xl7Axd5HOSE4rj
omO5nBNb0oUZB0owednYKkoGUzd8CKUYwX5VeJgHWZRtCWUXQdQ98P+oi4nE0PPevNaQsUVema8d
YjPMG6OZmDyNR4S3F3tEwo9LOgYhv7hVPtkYhWPGGQW8Y2yqtGNEeNqH98cyjpeJeTzKw15pbQqQ
/2/DwKme3nHohQRvJ8HK75sMK3mTBUxz78w7sjS1cfzz7TfLvl0+WH52JFGvp0k1rS/Ht9zx+vM8
q1wXgVmtXcUZ7DZGTew6ySuNUjVbzKriZ1tgWIl92cJlKsffAu0dhHCrENDv+D/IgvqYxhZ6dYcQ
jzMs4sTqcLYgs6QhX/aTgMahsCpBsDBg25TITwjuIP2jza2kvJIsgX8nf47dCFN6VVErVXoc1Ept
Crd1BNzsFjlS2YA+kUQd6tmKBqUNxtFj7WvefRB101LKSIfyfmDSwHP/p4iSa8ZVbf2J6/CbMA4e
jP0v663ywB+/0nTMzhETMmvEiKeAenMLDT5ViV1c2ANolT5ZKMWwgP0IG3aa0dfAEdQ8osiFM8hM
3qQY2GUtkG+I4Ky3fMww078Lmq/NrfH53iAnwHgSBEiMCKUDkomulCTOc3k+aZof0yDzLb7vozxN
3rA5BZL/gxybcJz7nYvkRaCotYoDiwFjm4qhWpcU8RbJllzCnSqi2QrttErVtEWQM6YTNHtwZHMu
OkWEM0hQ48HICgk2H4uD7mtKTt/XIVMzRgnTflchN4Lo00d6gvPVZC5LDzCq5SsQ6YkW99pApjKb
ibKEwF/JMEkdst7nMKxLGDY50jmS3sYGyUYBE7KL4M916U8UgxU3iuI4P5+kVoiS1d7QPL+aeP2B
2bIS7m2+0ndnIqJJNPC9yRWaJ/ikfao2XtAkMhuagyg1YAoEidAosybJQ+CLGdyl9GM3JKC3s9Co
vOsNmZbOb0C3+gkbXdfmlADXMRVBhmJy1yKyuu4fDjitrZWFr/PV7yoQTEfBQgF87xOTI1q7qnn7
U5z7B+zb7L2kAISfQ13JIyZhBwQFEhFDQexR7nn/aTEv8KYpwURochxNVM2RCji/FzOao1ldVZB0
1AqRqpj4hhO95UmQmXzQq4AGw5IbXZBu3ss6q8yKQrhS6RYesntj7VwayR5QYpcHld59rqQln/Tu
R8WlX15khgUeV45YjJnqE+gHDyNw7+5u7PIMjOduIi5+xV1Lo4vAYz+W051+bo5AuRsvkEk/yaTc
RI7HUHVGUIGJWPfes5P+gGHoZ6it/eowF3oZsI9cbxAXvJMnn1h+PtWSHw+YeNSlSTI6+bAkWFNu
4CEj58GrFPJ9Vz1VK3LpmZir4dxcaA7ak5Y4L8aRS0SxysMcjUjHGm4xCjFUdBjE0yS2qCuCpVVT
DkTQ8TbHPDz1r33oiutJ9kt8t5N51JjctHF7qqo4iqIFu+epUxWtBVJNP4cSz6zBnb1ZqoC3kHkg
BzVywDVw1fOv5cVQi69FvTZSYCPaPaH27FWor/BzyOwUHdk2YNg2OdkMaHLLzgJ1mOYCLR2mx17c
ML0muKh30TqZjbDg0i8HXZaxntqSQAXmoAY9yOTTnCFf/iwCSSkwyOf1ibQ9PF2fN4S1nvlqDX+R
mzyy4we2oa+G5IakK2Ht4R35oSH6Uw1BkS9/WsBM1VltXTR9hapdfg94qrnN4R2xj/8zUro5oSE2
b1PLI/UWSCP2wx1fBiQ+OgRGeSoIMyx7sAALNT6IEzU9qlQtiU9PfBC8LM/P/jpzDHkiTsVrzUWx
ZtGo7Vjp/bVeng/ARLUeiaaKgphMXPrqPyC5rrORAaemRfstPRdnA+gJMcfD15iewv8Ldc2lF4S5
mJdrvZN0MYO00WvLG3NriCy7fsr0m9MGz95CxUC4lgbbRjWMJY1IOFvWMwj8Dv48ny3paTV6kU/I
eSRYrTk7XIy5qxnJkMiUYvzQs0yB0oikh158xODZ+zYD3vfYuc4bqA22D4QDZKyvx9MXVN9AKH1l
3Nz2YYzTu+emP53WVPJR+MBkveEK61mKn3FPtprBWbI626R/SBQVQrCq5nCzjVUi/pBA01U5uiQO
RssrqaJa8j7wh4ygg0wBDwlBlH373aWSubC0K0NdhjulHE1udoQi7zsBpInHoog5fnQv4J5Q0Wv8
0DRg5lKBAJSQ7DZzjQNV6wKE6kGlboQHYihLtrULEx4oSWVnP5l/7w/niov30R/Toz/Q/kzt0Kpl
oB+IWdiKhvfwplYPd6CqQb+XacOZiAp9uJY87X5CFMcocp0b4GNZOC3GluFKQ3Abk4kz+eGgnojb
FNcWZaAU8fTruJaB/t+g4wIEFB43u+pZQykfjWS+arlD8SjCgcTdilVs7YJZCcMftBBqO3x0jzgX
6HjNTKifx/pAigy+kYgnaNMKjIppgVVeCSszivqsOWHy557kyjj5ho8LS1qHATjNygS+jR7vjaZ2
vvCjp0El2ls8UaAyo57hFsfRJGJ9V9JGCqkyQ8pCaw3YIZtEQ3y7wARof4IRSUOqr8Sdpg2rh7Qt
govye1JvaNUVEU6GCPehLsJUIxIja2lFmSyWsf0FfEcR69ef5UCDc9qVpZq1EM3b9AiAOAdTOLrw
nV3pZVRQrZgSRfniZM2qkfAqnCjshRuDYn4/SGjYEG7CPj1li5nPlIRbwa/CVoWZ457T8RfTRLnO
aPP7eBP4GYGg0YclGa0N5IggZgbyu8WRLbXITc9Jwnt0xrOIucTuRxfCI1MbIf/OJzpI4GAirMiY
IEFunLimsU6wUG04EiZk1aUP0RqOiMkXL9FEKE/f96BTsW3uaHZCID+P7wpoWBrMWJXZwy7CyNjI
iQzhDAXU06tN3NtGStDEYzDMCOxRExDleysLDiN6EDbPDE728MG1rjRhWLxh+C4uu+X1p6G6uiyp
oPX75ql6038kroz1wd5J9VgP67u2OCRZit4XMg1u3KZ7QYM0LaQAe4EpQmaggAdWA354LJ+ioNL4
53fmYkFvWOMfsF1P3ip3D7s7cum14owSGlv2+zDp5FWsaDaqNj0iqhfAW1X34mIqkkAoH8geaZsl
S0qj4MYmh3nVuRwD3dxT9/lNnAalHSeE2Lo0coVsgzbdZNosJixGPjYtFqnCIht9BOyHQQgapKC3
g96KHPBuAsgjEkCQ4DjxKXlq7Z6QeeeoXZQI1ntTkgwvE0OsIpZV0F67uuuYj+mw5bmzD+9pGOdp
D4LhgOyu5UjLEZ8SmgGJv4AG9P01vCc9Cm2O+BI2sHh2JOg5Fisw7cz8nVYbeP06TNgr5cjtlLUM
rH3/VHsPdlolrqujaPj3sPE0vsStjAzszMJPmg0q8fIWTrMudnHFLaYB22A3zIajBDM82JX+3xKb
e0AosvjcmbCqg6SIu7p8FByNLb228nbK+7+TbkL0+WuBMOYc6jVTHDq6U6QVi3XcZWz1L4+uTN7/
GtY3pKor25Wkm9zuhoi4LWOX1JBvbfJWtJgtFLSVPLfRHlq+27ZR+rQtiCgQggC8qKvWyvI/yeVK
+eZksNytGeI+NqGg3yCm2C9FIk/Xwa7c8L1m2LbDVCZiY0xSTbDKOOcg9gkQqJxB5WbN8mfXsLI9
vHqvHcVFD1OSa4ac1X8X6EsiyBrnhe6TO0cC42yv6C7rSjWoXhLC1xhuEUhYjd47ohW4ZNIr/f2k
IgagBb6KcrOrvAPO73m1q8YyU5NJJGshIj1AxYglvXHei59mspH+GQ+A8mJCK+qR3fcdUGfClYRD
cYJGPFBUcrQ4J7xXWT3AvlE6ZfxjNQA7l+P+/N17+WQD6iAB8+IMcLGT8aPPwB48wyFICp9wZlOr
xbgm7qZ1zNEaksoMIvgsGdZifvrf7UD/iJlbB46RJvslmsUAUi9mJfIGIACdfbt5ObsIICWhHlsY
qaIqcBWkFlgNxgWSUE924ppT1J0/NN9RT6KxaC3hBFcJIpiIio6lQHl/AdOKD9Pkr6ymf68nQqZU
2Z4bjL2orAkSUMck70IyGdn8879vIlt0PsIy7AbPAHQ41OQgFsRaGJEpXhWPBqrZcvjPRaKF+Av7
TnV5j1NIxDpgmEFbVSgVLXX53DtInM/C4nRlMiScDzHoCLeaSyRUvcBpFFAaEcC8Qt3vGoLfRkG/
L+/PXJjmY5IizO/np6PAeUrpKr2NwGTpcQHfAKKiLVfnReQXZzY21wPenhOONEaE7QXyCipQBwAt
AG+CE1oIhi5uZqFDGbnTIEBwIrQ+MK99ExtTWRspQtp0huyC/o5No/pEZFGO5fnBFlDWzBcqpo6/
mF9kxL0ma/tGoFJue2MmlrYi39ErS1QuHifjzArKlWC97d7mlMEtfF25Ic6ibxQ0AntNszblgukV
IBcLxUeVWRO8IvStM1HThJN+6ZXoHp50Kn2v/nIL6hSBlL0akRgMX/LSh9MfLnsAHVkO2EvTP4Iu
vlJmBvcHAFl2VKGKv6HS/7llX4bMWlRmUbv+oKL13gEtr19q7z7ajWv19P1A4AdRU9yryTsQhRDp
EY9cXkQWt6JjvPm5ovHPPBURUguDM7r+e4hAJ6w4SnbOMSyZEEC0AvMLe5e1LmkXILiVKqDX4s0e
kD8DAVSwDuxUVilfKdTAHymIfqrXZJYDk8MPgaqJYsnm1+cp6Ntma3+5qz7qSDWPYZImY4+BtlvH
Xp/EZBd0vnUUVpsfV0e0m+d/QfyEf9+5TwBVNSFE/RxPFVqN0V64z9B94zqJceazJL4xTfUkQuo1
4uOCQxbbXedwlQAekuO/m881nQIxBTbNwOwbJm7QIFh1mqWZo8Rwz33o2wXWF1BSPhq3rVaNyaKJ
0m7sH9jsLVOLnvvSNH7c9s211o8n+a3AuguR/GbRJZvSKb8u/e8wtMa3K7HVP4LIz9LZwOY0prdu
El6s0z9KitUu9LDzx6kYmP9R0Wx8/pSkW2BRsl3oHFGkhZid3aiXo3ovPrB7WojNiKckWn7FhIar
QDtsQbgVflnlqQGf9/qYfSQ/oXFduYLzpBDDV9mnn8CGHSzHIq43mGzRo/54VIKGmE9Tqv+ax79E
mT14uUtG9x/AL/6kSfAgxkLHqbXp/BHAEn+u8IOUuTOtFiF4EgwtQJqaFyTbG/IHJZtXBBjIHuBG
+gXuDwhDrAMRZoHn76SiodBVXJNkml5G5hgwuprVsAipl1defKd2a2MDY7WeYwDUsopd6YDq9yI9
WdB6/KNIj7Kqva6lDKuxdB+Fk0HoXAeVSLEtDgYv96hCARhLWgf4HkFBF5rW8lHctvDrcX2It75Q
TtRvQvf1QLefQ0aEbKPzQ7olvyyeiNrYw0uGnyMi3F+qkvnCrHASZzMosL/f+A6tAl4hlHcgtgXQ
KWq09jUFihwff0N0falK1zDrJm+piKynVLRx1v+n0euJ9GqT6acXOPsTGvrU0E+aIA6arQlH16KS
ZW+6LOJOJJeavDAMk2YJ39zfoJUtB+JeWW068kWM8PZj8W4hWtmV1CTUwS3j835XqoTrD5DuYGaf
SdeXSQeZvHb/SNIWmLlRTj0XXRFNp6qCCe9Le2lSKw8eptaHhWKJaoAG8Y8ZY0Fse1T3oQlYGg+N
P/8GVB0dQh9jLp1g3KSCVoxTbeAl8AT2lqBkorzAJLSarbKs3FqQldLtfnT8B2ZuPWmbZV6dBMIq
6G1W1W0AVxRVL8/yiANOTvFMyx0blTMfllycYyY6uoFOwHuz4JZV1gA96n4bgnrnAM7xUDhaXl98
qCUXvnnd0Z/pIhQvu6+SA9mqZsvp23NY5v5xL7eE7GxthhQF218AJB0Vs2bcedTvkVBlSL4T9cqu
42TFUIK/72+bxH3r8bY4nh2iDzRWlqLvZkUBsfAi0//2zVniHZIhy4ful9DeU+dPh/XfX1oFIgIg
FmqPhVwmu3uLerV+AFjgodDjuiwDDzFYVHuLZOuc8SNZKXa7S0V53LPIzhfoKHWcvLU6D8uVEhgO
qCgarSx4d82CqL+gB1Rnrbhd6vzCZQ5ygQonI5vJXIE7d4nkt2OYQiUeKZ6mPP+gE8iwPrd9tv7E
Bu6d6IOsQdrWyzYBkWfD0RLyDH22sD/Pr/Wg/EI6iSaAkOWc6S6oIononQJOdvNMq4zvuQTlfUXz
t48y07RfGMWXdmuFTv7LVqiUf2RbNaJYgn5vMkofuDtLrVTjzGuL3L2DbtoZYWD0woFeOJqEBVxP
IPlv5ZteaYKqNlr/uSCvz0WFNpWb64BpTixNTY9L1l7IAEtkwVrrraeXpldlHenEgSoqPVybXUB3
4Z30iA0/CJphjiFn2zt0Oec5swKqTsP45G96Hbx3xzQwfYNlPHd9S2fhzR1fkBEf0NzItM9cxFMK
KoX9dqi4bhmyvYx9bvnpxQvGAXm3HAhxWPJnOrtm7/QArHEO7vV5686f7UJWeie9bnGPkfCNSGe1
JZMPs3uY9hey/sRQt0KQLScpthHBa3+p1ZZSgneiug0mvnMu5LkwtP8U0kgcO9OHegaEp3ICoKjI
7zgHYtb+B+ep4YtSqPlZUkzzrhcJxn4dj8IDdbHECcKJyDF02RpAqClexS+ITIjPvIcxIBFLlT9d
K+Ggs5gqnszJQqFwa8+RRnkA3DEK/iusbowM9okvURGVHyhaorlfybPXapWyzCxAe+TJ0KFtERVr
S6QOLVuXpXCqgZdWbqTUd2TmkTXUelM73W2iiubW1TMPtQeN+mo0RjHgd+knVYzeI/iWbRr5c1iD
7CcRhkSmsMGMzNAvsSCp2koYV0IUauy5h1sEzXRYsUZU+J6sRHApPX55G5I7XIHY9xBsCIn4IK1O
sYeuRuYr9VrZLlo/xzH6+aIoBx4MZY2sTFWy8lMw9KDGOSrwF/voLTxwJYqihoI9y4iRlQuZJhcC
pVL/NLOgtP4qwygkvSmALWi7aefuGoyxN/OLSt7oasqT586FeUbW3XBiXoIrwYP3BUkrXt00VXK6
bKwd1iHG4CkrWCZijrc5erVnLsJuJv8+P0VluQ9XRBAs2aZ/myEiR5FOgN+dlZQmcr8zw1CGXpqu
OVAZItw3AUYTUIsgryhESpUmBCFGDCH5um55HX9TP3tzDlyVJGB4p1tH1R+bH0MlBXUlkxTv7Me6
QAPob5uOnDa2okzCKZeC2p1qAmxwU0TZOwKJvLdPV5Wqjc4OFA43xxtFR7D4Wd1GKCnaKhek4COQ
12N2ETQwr3KLxGXmeNj6/9ndXwHD51Rqi4zHf1lzIEiLhcjumZH7AV+enVVtG2GtA+edmDXrgWQ8
BuZIrxJCn9bu5H3qiV+vUFTAAzoRojGpGzphIhjiLOd8/f1YrYpIOlePjr/nhPXWEe7r0LcD3rpI
Ao3RTwU6ZFtuGOBJFt3TyLrNop71MgJzuhpMclKBDJGi51hwtrbkwpZOaz0zSjl0DhP7icLV9jSZ
FjynI9kwE8MJ/2xvgHNBq/sR2elvRvwaF9ydco8RWXXCjrG8/luSBQy415aBzhvpcs+z5PD7csZY
jQSdORsDSGZPREclFJ+79ZhVwZz15cd2/WIqwh8vs1/yO/EYiFIdhKC6IZR2w3SyRAQQzYndLqjc
WnaIfQ3rciwvjntrjmrU2cjTSLFYkwpsLV8BgGjZbKGfT9/LdemoblwHJNTgt7Hg8WO/rUkmgf73
PEP3VIJUwdOx0BZ+Tcrp++SSeoZSCP5wIMUQHIGcmeCrZIh7NC69hU9NsSY2Etd6XxlG+xTJmjSg
HW2TZ5t89aLbCTuZMdJ1Wr0i1wIcVsWZtOmgO8G+i9+kHnq2ZUIxKNok3/eKtAQLl8NZKYzBWi4n
B8w7aGylKsSSO9/UpYLBsgvj2GqmHbj53SyVTuDb3Wnv+BMUVeY8GaHx4GUa5vGl52HdqOll30Lw
N+wUBB8Gm6VM3tSi9FVL0FphVYRPfZYQkU58ohnuHgvOpt4RM1FWRIYQhZCn3J5laZYITMvbTZKy
42nWMYomG5ud4VSopuqLlb5/2Otm0bHOzEO8McuBsNgQMTwAmPsMyOAPNzNDh6fR9mx2F2vdsFTP
DZQKPMZl2W7RU7p8z7P30mqL2VdeCr5CwBongapgPImWKLE9oQNqUrrlj5qgAEGegcGvWtuJY3gC
10P6hYWmiEUPk2VpH+s2FeeuVqX6elaRBH9IwaM6a+wVrbKVhRvxvBm1r/5E0E502Y5GfcXpmH7I
XWf3DzQ7cGUBs49MrHABKNz8iSdx3hESK0roe4EcOAIFAHm50Zs6Pe+fcfLmCSm4ilVzfwo9ZAk3
ZvQkk+CVM75w7KioEGMLKbxkRpNUwCCb4RyRwvzJS0ldeSWqvIzLX14lYhqigBM8CIYJo+UA8HoN
MDOYvUpLIIL30U6ElP6hxEkwp6k4rJGjrJcuz/n/mF7itgmA+KVwDCCIDLX6Qd11Rgdfovg6AQup
swmySn87nwWJTcaaxx/dWvYjwvHHZ70rxBxntjnWYsn8t/oi5UkZG9LEGYE1kv6uowopUR9UdwmH
sFu6pBZ25jNclekyE6fnpKRxlCuhObR7qcPJMJneblxW4HShUT+iBV/NtVIF3Af1Fi7nOZk91APz
7kk5kdRkJBab4wu9C2e1bAWjFWI0b+dndSH5EGQFNUVkFrJ9tiCwaTMrGZFhokaykVJ7kmOX+tQF
t5k3TkAHD/rO6rM3rCzMrmcUL9vtVz1tyrZrVT7YElixcJct9rTtmChiJkvVni7Ncu/0bO7wHsMT
deM25fk3JmnilLOJiSvZeNyrppu0CNPIo1l6gBATP68umX6k/j7d47R+iY9IRICmKYH23+DjoHZV
hgePzLR34hH5CpXs+erLPjb9o0TgkK8NvvO7PkCo2Ft1XUxlIdgk2HH9s+bmLnXi73lHSR6NkTMp
c18VLr6kqhXpHW0C7MqH3nm3KQ5dfbaUV+l+N4clJwaKgNOVAdLvQ8vbJWR6g0iwHnKoNItTipSj
bjCk1drRZ+DLZtfs/PtyrrS5pZH1iEaT77dVgh6D8C4aDUsBRow7HRyeGudEgy659JcQYGb5E6Os
BURRM6BtSAwgRXNHAmRXYmEjxUZ26ozeAMp/vufyvCCcPBYItk8HhQD0ZB3AWv0obdZaOECswByD
8am6zD367sElEUsr6JTpyUJ+cU7lKIkwTZNGzrVjusDHue1c1qDo+Qw2CGRFlPPe3z+FCeicb7Ry
r16froo+Gd6DAxY5r3aXLWnYqQE9p2yYbPEq44K+IK+9AqOd98Rgfj5OAhb00i/84p1XVyPVhZgP
Z2J/zUk1IkkuE8lFOmZrIvYbIpy0L3ZSYkhRhXsNzce7NMnrYlah0FxVa5vflEgWXseSyjoCQIBu
owvJ6oFJkJkIEt3YACrwMmTPbxP3rcAImduj5BktDhtQ76w+1oOCQeO4Ltn0byCNWYGZUF/UpisP
8TtKuwa3/3dwPKjzyx2NZ+EP3eAwJvH8/CZ/7rKgb671RXzimTWhozc6mVPuuBnaEUO0D/3U6sh/
YPvI1m2+Jka4zXlyek+J9FyZ3MQvZLFzyMG1tXwgUCDB/xPeVp6etyjoFQglLgN0uL7M+o9FCbzc
pmTt4zx9XnOrgPOCsziebBD+7BuwyxhHGexBE0LP+YsT4N3YQqdVXT068/nLVKCJatCnWIUfZX40
y6yRwItpvUFENJZY1nqHL5flwYnBTioks3eoOtuNCQql+/OmQczJuxVjVgGCAPnAW27xz1hBqW9K
0fv263rOhUk5WmyeWFb09A1kwRrT5+lK72e/xNPF3ucL4eh+GtgFSrL6c7rYBeJQj8V6oiYVlUi0
JeazecUSA/4ArE4s6/ObrReTw7/U/rWx6Fmn5utKCN20e8HuQOn41IhSCoIlLKkM7z7NAOJnxR3+
HJE2NTUPYk0UgHVrhTBduKcUDowvC7s8NNoMLuALklWYKV/eYuFXvbFieZubimAJRQLxB7DN0Utg
px8vXy/1+eJcY62QxL4FI94tVZerd/KzpePtZyxufe6UNultjmUGyJZQyZS5y5sAWwWFWKHgIxHR
pEyfrAMN/qNIIIraNEf1O4YlTwndPEXUUyOxhxgf3Djf/kthdzZDm5pYeIUQcdkn1sb7knb8ZsYG
OHpVkXuVtecU0LFkiB5crzmwpgoUXSv2F3BdLqbVU6JZhHqcQhefX9wfkB/Fq8S/g4u4VicMvxAR
KroBW4dJVXBrjMZotGCStUreavgYw/IgH94VQ8ru8cOI2YYUN/DhRXuVuP2iHPH5Dnj04ldW//87
tM2l/zKiu/d+cHeV3jdSl0MBADLJVI0eo+hUqGhKvy6v7TURD77b3qqw7L+a3hICgExNSCBF5FY2
hJOQmvOvsEK0hTdRcOdiyYvEQZaIbEIzzKQkNR7G8GAjGd0GXi5wXeNrz4hggk365b1yTJ3ABS7E
TpT7jHyLAB0eArx6ZR27oi1dohj9Y7GQVjOhQyE6zbsoKn87Y4wGhVpI5O7jSj2ybzi2HSUMTw3B
OkXGuOliva1L+wwqgNEyTMX2ypD5e8CxUEx10QHuuZAMNH5QxTYFmb2QyjLRFOmv+ZpkMDnsY/ih
hafVa8qMq8SAbTlkQQp8GOhTofuiv3ul+CA4zM1XZnsqDmowzTUZUVsxrdHpIqi6+wZkR+nPsHkl
GnZn94YnOOtNQvCdGE7DR0CmzWNvzREvQX4Aj/9cyYKWPhb97YZ9zhnF4r/OHdAoes06bdgX1mHF
hB65WVTiC6f69Hz4knicJjYvHxF3rcM68kxhcuAIjVF4WwxFKWRl/80tDEgEUxzoiUW3B/MXs47M
YqPNXRrMF2vFAvrfsVptKC5D/eCW1XR9WfE+r0B3V/MBrLtywE9CMB61UWa1dNsfZ7rRlPuKHHYI
4Mv4/V5N0B9ttUd1lQw29cgS1RIyfVPmuhyxUkM+WqXGmjL97R9xfz9Vdz1XuY2rKljzJtSu5piB
4Z50KrRNIDPdPG14R8AhIMVs0WPezpKcgsPnARdDmQtkjgL4sBKhPwgZiL8b5YYpmk0CsOYQWRP7
JTfMUVkNSNNHqtb/cJI+vWwT1I0eVEg+FZR0jhh3lwjESEHfTvtsKmrhvuJ+SkdTWmpuzFPpcyyV
TzdlwS8WBGxTP8SweROxwMwk9TMCxqxzHOHiovX74J8oFV2cE7MEtF4vddHCECf0qnURwycFp0Ru
VU4PPwJNvMzLzHpTGToYpNaZG+rgtqYMl38V4x0Kcaookb9vIHV8sIJJxkRypqBvDzyWDg0zl/1K
NZrLBzR7PC4mWByTFqiHT2sYQN5IBS0JR2a5NABk349kv0GNiXSCRz8hb76RVyOQ98YCns62mJK2
zhMik6rIulvcH00/1LDvb8gYQ6puaU0Y3PebgxQ2Jgn6SfwKHgNqxvuXEu403BLf6K35IRN3mm/R
J9aPgdgD2ZVLtpzxUa79jR4pSJxgjVYQO1Id0aLAef0pQQPr94rsdJSiCk9J+MJwg+XgVYD9mCNx
QdopCA3VccrsGeWawg/5iWWBZNnHOwSiYsWzsjJCtTdwFyPuNFfJYxhl3l+MSdTdUrjLnUTvY0q7
kxNTUsps8+YX4wDTjHeot+/m94kiHbWpQH3kZ1q869flivz0dosz9bbNA4oqbq+tMKsZeSvkl9pB
zTTceOZcFxR8XnaqQtqoeCQRFquD3OG5tC71hmTR6PbnO4auNrLR+vDJO9ApDVJquyVCkvYOxLZE
saNqpqct7nnahIwOaGSsI6xNm8vuxbi+knVSBAMwTu3GktnH2fmmXQRJMz0soJSVdiAWDkDA6VH2
V8BrM2daCNOQsKiuG8FKS4b83NxdAAJRADFvsXRV05eQ4F0WGa7+RDze9ynz/LRtzkZa8w2F7gdX
ZSAFoPSOVBymR8T/TDrqAlqnnklC4EHRzX9sa7cJt6yb6PQlYA2KNfKJtDsZhRSM1hOmQhkkJ3qo
3ExEL1VRr9Aze74hosgZ/7HQAsOB7caUnMBD4Ph6T+AekgrBiHCw6T03tAx603lCugoephYJmdWt
7bwbyYAmKQiwKkjF7e73jiXwrEdDrav9HrRpxMzJBoHGMkhIhVVAnmkLFxoWqRvTzaKL+vjne4j3
XZprVvzuQ6LBUmfxtoMdl2tAvpAEdl2I5590Uzxex92adCuda5LsncqyHZCz1Sr7JZrtEAkcyF5O
sq/edZXwYpLw5yuERILBeQirLSZVAqHrLyN5h6vnzPzgmNQsLoJ5garQ/wAfzLdA/J5Jx+zSOoYA
sjYq29Yl9Vr2dVif5msAVQ6zRes0iKGe/N4Tb+yRAydQien28qx2i1xwnh64dpGCjLDVLyGL2QR7
0e1IDuj6UMg9wJhmWIW9k1+tutWW3kNiuk2Yql8Bw9DudW8ZKQWbODwBP/12mRGkxeEe0/QkduJT
fuvlMO36VUF2fBr+MTUvu4hlKkuGcTWP6VVPWNeOUGHqBWO99c5uXkv5+hWXs8fwKrtQapT+A7+v
vyDwl5yldZSICgs9UuFCsf3yBxaFIV3oZNU9ps1pfDLs4dXQTnbzgXV/hoYFMwSdZUHqqyn/lBN/
JB/GyfS73REKmzeMLjSXvuqmqUac4GsutOp6dkTrc1F4xxcbBCkXhr9div56o1bpBPscBHVJKnUt
oxSmCR060MuJvStnunkUm1Ffv2zeeOdO1UMBKBUNa+WwWKVloKV2g6hgSHUPpGfgOyLPUOIEmZ8P
Q50CQYr6Vqq+pG4SetAcCXsQP7dg/dh9VyYY3Iu2qmj9N4xX15HHHt7ehoP8+SbPTnIXbZTKu01E
NXpWwzAWoyEBlS4IZFtZ/p6h4Y/Nf1SbMMfQqhND/0PUDbwzV8LonFweiuDNjJYOlx9OTsSNGIN/
W4vRDUZURf05x/B5HOep0UVFzdh8AITk5U+Y20Ba703uURB58GnD1dEnO7lZ+n+p8fCvPRUT70F8
UmURPY9/rRcYIYgJyEBogT89M42ISD21ztPVVVlogkPxRyl9a95u/ygzBS2qbEwJL0DMzLZKQOgP
RcR5Y7TqX1Ryf8OQuTlt/VdrfgXMRWg2Ios6G9aM4uFFF0QRXXELvj2w40KPc+OVg48bk1juOihB
DANSWsCDskD5KaJS2RSVUzM0ubxfpWGlWOCiWc51MtyJoxSwlGrcMx4FIh3rJ2RbnoamQLjZ42bj
hOKf0suWsIjjC9wET6adkUrnv1Oqa4jZz7nGXJLXDtjeKS1owFEiZQKgizGFU3jYrHC7/HgJ1VD3
FV0Rj5wh5C8qL8bPe3p1gffOZc2N3070J5Nw6qrITUlU4YP26zagiyoqvqax6lATX9zkin8GjNVg
PPCOHAQb4oYf/yA0Ebdo7o4Dy4Zbh1+/tX0L3optaVeO3fgtVpHiEpf0XxdwFLOYjCp/jEyTmkY5
l7On5whYKpNIuBOh6SCnCM9g0OQra8Ghag9fc2rtV6UDXHjhv+8Tjzmlp420bhAz5hHVt0kO/tam
S8sSEvJQ9vNu+cEYsfWZPLj3+wJShNf68C8LEdY20i63ALl8OW0N+8QLvXPPpXFnCWkNNkPLS/Gw
nzOlPTAVtwrazG1keAslMkDRby6FcyNy5/Sx0kAMzeqSnL8zffX9BfjEeX1W5p7R04naqDTlkWLJ
cekjezKoYtDAaia3gQYmqgNE9Ms9a0ppa9Ds3yFw9+7+jgpQPX37cySAOklDTCGJaHw7hFF/D1dh
oR376jXyVMdafA5N86BjPfMcpf4kLduL9ysJhvm0zM5HU7WY6vGq5teCyXHGUl49Od8hzD0i+mMC
fCVa/8eP3kfm8xzrJIvjI5oKdspwB29ycx3pJ9NyHhjQWFSmz1myOq5bWyPThoRUjCg98sQG3Sr5
W6lowCaB/mJX4NVUYCr4Mq22jgVpb4WUj5l8p3XZ9Nlkn/Ev+qZ1GAcqpeBp/CgYm6mY9y3VqGxI
vI9JcuKaUl7+gAwpCltQHbNsxBr9kz0oDJo0Urfa9XqHe5dQ5zsJKMHmFc907XjPoxpv05qTLKJo
u00kx0Re+Moq0x4N1BcO7tm2NhHLb0dCRuo5Axu/scviw+i//cHBBfCFLJGgsrPwJVrritTVtWc8
W0ocQdhw1JaiNx3+SupO09msn0f0JlIUBI8WfbSXlQsvDcNmubdzJJl19qpkoBbx2Gg9ZzV4vmUm
eLBg6Ukf+nesXFZdEbGmwpJBLQFQxarwf92I/pZwDZyE4HH8oqopDwiYa5bbfTBRsZFq7sphByWl
jRvyi/2XbSdvfyynHq2Y3DR50Asn8QZ8mb5LQaNKqLekDhtoMqxnRUBtAiWZo3KhuAxdG4+MiUeg
Umh3jeYd0yoT6ffhBiDgzwTtfNS67K17NtXeb9awclHweAzjlKzSdOGT17238W6cAMYqLPMy1ut/
5zwujIf8icI3GE0zU9LZkd5J+1Jv+1pTegoBJ9d2PJmHe6Zt5AU4IjKW1U7MHiGsqwvZ4XBXNvVr
R45XjMU9e04K+T8wCKSVph/4oe/Qmf9LBUfuua7XF0/GKFGhVa76FALXcLf4mTfp06mJMM1x4eYq
j7h2IVXDZOxmFTTTG9nzVMSyYMnJ5Kbij9M5FE9ZpiFNweXp/9KcRmNNH3aWLAucKUF/f1MwrhH2
KmMjaOfkrqStS/8z4wygF291r1exIXCK/p9D6azClNNfcj5HIlMRhEGFfMgIsbZxCSok2u1CekLj
G67eY6jl6qX5jxpzUqS2Qv/0YkR+HSQwfr+8TwsNhGeVtZzqPahT24BquTSQ5Ti95Wp9dniFwYRk
8xVam16w9ecVigDK7yunTAwMpq/NHx/UTbmwW0QzO772+6jR144NxBPaYW8WWGeLMTPeMlmvz/Ml
y6ws1mnxPShOXA/Q1JMF2UHqnlO4aFje1G18AKII8qPJMnJ6agyp/trx4gyh/Q6hqv9Q+S1Cojvn
ob4/tKRmpFv+pKdA9vGzcXvjkytTWfjPB1X9XsfueHTP7Ugu1pucqkODPEvkW+i/emB0dSSOJku3
tarApRH6LG/AaV845fAXcg42v9FawKTNK4igGg45SK694vC1MbrEu+n5QpA91EJUnMjQwoAKk7KO
kFpIFT7+PKdU6b/qaWvW0vD6UKd0skWhxpFlEAgRcfeehbeh277R5+yf1LMNw7tjuJTQzJkO5+pl
8jtblGAt3JMM1mvWDR2rgBKh9304p+hmWCoJH5hyiEQ2V/Lbj53FFrjIFEpGUNq7TuyoOO30IMiT
265rUFwfF8psojQToLACEopLssv7S4UV9sy8BorO1sPo8pEvgQkJPfbvYL8GReGzX1sJYrXeWlb1
6E3X/DaTCafXIpOaBqcWgCzxkCQyVRwvtkSCZY9jxIJOpjkb+ui9wct+zOCV8JghNoXmPkbOYaJU
8M2XunJW6kh9yiLDHkEoIxsRrZ1KQYLu71bTbmlIV+OWRgl+T0qis1mO3a24qMEQytAQMQ55NitE
7l8MIAuUooGIq+Th8nsEj/DUkD8p+LooXsdYaIwK5dsn3cqCxVyjFLG+04xuTIP5z8PrdMrxr9YQ
C2I4qBjWgdBWVBQz9W4NIIOwLhPcRB6kfedb3f29d7a2zitqYi8j0XA+T1vFUJmuX91u6ekPCB5w
0Ej4MRkq+hkPbVtNDPL0/agLSbe8cPxL3WL4j109GWYyIfR4FDGLiRN+F91XXXs40Fy+ST5hOg2S
q8Jd6qPmiO0gvPK9l9XXWrxy46gEY8+1wR6YszV4onETZ2V659bHh3sufpDG61IAU+jj06MAbnqL
b1C7TU0DG5cOU9Gk31u6rUXY8j36gt0o+iQX4DFqPAzwYCg6YOeHdjGOQiUz4U71NgMz9bIdQj3o
SBXuCMyZOMkFyRGU7Y/fkLKgmuLRIJs5BtprF4F4OqExybkKdSiz69hKGZywIRfWTgBztGFzZVhN
9a284ekJVrlSyFRDFvQA6XqfSg7LIwEWX9Xy/fWY3FPAyTQ2tnQwi5iW0K1zLw1juc+InDjjuuQy
dvdotZfN2hi7bF+UQqjsZ1vNzaWcyE4cVM9esm7VYkTx/xoNdYLq8GqS+PnZnFmm3JrC1mnsTf0s
wwCznYEcOw7BBhzOe59NdCujlXtTbEtHdDsF3ePH5/ehKvvw1LBz+CJcDwRHbZHdA29VtgDi+QH7
HJeR0fhajG3g/9AY7TTPykhwIlMlCJhHHioZZFbOKi6f39zou7hUusXu4N6e2BMPRrFnLNMcghli
4CpwZXfSLX/qlii8Za2HeetgZ00lpZ2yfw+NiOd5KmTCpKlhRWFQLWyxAFhZpMbtn9g2AZaXrluc
graprvL6IxIENOSSD9g5UwVgBNtyv3XOJX8ZQe2w8zokJExJk/fbtcemA7sBrSoN0wMa4tq5z91I
37NWeJFg+Vu/ojSBE0xmBUbcQNNrC0fz9KlVVPHcSuKBtGK7IZthPCX/Tsv4aIj7U5dvAetKHHg0
AYF3T2foc7akmPipeSA5VHIK/+Rtm52KNUb6BXmEFBKDAqOFFCdP1lMY6Mz67JgHFgAYqtlNGCxj
J5e7Ijfw5CA5nlt1cQ0Tud8vuU0ArYGvmlew1zws6cZtQqBIeOzuZOKYaTxC4x+lclQV3q6Ba0/t
cC8OhZtSkbY7cP2M8dHsC3t2sK7rXYUjBgtU/lixMYUfD/DIK+kzta2/6tPCoJyWPhtrqqy091pW
flswSNqr6yBU0BN3BPXSsjiJR7xsng76C5rlUAWHXC1LYNlDjCohWmgdqSUOa6v1giPkxOOoh9hr
PbLxDazQ2PnGS0hZF5LDHfj+t9kjfQXQoUm/97FETEJGbvT8uENdqizKPyCxn9o/p9/jZDj70sT/
dBnTurIAY43rz7AFKBgdvpFhSk+w3UcHMLVn4trioeyW9ENYURdo99SWFdlQjyO7tl7kAI0ni4fN
Y0TB+6gRIWH44alJFUZLgoEc7LXkRNJybfTCTB11TprxgTMPueNZzBLqoMGHy3TmNnHd5pQV5rsa
Sb4NdNsrfT6yWAcssAXesU+Th3q65KJ12BNtGfy51R8ec5q3eLnBYae9svI+53hs264SK5C2IT2q
NPBbEoz3VH5hf52dXHL4UuADnTFkJPXKtbxoQIKRARDdpZOTOcGPkvP0ElUfAZRzHridfan+9F9M
MHD7Y+Ex13tJbhpZlVzQ4LnAVey+4vQ7jyerrtFUB1btfNQuOQ8/sn3sqfj5SWd5qsyzqjnn4PWC
Luz0FyVEfaUZU8DeN0RAvwGomXcINiWMxGl0xpTrtkU2wJ/2XDGHUhLu9ZtX/T1UxMxAiF3DEeRV
60QARsGBcBMJo2Hzvdtrf3R8xDPaRDMzy9nRqOpMkuh3YAaIcFGYYJzpeFPSIEkQgD0T+BwlE745
L38AhNUk6BHWBajewFLX69GHQ/d0Tm1Oy+e6WeVbT0FticDRQvdhain/XyR95UxNp+PBbOmJwyA3
Zgrj++cCoR3eejAGBKw4x0FpxSE3S3cWHemv7GV1DEbY8vfQWTmtTsmG0ezkEWlrELfgr+GNDMVq
Nrt7ThEhwGpmBa60vbW+zdgKGjXXmnxj+oq2oY3VTo/a/rvMBDRhfy7DeNOq/xH3cy6HAKFE/Mbe
pYUSk7uKsz9yCTKWnk2I+Fq9N/CfuLIxj2ZtcMqsXhw1Ryiqi3Y9dMJnvVPa8ISN9eU6z+Up55Su
AuI3/ev4U7OV132xlQ9fc9PI/08iMht1PV03KFmSkXrlCloQDzJ1yXb4ZNjEI87DJDsJovUBgNNv
4kfMX0H0pKQ2tMC4U/e3a6TAIrWN1Ziui/TDz94jpDMU4lApqfPyi3UaD1KryzHiG0zMkcQpS8nE
zzt6Jh9GfRzGCx0dJkxHgnS+H1WGwyUUwY65gsjKes4BS7tI4z2qMmlQg7Adn6DIBTPRGw3zzpbo
X/9KiVqbieCA1VEm+JKZXCL/PTlCnxk/FNA9jJyoSIhQbjSWR+zOGCCGlpgzeS5KxSSj8EYWm2xy
H1BmbNAzWo+s/da+uOaBsziJ4gSpywlr/F0btHo7n0p8j54Vw0fHbIiin6TmuOdWzptDGeA/oNTm
5yUHj/o5ohGcIwWQIgcaCBhg6gw8BnXiWv6AmZbalEIGwBQe7nXNQHjfWTTTAchgtDarZifNs4Jy
OXcMEPLQvha1sqmD7dq70UfiFBhJ5OdNKMMzZpKNMfIQi2stGDx7Rspisx3TBP9hBBm44DK0x4u7
jN+hSZui+lhWSZDowxAEw9V1IHw8LQXoxpxV4n8//HPpUr0wSp+EBM5TN1jgdIThmosaegXmKayF
MAV7udPlC3aabqreT0BAEbBo8a7CJLWSr0mXNcZZk3IV4LeGspe5UG53u34m4GLBTYIDyVpDjWvB
vJOiuec2IW4la2R+vcFO4oWLXHMG6yU+knmZyw0iSWDhvly2t7yXR0bjJ8kYKrC5i8a0MnRUN77e
y1sTmnQ8JnDI8ItMJYFirSaHL7YcgSYsfHJqfDgFT+qqyRtFejWfoBdCrr04C5mHZDSEOeidMDhd
xh9wzqLT2vxwdP4foNUBBGaHTnq9qQ3MB7ALbMkdLAbfo4jus3zt8lAJo6WOCjnqixqgE4wVuLGJ
Fq7awCEiTlfDLHd0J0SO0Mlx/tuYlmIsOCERonsLvUYAfZdpHT6F16uUikiGLUnEbAjxiCbmHsBt
XDFdYt5LTQ5jmA/gH7OGNgZbH5N8Iw86SDNIqGI+XQzJGxKu13S6Nwx77HlE/5Rr/sBD2uOYt+7y
tlGvoa0vSS+f3Z0INCrXDpLtsyXwomrwYFm3QZ841tWkp7Em17S9ca7SNJNIb+NOQjtTvplUETdx
LpppShcR0OK0dC67MH3hcdKpCZbCboDmp1w2kvje04uEgX2h0Xs8gpLQsu6+DbttymhksNjJN5+N
8X/zPuAgnbjF2RcOddMJSIgAaXl/RGNaD7Vya0sZt7LsDb4QIscuQAefUNjuwCvu7kX9mvb27YmF
JvIC6UkTgqHMQCcdd3w9A4q4hw8MLb64+O0Oq5TVVs1bFNg5UaCnpbeMgrcp9fUVWUVncned0j5T
w0gGOgrIf6XOMdIoB+UmyYydzdLX1B4WURdcweoKJQa96CpU15o/47Zv2Om+14/D45WYWrR2Pp18
mYf6kfmg+IdL5XLw1M1k7/7IX7KjaMp3OZxedtGkoqK8C855o1wpzxnx6BqrXoTc13+qqTNOelhy
PNwkjT3z96Oo3najjFWWHJsLlk5A4v8MpwH0JUDBofRifMdDwKXt4ZMpPxyaHC1uobOWTjfnIFLW
dHULihD07DUjyMSv+yEZuddsFSccPIvhlv6RId9tS1GJDc8cxnvwOlSW8zzjqIUJDOiGR15oM9tY
L8wW7TQGNznjEwOfnt2fbdQ3uDMFbv2/0b6WHt3xYNg/KCjj+ORWX6jQTdjgd8lg/42gmptGFeJ4
ygfXt82aQmuZsi0NHy85HXuMpwDmqt3P6SaSTEMZeDNuYBi0eDy3ZV4sKdEfFUOHZsKIoqqH+Bpr
VPQKEwH/+t42WKGJ/ibSKvLq8IOyU0EOl6OSdEz+SvMuDlMBSzMoqfJvlPJCv6HLsGipDMouqNPV
1NwU8ITuffj+J4LSyNfw3mT+HqmXGBXBi1EMKmny7P/JRbOM7hJC3rpRyosFizLYCz652if+8LVV
1bELzCAXoO5kEPCuowQOQF6RzexLkzuwfMCn64ze/5u33LSA/w/0OIDwfAJB9qvXEeImGbEjppcs
oUJqseHsrWIXqNhyH1e8gTySMMpDP23V0/1sreKuhnDRlxalKvZTqXe+wgyLH4bvyzjxLZjHuJFs
QDBzcjGKk25/zS6f4UN7WA0suWrMBKyI3beZUMSQqWCLj98OIO3yj8jcB5pi3Ucki8x9yPXjDIXz
Ds6K3+5izaNwKHEbRWxRcD9lvu9aNmkJypyj2ucnML32Wf4VdvbvOu819Rh3g+ODR/hzErO2Fs8W
qm0rxApnYGzxwYMsrRHdxXGUIoNJAF4ukT0E5CiMcqT+v2CQoTXb6D9vSKj+Cb+59m/SssrMGJBn
ePsAqTHVBbpyspreUZ6HCT3JEz5HJCsSJGNwzraS7H6SORt6ifOyE9px3w8Dd+1jBExmq3nPRv8K
Vi+kpJk13T/IA6S7eZZtwgCoOb/WSuAkUR998gDMHzRGyCAqC6jGEDtuU4EO9upy0MFH0Evijo7p
D9d5wPb190ZD83CEMFqIYJvSFHT+5poU+zFylEL4diwqusYRxCrwUgExzeepxwuEET0uho0CjyEl
t83kI/PfRQgqmfFFcQ/hUZPgHtCdPJKnC/fA3MTfHc9ODy+OfPsNhKHFf3iNIUXbdhEpOGFKbK1z
5GvLZIVSH5Op0q9msikkS95+Vn3olNXrcMYL+pCVgklsfSnZJkJEjhF3zQYTwthBeiiB0rSb3TSH
xO1uDlHdE+qb/IvI7VPQjomAilCxssCzDd8q/U9B3zE/ktuQZfnB0J5P6nRTKa4du7l2yF3bysGR
QfHjqNdeHwNPUA8xcu6yrSLVHW7i6t1bZm+iq9m7oWYF+yqmS3gCr2qzLFcGwbvCSc167TbGdwk2
YZoae8qSsLqj45+KYs3MkO4XSroEfy+Y2KABPApGawd3D7Q61Nhqp7L52GqK8D1lrcckVC7drgRE
Ymm1aPfW93mvb0FOGyXxWOx6Rs2qiFe39XOZZjq6xc/Ao2drGHgp/3GTWgraUYza6wPoE6l5vGuH
ujUmgD42/V2ob6c2SoF0I572dNH38q9XtGcGor6so5oGBsE95dfRry2y42hPx+iS4S49jAyRGWOB
Qs1qkZsta8dmgvpfhJS7+WQGCDBzG0Bjbjaa9S1/X7I+ifq7Te5mBPrbraFj71SsOtPAN8UT9nwG
/sxGALkdMxuJTLBHvIph23e9hKrwsk0q9D4fU0KNTnb7Ckpcjfy5CGsuNt1xLogqI6GRwo0o0+oX
dgYPMmITwPhuAAVEv0E/9aXsOWzXxRO5IKhYucczYsHr/YHE+IP8id9LxQ6a3zoGpaPpTqCHO9JW
ivmMMBrtN66h6xUQlSnCxtAJtnfdGt6kJynmN2VH+PqLJPDr2H6bwOyfZKJ9PvdtWVqDZQVZ+PhQ
cnGPfpn8raLjnM0xmze2u+Xb1nnFublY2HdZpiNTxuhW0hkEwBDTSElTNnAvu5gl2lE8UdL1WhN7
3EcoeKnXkmn3aIpe5NEIKQk0bMlZZcUs5ZcHP2RK4SwHvxv3jiYkHmsTM7FPtxXHIJJZrN2pmbhL
mgLGi2PGAmpB0lqQD7mRHXMcGzB5yl2opv0l/vy7CAGefRBAxiwvchC8NChKecERpGmv7zuQ6LbC
96VhlzGt7S3OPkk1LX24KDdGplIPesEzv53uSr/oWBOeZXHfrOB49m/hFulWHtXtZi4u1SSqgmoe
nNnn3JUVNep/Zmc5K9S6uFmHWgiwkAlQD7/LUHBNBPXk3wD/d6srg4uOIpnMRrL/bAteQIRtiJ/y
cS6jOT4irDndlp4xiBLUvsiuHUasDKbH4ls2aPaOAaUHnP9WrEWerB4/1IDyqXI0sWgDCU+Zd5Tw
JXXtyYhdsxPKZ0jXUZZeY3e73q8Vj6HAMBdH+tlrNvaXnj4h7shu4yuOuDdW7UAZ7bpXMHU/rjiH
lEx6Wdg4sGSzHiBU7Ax7PJBk6Sg/H8U1gcm2lmhZrWZkiVPMornv9R+wp0tjeg0vPYDJ7wBYSwwz
BDG/hvrATEXsXIL6CG0PgBEzrxVQfYiHbQxm+BPcRpInnA9s7AWaUbW8BUtniHSprMlSBXQuMfPP
NrmlY80FmdryCW6+ZS5Pvov8I+A6uUXOt3dFWFeucBI1DJF2xBrrr+hlGm2GN9rTsdt2uZHHTKLx
0pUw8gWICHcz517JuQbZkzeY2BpbCxB2N8txVjcMLaEx/UORD+Vv+j2fuShViwCCCXwvBJhCtbnR
gyHsoGG961NkQTMYHU7+ceTD41LJEUgHKoHLwncZLQSPUJSM5Zcq5M5unvK49Imxk5IkT5UgWL+p
13FyTg919TbySjh7bwY5xQoJegSW0IzehXLcDrud3gCxkIqxru8iC/ENMxL84IP6rbkvXGgoFlFu
ZZCcaDftHtKWr3ZuffPI1QPo0SDMOPoti9cyiy8l0/T58v5lbwrqvyO6Jr/6y/SSsNp/3e+YNdrO
iB6pPwj5bNvPEFn9rEaYcKdOQAlOEgoLjZ9ZbitlfWn0ClZfGFICGhbcTYDBGCW/GtCJSMHdd/qU
NCjo23KpDt+cyF63VK4weAqmPAqcYvhEHcE4W0gXGKQSmi9gtsO30HIqK8mT6clXxcmGzFn2mudz
IcpGbA9HzlL/SVDt9CAl6mABvcn+52IyRxpTl+60+zQ8Vf6golCiMs4mYSQvFCbsFjHidXpHKKod
XywjO51DM3OvM0PqPR/0QwugW+YKClKs7I6DJIYHpnsKe5y0RaV2/nTnO7mgjiGWpmatp0y9OjRz
66nNa9IvQE4CZvnEyHDPpIZICYW9F688eBsCiPzS4Z/9AbVC4etM+XjjFX65XBaHMnLZuzIdEnH8
UU+evIQqzbqCKuvrnDJyy0EhiCQSV2YAHXO22ez/Fkx4yP1YOXOI/4ynwqAYVBAAXOtUbIS2YvMF
GgCLxxlPryp+fjwZfCK8fRuEFha+clZIfcDgbIQhTPxZNeaVLmy1KqvBonIu828CopxsbeUNNmcB
Lm0eTGrQ8L7P0h9dgdezoQ14I1e2KJjAwuNHoE5uxzbbMqY6GM8gfqE3hGrVGo4ptPn9GyM9/u4N
OrndRYlui/qNaTPWtnKxNP7v4/ylXBDpqMrr/6IUqWiz69AQG/qKqaiFI5DrIiBVJnEwjtake8n7
jAjv/+nUdGTJUwbxH+aM0jH4KlesS5fDHYe22l2LSBsC3l2JopcoSesrMvEHmhaKNKGwUBhtMRx7
bQ2fTNhefBfG0iJWNYxJKCqIGnBCiFuZBNNOCHlxA34QD8Q+LUJsFFa2s021CbWijBdtd7aLU9gE
8j8CT6lWQZ2Z3cl2/TPd2k+klD+Uuv4fe/HgA7RID6UZUOY9CSqZmdesRU3m5o1RfGPd29Y5Gl0Q
7ZttXZjGX9BLp9BjzCvl04YEUzz3woJJMn8ERVK5lu28Hlk0tMtUwBfKvYnMfyKZpMkydeiOeFEn
URIpoA9eBLdfGR5EPl/2CTqZVge30sxetQvEeOzUMH5o1Ow4aOzCxtjZOS3TFkp8s8fccrVFwtkc
gFUgLarrIBCi6pImNCP5DTKCbv0DAaXqwbhQxBlnBDtrBH8VUgZLphHn5kCGxpI/UhoUoNIJDUMg
fuBrXwsFPwKKPDaa9RkGcdURTBs3VTHlSZubrFlnBRoHp5FlhE5MrHQORt6h1b+Mfv8PSqulp/UT
RzM16OQ8Y3/fgzZr8vaKcD3Xr9+4fm4JuUprlRgwmvFYMw0u4WPfdVuFFSH4Zsi/pSGCiX+BHVYR
ohJQE7T+SDopXCSKFM2fvoUZJFsOyKZCuYFa0k8aJvexLj2hQqBmmfgsnQqHZfY+y+YfkyEXOUz4
9qptrYW9mMflkBtDRrfK+rmVJVyEKeMEVYucw8clw2Q+6nG3V3kTx85o6TRnjVDfgG4zSqfS7UYB
VGlABbnt9g9/cPMpFfEvME7e94qo7B2oS7hO1TX8kOm5wivUTUArvARLElwIbXBKcADCBYiuiRak
YZMRahe+YCzTYGrxJx1oAWyFPMGoCoYCo7iif4vlhiKDJbQ0n7x1B94+LVYJ4QB9RK178oELrAn8
45Sr6MVgsSVbscFwT8TQ8qFz5xoFZvyEy7FqrnN/2EUnWRc9+kHk5ofFORk+vO67Cp4Zd/3S3Egs
mxKige1X+74GFtyebeS8Xvx/GdAs/BNhqRKVwPwBzB7T49gLxQtT8uOe77JF0WSv5B8WXqD9muW6
R6Iq4NRBi3TaIFQ5q1Bimb48ltJ3hIxga52v4GrMubsGu+ct3uV0TmAqzqU7yWL0YAQJtbYSQL4o
HDYkCiZBavsj0gXhT5TTagWpyncF6GXrlQcNRaXaNnp6DoSWv+2WQ0osdZjw3mrySCOEMs1e3IC1
pqIYg8vM1zA0Ku2nBGljv0is+s2ge8TckQ9y6LmQenqASglqLTQn4DXJfQ+UJUAft+5Th6U4q4+t
6hz9LsJJrw1dChBxkAMZlcZ/1MymGT64CSETYx34yWUUt60SiCG6eolLX/j7vvZKG450ym8H1NuK
g5c97AkrRRUBzXWqtQHiv6jqzv2ksENOW87e+ibOQVbX3Kw/nB6DoOzE9yEEIGC7NDNqtr8xiepb
QyNHJB+SiwV0KRrBe5k252i9QzNKl83nrY4HzlfRJjG3hzQAwMXu7H5HKdxynwVRubvsicjp2Ism
KXw0jLiiipdkI+YPq7N8Gbl7SXb2pZjbAAtZhQTSDCfCZIvQah6K8WUhr7MIrPlxmwmedL6m8Bwo
3v+artm6aCCZSgXQGrFREbema6rSdTUBlu9vZCZ2pRj2in9ipZziQW4EyGIMr6VVr7ZQOrIy/irz
GZJRNeH9TKCHpJVR+zc6k9Yp5F0BV7qP42XSGomNm7hnTvLHRtI43w5nHIid9dI64asFGW9JWyzk
oScaPMgQYOm2ABBAUatMq8R0F4i2hdiXc7X3A+Odt1ypnAiui8WgqHNhHZ/HMOyGtzAhe2Pkt+Pn
gAWsuGpK+b24PsdeEjKPYlvOTBuaYLWw1n77jqix13EhNPmCJirWeA8Bj1KQnaAU2vXqBCvpDM4j
fl5erSAUHlo3/RsOsHlWdZJNWzN6irBnfYaj05hQwKtxyp542sKgTDiNTKo3x0m7T9n8958xGsMx
xaaYaWmpSPjbfj5r5CeVu9idk0acdRBk+bpalqS24U9tfOlq8RAhD4XqOjMHoVwBnbit+HoGgFu5
XAdNpeeYv50jQJ/1Jm+lKVX6xvz9eZXZjGf4qAhNzhrsWs5OA+kR0QoIuTdGj6tXpuoVz5suEYB8
WX6mcQAzoy2311NLsg8dqLQxxAJwgCME3n9DyqbyFJkPUQ/1OsWGurha0D5myCcyCoYAMbxpB2xo
6QRbXrq11yEk021aM38NigyF1+IHE831a/UBcU+jMlWI1ll2DyCz3/vrG8eEd3N9x9payxK2EQlc
YQyT2DYIKvcSnuGtSSLHG5MO2TiIosRwCiQD6QRjOGMXGd23C0hs4QoL1usTlhKZFeAd2IirIAr/
iL2XeZ0NNXb36GVxwrXzH5G6VilfLRy7Y08Ee/5Wh14yQ00okkZfqCEi8cVpySMRSMiWBAdJ8xHM
o71S3JxhCV+67XRxhuPOZx0s5+TWux2Bfccfr44ohwgrDtpl5N/Gwifbb2+N/1lQvKEp1o3ePXBx
xqlJtwWWvRq9C5hyfgrun0Y0dn7dZRYoIc+ZCjA3vmefyPA57FfH4jdO9VaZVqwjCluDBN56xfQG
XeBLILXWvAioh3zA7rjy56CLGqOS1hBFT9S1qoRYYgEDG0jISoCdjVvC7DmO82PG96rZoxk7LLQM
65J2mF5v20wG6hF9qzSmkgVw+paj1FjwE3rGaW+oxJKNz81MOGpkIRfmy4E4ASA/qBnERRVYftda
Aa2D8zkfXsbthXe+egJnk/UFziEK9MabS6BKwoVrDCXG7Vdzfx9bux4LR/mR/tfF4oaSERXyeox4
3ieHIbvNlmjA20LFheT33iz5CsTC9wZQqRyYnzCMpvVAHqwp/VxR9lcrb/91F+0ktAbW5hwjYiik
LJqlxAg6/xVzka3aBfD6Btj8wuKF8/rzNYQd2exkr3ocjq2AAOQ1Joy/Z4/2scoNh9SQduvGonrZ
WkgohV0ytva94I3lIs/27nGGORmMggi5UXLAVuM+IQs9Om1aPY+YfKp9OSKkWlwFdp9zJ7tAzbBg
nlbj8yypLNMCkt2dOurcmmPLqnLq2Rj+xDJdRB7AEpXB+QLE0OSVeC2T3czi9G17Z0Bha42MjQm0
z7qcjkKDKB0bGT2x4cFwwHRo98iDCuq6YNi4qk5KK1nP9UI52MY6BtLMHGfrGEWthoPW7/4GMg9E
6TEXEQg3xQY+bD6+I4wQf60/82qwc3OwRtsJ49zWA1Jd23baKvPPSyU39e/rAlU8HWCyR02V0C6K
DBhbdntQrayK9eXui01Etmzj/G2nKvLO+C9hQbJ1QYSz93lC94W4Y4IeCwQeXTl84eoDmubj0rLO
MeZmawX+9BhIcyA5m0DrcgtAvkixdHvyM9a2+7ADLjzSaxFK17V/AsJKRvDYAjorc3PHJmJw7HqF
6iC7+SlU5jpXEHfr03Wy0soyDZgpwpI955SuXQkMBWw4Dl9qUIag/sv9+zLzq4M9xxXDfzaNqrzp
cMBoR0zYiUq75mxucDIkqPE+Dnu8XB3kv34/VHrqcNP3CZ0FftwDREl/dbsTuC3sEn5fKj5KSXmB
rQzqobMelUV3VTp+kylE7okBtQlvw+n7bClGujnZfuAhAnLcImSkNu0NptjQXaNxQXpyfTBX9AVf
c6ysUsxswhs15lMystNbK4ZW9exdUGf6Iy1SWEdMGZ7mjxiQkGfpNHvJpyCorYpACRIoh+mNYtPu
Rp+UdtkSr1JYWwBY9knpAK3sRl6uCLIh+ZYtzzpXaEj2yttwhpMVjGQodvMoZF9pycpdzO7Nu6Eo
ceMQ9LbLbnTn11e5Xsgy65dVXx8li7hIsb4iiW9Uv5hAZFwRy0XZNCwdVNnPu5U3kLxsb2nx8oLU
x2D5lvPwe/+aChRRWtZgq2UWXx7oxp0ZGth3g+Ol/nWjytDbywI+GYwSHrXvNY4aUuBM15R5DlOc
gM1sM2EdDqHZo2S9uTcWVGOV1JGp5VaseLYXCZywHcrUFNF+TweQYAt7IwvSyk2Dp9Z5t8HSr/Wi
8IZqgbkEaEg1sD5aKjj1QbqSCj5YFzNY0Wiz4A5iRrNuUbMMLPGAdus/m7PU9u3aC7dwStP641Ik
qcpyQ75At65TzFOjj7RLYQUDv5WETHk+CfEyTS8wK+HhifRrmmwQN+GQiDdEiaqaalki7E5RJQxz
P1wpZDVrQWLjX9o+3kPBuQyMFsHRWf8y0SpldePNXVQ/d89ug4Ln6Qj/6rcX5c5lqu3rYEvWaqxp
cYM/aO6TkN+F4jUlhxyvPW7RDYU76jhHf26+k5YvrCGXggZ5hWpXckjTCmIRrrt+3zBCR4B85VfE
iWeWgh2016bUz6EYYY+nLdO/v53Whow3DaHjC0LwZ5td5dLqauWOt+XJFABEtaufzdfMkGR1Ps1A
SW4ZEfro/ahOsV34iwB3tRizuPiDYNFMcckrM3J63LFLPzg8llooCQOicD+Vczvbw6AHOpxPARRQ
9m/b+xku2mg446rMoGrXBADBKikymwgGSZqt0qezjQOpAKv9gVv94rN5DANPE2Hc1PB1zEcqFvBo
9bJVyn1MqoIPXeTfBYPsz18zP4mgRZ5iiWnzGWQ7v2k/58L+VSrstFz7jtxqJcv2VGVYxwfFButE
Q6Lrl9nuCBvrnCPPP8y2YZ35dQjz0+2kB9HsFzCibL8CT6Bg61MV3vXd5FWho7jI553MevvHy7ta
u09IwIsh8TmFFuVquKe3ZYUGMFkufM/3JVAtL0mui0iOmog+487PMGFLkkQitY30388AAyNURDYB
9nrvSsiuTYRutaVX/DTBYZuWA4B7QVn7uNozHz4lJFsiH40ab/NdCpYLcM/eZPi7hlKl7IWYGr6f
x4wYmZEjClVh5sTka4NVwIiaDowI2Je2r2ZoMNzMJjDs9YiZacnybZlIXugOgy3LOPxuCYtjFslu
0ZJML4DYAirqkOO7+k1Avq64wFNjVP6xJvzJU6X/+xjMVRssh+UYvgSMczT/UguuwCbMnRj5vsYO
Mua2dEbArs5HW0sBTC8H2qxpGpMR4kOvjz58Kns0pDjCo0GY9mCl+r3i8yN6GSYGSrPbc+SyxRoL
FoaU1rrVL+cs3+nTlsDUxceTgodRUptNIQHmtjdS2Vbx52u3Kn+TT31I0Hb4Rsdk+Ba0603gnGob
YFVDFLpe4sA9lSpStf5ksUmJrnTvMSJSNZuqgk69Oa5zusmeqaAVPasTQK0vzOV0aIYvqV3fcTag
siRRvOlPcFMyLtZvp1oiILINpMcCc+30zrJ6S1MmyI3Wx4120J/uZkEBcSYgEY6lkrrRXHisfhFZ
YH5Qsvjj27i91noKAUFtwPuCg46mJ9yzDqaN/66VUPhOOwNPwJyw/zunuQj1FWjlKfdsyNNeYnTo
aTwuq9Si/RE9Eb9TiQ5odbEcCkWnifMElBKVrsyS0yDyok6PKJGxs7ddO0G8/jin9krycgmMkwrK
wgsnoxerjoycnjPT9DoW+I1V+Ivgy5N89XbIl+qYusXGxwLtN7bY7NWEBA9E38Rhlu+ycS9/s4xU
9HWl7fxXCyn/Oc4/XBUqn2JMtWRfpPwZMC8RQp6UMBNevgZcxeSbOKfVh5cqT+JttIml5baE3IOm
VNvhzUGQL97nUCzLfHIhLuQAOrvaH68Pl5CH9RShL5yJ3iLLsZtiZ17VzMusrITNZwA/8lylZZ4n
nisFuELQbyBy83ZXWCAeY3hbPuh1hKYrEMQ+rbEqSRUC/J81bn0j0vsA5b9iDvj28X91uOc77PFK
C76UV4EU4jKlIGT/T19V+dnx8SLrqHYlon/6yCZdMUE5yWFEvZUAnpi3nFXrcmjUMYvlAX8MNzU9
t9jk24bft0/rFOoWIEq3Fk4deST+9A839qxDmH/Zj54mhqeZ9hBIY1ebBvhpP3U8BZazzerCx7LI
5X/1ukSw4FsDX9sRc8kvNI6vIeIv0WOFIHpjHGZdpqKFmOby0u+m2gSMtm/6ycyGQWUR3PYZEOXL
Dk30nKLmUw0kBCOv8+UdjO/p4Ag43pW9jWUeokWjx5M4ADju0tz89pBfXq6zJYTuO+C0CtP30TN/
qNspip3y9gRs5NNgqYP51edMiiPHxdHCMzPcD0dHPybu1WNVITIf1XVOJ81l0u4I/VuaBD+2lEvJ
aNlHPJYofm9U57RSNLo5cAsI1qmDH47BtFVwNJhTUdheHyCsjy/r5joULSnKD/VHNbF/t4K4LsQE
+WimZjCTkqIessR7gZO1B9P1qXprxp2Pkvj8CgzYGv4tfGAYSxcZrcDpPoQzu0oAVYrbcebEMs4S
NvFolA7CtgbkHVl66uVLkhA4Yc7n+uFkDkINVW1JeHDhFnM3hjHIAoX2EVbdfddNkdmBQ+Ri0FCo
4qb0TkKBdB5yemD46NxkjndMdTSqgA6k+LzScNMJsVLM2ZFrrb6RQHRtsoLSTc3Y18TRXgU7TvW7
qKNWLj4ebvZLugQwWe9qErIspX56QroJDrh5C1L4k0CmPYuWGjgBg7fLuXb8LQFe7rAMxoFDzo3k
jzy+pzIDQDmHbl43dG1OepODT1tzj9FyNB5RNZ8mKNmmvHIkVVYXhS0dkqFitnJO2K8rcx7EpJ3S
JOl5czTCG+O5TIf1/wCWFXcrZvOQWwKOQ56AnvwYKi2EaTF4I+3oAGoIZLBof0O8+HsQge4Qimry
5uHHjnzeUW7/83zUygVGd1BJjn/fcRG/kW8RbQPpF9X/w49HqQ/kSbBhU23JFrWPRMYrPB5UQ8B/
kcOLAdvL/99btUHtvnfbQGjahQoY2BxT2/+ewud6oGB+O/oggexLGD8oc9lbbQSbB7Xj1cLgSOmh
rqQSgXA0rZ1tqE7CxR2dO1X+Yc2eKR95Examls7I+aLTEFn50aaVa6JkEmB3Ty+44PvPWxl7T8qJ
DNvVTk/uxjh+J/XyXiGIzlLLNMykoR5+8uClIFz+Z3ZfY/eBA86pcGX/YAJ59aLaxDuPcvsncFu9
V2jtdioUY/nxnJYVW7i+0gzkfN5N855H5/qGWAn0/nkqm4jTzaJff0qpCi4u4GVuc4illkLavlOF
6LsLP4s6tgt2ejjlWrRTXTHlNMRJhH5CGTCYc1kOGd7Ze0DM8O6Q9Pl/J2znIIqlpp1TdoEHq3jp
AUqL2IcGCR+7zihzsxmaa7nSvv9MfvRwjWLOZGDxxXW9IZivrnDYIUnL+6aMeF82dYv4ByH/uO9M
DW3amBF7x2maZmQmyvimLlAn/gRjwuLEcXxyN6BOWNto7JsMICc4sqw1sr0ehBkuFUSfH3BxiNuu
iH0Q+/GqoVuk3sspHwbXjR3NP6kUc9Q0ukyzz6RXLZ5C6fmr1cmyaB7NJgQ/KjvHUukJPWdDogge
HUBJWmo2Pw8qbvtje2Y0dIbfemNz1e12KuE/D6yFB3ZUEfhwQoXXIt07JnNtlUcIR9X6mM6W9VBb
ib6i2CW78X5jVt1cZk/Z3yllfrdCKf5sYEfBnTJAMCUcAtxbs2RBgqr25RVyh8axbzNGpCEf5isy
IaIKTPnFOxzeuG/GGdcN4TmVK/9YogQZFU/QQ1a+gxuOA/x3AD8OwlEfSLkuS60+l8cA/TBmeftZ
dd7bZt17t49JO1vNDVQH+uu2VYFEx6mmkflO7v6X10LkvYFqxTyOl9ukbxGogy/KaCgBrACzrmJf
pbxm8oRZkMFQSsQVfOEtM3753rTrAAdMAk+Pwp1FRfRC8WalEDklJquDTL6BjtPEVvEZ2ftVGsMD
YKUi5f9IkBacsBJ3oApRI9sE4gxDWcgtE+z7hTtXBtB0iQDk4vnLgES6SqmbPS24N5PCsHZorzOt
48rUmHb3xQwUm4wa1AgjwygBczYecSUIGA2xfgwR5lHR2rRXZkpWBqgZZMJwEAsrFHvFnzt8Yqy2
596LGr9fVr8v+7oT7HMZ4bRKQ+FSW/ud/YKczdQHqXHRlC30IS2zrxdRdOSGUzG8cyOWsX5aCn/u
8WDb9wq2YTaloZjJy6rOJa+TgFL9gPAcJGzSY/9R0pe53DBEfl1b8VJhXG0vxE9syfoClLPjftn/
JY1aZ5N0/krwS/a0gKcki3PdyXGuM8mjgOFnGWnoAbxfGZIG3730KkKEzyZVC79QUAHyS0qOyoAE
CrhfPPMX/Ah3nW8RccF+BVWwXuLKopaNICniyxT5cfIYqXQ2uafsEvkoNou+H+o9t48ml1sQqjWE
ZUdhzHXxSefySIWizls5el8OXZ9MsOnFe/QfTJ7aNij4tXnNEY9AD4NJ3b9Zgiw/YtQKKUZuJQpV
4gCx2AkLnXBIDbwYpsdFu78ZP3wOX3+OOvxqd0+m3yOVUF/NUKkPyoEHBa8NhxL1K/BzaKC/RmJi
UfbFtjbEbKRWDXdEQwukPaPFckIewO0tBVA7WL5d97e2j0/t0R/gADQEd5r3jJchdSk0MdMDYP1b
RTUzgzvTD44BuRyN15/4P+Mcl6HZA0jSJry+HQRWOWlVnNbnGaEskUfJE/l1+Pl1nePmTrAU7TlM
k+dD1xP1CJvc8doJoXKXgf4LX5pZXTnoLooSQI+Burl4tVHwfAaPIltPNGhVqZqdy3kWc9E1Hg2J
rUhz8NvIAOfsE8iirvn0W1B/sTlXmhtiG4YJDBoCtyrwizvwbsCm4GvYMjZai9RgUai54WfdkvRl
EjedHbhaiN76TF0WmKhDTu1+d+mLd3+XxdTnsfQD9Kdsk3+h/gpPgNnG8eni1oh2RZMpLdELZovk
miNlzDkudTFgPj4Dmk329bTe9xdWrAzC0it2rYmMFO37nA6LIQ/1SjXN8StKMhjUut9hTC9Tqs81
sSgPEJHNaHFgDG8UnL5S+Ay4kebYh4W3KcpIsDh2BViPFlcPa7OrbJJWdIbD4x9Gk1pG/nzGNKnV
qhXKyqOrhZWVtUHLNf55JVxVAvWoqikVEAgVl1t18PmXLVuDAM1rA7+oxUwe0zOyUQXaVbBnvDf6
Hjv0VUb3T5Ri+kvNG54YH0fiWifH5orNdf/s+vNHisO8eRPXGEWwtyWd4Gx9NG9+KHSt7PGZtjUi
96MzGw+Q8ACp84yLF+l8Z68sa/vsgc5IR0OmBIyTAK/648MjWZj0c5QWg/y8YprNOIysVDZJu0Cd
Nbyh9z5cR0keZqDNFGr2/4EaBZLLrNPW/+DjE/CqgxuMP62+KHu7Pc1vik08hbMcAs3iz61iH7Dv
U8rkkf124S45nuPUAfxI+P6uAVqg7xSA70yifAd45IE3SpsCkaJD1USOi8TG/TTWnZCOne8TMq0b
hWfvlTeolsZMnXVn3KGRelv8MugtOXpOZlq2zNbIJJSjAuXkfmSYKyXH+Nd2YOchYjDPefqQgLSp
vq6ppO7H0epCxTzgQvClMvhj3w9Jeth37BAqd4FlPNhpHKswvkAU4FxhmdbspqVGhysTmUHBn05g
IHaz1u5KyJbIHf90JkkcNsSZtZdCQDzJBlNqXvbyD3InDe1qeEaBvCurz+scxg9ljEqiYvdA29ls
rHbPYsYHPxcN6Xg0R0lXJ0gPr5e8Ot1ffBUohejmr+tku6NoVBhd7pBdsr4bBQuOhw20pXzqDC8m
vCBs43NgmP6n3GyaSG8gEEAfjULzWtlg+23pfsQR4lmd1Cyb9r45hTjcrxkZi8jXRIwNwaujKfOt
ZyXV+xa6TXMn7SVclDMSQLeQCswGmFdlJzi0y4RXtc1Nwq/FuDKlHjEU4PGKmkM8WdJLv/m7vg+b
MnUrduIUR9wAAyKePQIlY2X8ZTAuP3gXp7j12mlg1zAgbQQn5VZCvCR090QfS5GKlqqzfS6nhvRv
RQSzFx2rnZQyDlC+5fsXc/0614re/WulhFLgpBuiB2Scc3DioDAMkh3D8S/DtroHp9EDS2tqz/dn
LFJFEPhYywYILNv7+89h/r7g3dQK7hostohNwMHUCledqrKrcMQdvcNqasfzuWF0L/Xv2mzsZV+d
zykhQgqJ76ib2H20KYjAcvTZTAb20uDOfCtuIazNC/OK1H5lhclXf//VI4aOBeUAKNCsD4c3Zmhr
d41kOKJj4TG9AJGhmDvLlDLqloQErbK7Me17WmKF0+wIi7kEdeeVL/jeFTM3QBMDmnICF8JaA/F5
91QP1v1o1Wwchj8C/K6AM8Y+2swueA5sjMrQNRi2WGER9u7xVkOvAHW1XOMlVjq30f1O7d1RBKjb
TczzWFPLgpKtXjRrxlmLusY4k2hXpZI9pi7lnN1oc0eTyCc0+0aOM5NWjkj6v/7/Mbhh52T8i5K9
WP12l9WobXB/rM1oOJPVOwtlJOa79Tj27bZP5QUqDo/8ejjxk4ZR8DzQCyzV1zq0a5zKaGuLXCd8
YAMZJdBrS1LKs5OyyilMYodgKS5F720G2NBaiZVPb/Yh9vh0KiTS0U3KPI9+LcrYo0Prrq8K5Ybx
nKTvWk3b4ZGMgKhXYqBsMupiWJTwulq3VbDp6VlGanVRZp67tuCNH5pst7t8arcjvDPx8jPV9t9Y
ob9bOQu4QvowPJxtniYKTOasTqCBvptZhtM/czcaaLc3sHNyw/O01D6PHykKBHW7ykHYkr352YlE
+XwoS8XbD2pCVSxxe4m3iskfA/qyf9K/qKuBdTE2DWUu4QbEW1akhDarm9/W6HKYe07lrehhYqzx
g029krAruARuE31S+h8PdGJ+6QI+a2IT3AQz5EmYLAG10f4OVOGMaFiRGo5cjUH6dVfYmnBBsgcY
6Nlu0V3C5aPvylp6rQYZLEZr9SLYM1dfy/VG6d31Hl92flnV15zeOl36U1a+wRfayQGnbXltR1bf
XzcGqcxb0C20XE0HZghFzl4qVnKNSYBfpolBUShcUVwH/QkYOAvTunAqXFInoL7TgWxC2O3z69Wk
tfwwolUqGVt3aQIalc+szbULs9/9lAY9ukV6HM0U3cfiwrqk0dhDCgSk/ZPoG3Y5SrBo6IZTZSdI
sl66sHGk7A7gecKElOaMt0ykM5z4JftAzN7d8h1OMAtV1NGDKG74Ln+Rygo+Ohz1ZbXfFKQ1qo1t
mErUuAra66EoxkO8cQ5gUVyeXGZY+ITJc8EkAzZedsmTz3O2dKLDPcclMSZDD2VKYUjvUFcgYcch
+o/cc7G1Zp5Qj/TZVhILm5l/IHJasVhCYDeffLcGuiGVYTrZssjGRMM8Z93XW88OGFa0GHjeDMcy
6aJ3HMnQHO/lXABN+wlv8R2au9IGAp0BCBnRRuHHqvL4YoVnDClhaN6zWg7/KfXcVumrSWieC2Qr
Rmgvy1Cb0VHIGmkpBbFDj7boUKD2KJjtha00OHyypDQE3iogqKNAV5DzhySNnRs1jmvMYv+DQXtN
Didy+/fXgCjT7rpMJzDJBvryZrkXLEU31lNeY7oJCXyUMc94k6vt2ufuMFpscf53/g+ZVRkYmUxj
d50h35bP0psQYMxNqiGoD0Mym27w9fqLc6rZRf5QTubFW25kuQWkURxgxFSgfGA8UARFVXLQj5gV
bXJyiU16hE9EdIsPCBIi6UBQQFv9hTfsX4NoVwOm0JZZXJbLi/RyRM7oVzuGhoQ0UDqAeFV6Mllp
puGrgu/YLJiWC/v/JZoOs3GpXKTwsP2uIGV32oLbHao/h53dwlz1OAFcVEdqQgRqP/mIKlTqpSCc
dtt/1cqnGn2Yb2Fy54woft/2fSmjgsHmSmm8fzQi6+u7TemIZvsAnLq3De5G5dSKjy9h1Nfr1hbK
lKntG7m0pvIx0hoS091foKG7AufElMpi+cPsKRO4kY2pNWxtQcrvX2rLyFOx2fu+GYSxogTdlv0L
aa9812VDTS6Us2KFudYQ77bBi8ZJus/DD1w1O3AA8Aoeshm0Oq/3UOFZWa4J+kWAWmWUy44ZKxAu
EMW3z4VHmx47DjwRVDbXrS4Ym2dw74D2tUUbcDjaNHFEEcZehhAPNMQBDvv5LTtSDe4shK6xQBsC
JqNIKQ8/Z0ZbPtuOipHQT7NkYeeCNKu2X08qbRenCemTW83ZTcKSDVUBSsHzyykAm1YMdtRkgzgE
qyuFpf6yCofc9eNGqM6uIppUSKH85VhExBelaBKwnd2rDZi2xS3/jq6Kd2y2yogjEPADk0ZGcIZ6
QejQDmnrpEHjxSktuhQUk1mRgaHElrwl95JElxWf9OGopsLbsFz18lL5WtIZCw7G4JdTBJMx5nXo
ZReH/T9KBKnXwdftQSBzJBUaZOZc6ri3hYmp5PWBeSm1v5hN/FBTdoIqrnofZH8OURunwhdi7xvc
LoJcnpuAof2+pIvzqk0u9qQ67I7wlksJFlfoNbQmUOyUR6OJeh75DmDxC253O1DbgpkIpxOlvEcM
5BuGRkeJwr+gGIlInDdlL1/+sv7KMOG7t9kL1C5wUHpQyVasGA5D+9eZ9pudxsMAUtx6pU4vnq8G
Az2iT2KXcyiicY3hCYTRyB8DL1PuRldnGlelkEIa5kV5sSA4KHkxvw86hbnUg3dSqPrYendIV65O
8iccvOFmlOtbNhkL0eWFhOKKy5Mmj9ar8Z9rTlNNqtZmrqcJq6sMNvDJRbABj7MPBYiUy+qw03yQ
4JYq3R9NIMn5gaHqQ9cTvlqErhWQ1hAwj/3JnssQyezItilICrzWY6fg98lG36KkxQAkFIV8VOBA
j3PJyYnGDgobpPfILR/L4ROnJ4XR71W41HwYsKLsZXRvBpx6T4/xLDBr9t9jw454sGcqWlEpwIEi
6skXOc9IljZv8xPpFA3/XdUiCpeO8u2RXvQ2LHioEKfsrExAG+Wqjo9NhtrKY9Pw646VoI6U3+Pw
mUORD6uPciYj2xbpA3IXCVTACXtXuNIaqgXiCcXUZ5eLtX9xobSmuqRiPr/KaQ1m+7ToHGsZZhle
xQXPPoeljYaH+GbHCmcDiIflCgIXvnM3/NqgOWJSdcwU2s0F96b/hLCSu1QqPWpkSJQZA9mScvTW
tD2pN8ohLq91WhRKTERFsFx9JlcyToBqzzKffZSNZhK31z18kJUG0+Ihcjzy6uKDy1Qd7sKrC4kl
gzJQwXjMkV/4ppbTGew+me/1f++/+Ml752hpZ6UhscqJ+3FVbc+lscAp2c+FVhXb0xYO1ewbALoc
oGLIqKp2JmjCC7cNdT4arq3b6jrRJ6nIxRe2jzZkDICBgU83YfkM5SWzDVyv3Ws1f9FSA1lhne/m
Jg4zVpeOYrITmkJ/fx3NcgeJF2DlMl+AbSEiOucFx8AfucuQmCO9awhIOmZp4Mg0f/UpRxIj+2gS
pWKK9pRSRd9/QR9gPKXJTAnUcaPrax2ohPdheRiCt5EUmxQgQl/SCO1wMF1PdAZ9O1ynrqO+KA+f
bgGrLDJ67XZb5igDywMJw7NCqrvPpUhFLuyYl0T1ADlqk7mdNuwnIxVp0JSRyskN/McHE5dU+WKV
ZILglNLrFR/mFIoFPP8Sy63g2WR9NoW8aZ5y5V3NbQvMG7CJlBLJOLdGOIJ0/AKsSR4Qlkmo7Sak
7dgTr4jUPWkq0qo4Hjb6Lm5bVLVXoeS0WIbE2Ez5lEkDxkUip3Zn98E6AbMT1t3MuGgmdW9jj4nn
Gb6ZY2dHTNsBEwWiHS7XAlpQZSEMXKtwtWKSwgirW/3KcLiQw7AmXleS6SnunQdMr+c/+kGFy1YG
1Mz9wDrDsl0Ro/Q+J/dX9uopbBCtdfLKBOoNv0QBd6hXpSfRZpJ1U6Q0tAcdL3D8/b9vP3LcHZDV
gvXyKctOTwU4bICsjQmBqKCmV07Alu5WLSUkVEeoN5ZeZh2C7Jk+J0Hxrj8bx909NF5Fsv7v3wLM
zJC6hVwtp8ybQ85yoO5VbRCVdEKw7ntoiEEvzByYrq6QYDaGf8OCFO02aLOB6jnA96/mWrypnayj
UNIdAcwcKXpthySLoPiv3xog/2pbFyrVPJvqUei1ehb96OMlj4+uzhCOXTwADAwp37FRoNBzTinP
9micTZnlFuFwS3ud/RfSPm5AtXOH70jra2Qo47I/JgmC+5HhuZ5RDT/FY8ZXvKQGRMGaK4558za7
JBI0W3YGwQt9Pc1N5asIa9jmeYC98GPxWf+LLjvah19SZI1jGjiDGNlSAnC4Ywl6lTRcZ5jYFNrJ
hv+IFt5/VO4Gn/pbFlzUa+gTQMY61aRh59s0Jmj+sf15GJSlLDiEWbfa4gkRpDyNjBfR1cpnzANR
W8lTBLA2W02xYKpGDyexnLnkug9VN9ldXoH/OLo0LLOKGrJb2OcIkRxH9e9MjY+xlU5G8Ze6S9SO
k9u4uux1NQMe5NckW8C4MKs+k14D9IrYS4ANCON0kEGtDF5TcMFz9BX0MjrVO/aDljcTrqONLgRB
PKUovYLT8rJNNa+WYci6yTcTw7anIkqKTKJ1FXHZiC92516zbKGbVwRRAwwlToiDG8jcK/E8yqW7
ro3ABwXcmHQ2ZlCVDWYtaRNt2attbgPK7j5zXSi+lpXtN9ITJT+Wt/uUBeRX8FTAseudITu0SN+m
yeIW/Gg7TNE++JMvTJrRAUvnw933XnbZRKu9uRYTPcOt8Zvn/0SqpI5T5ZnlfFmIFL3DEqNxqrvT
tFvDS1UfOL9XqIfGNVs2PjzX5wUfWl0IC+4b6JaltGZiksMFq+HOky+JlGL+JXnIwUQMj0Yk3yzM
Ak85KkaDSu2Lg6qXNd2GXFtYWc4R2Kh171X+iKl+gbBaKEu32WQCrdk2GBB9yWReoJtcP0jbDk+0
xcr34msI+oIdlno70y0nKWRZxbfU6B04bTVMjr0M+wUQfajfMAYK7pHCeKwgjl8NSD3c6XgBd6z1
wusBTh0Yv60FRkIn367McQtdSDvyMbZrj+XRs5wey1QkbMOqye54TU62wGs7no74uinnwfDlRR2f
NEQXb03fTonCHO3vAM8gIWlexAKk+eA1YYUFaD1EqmVBGuJBLZANpZ5+JszD4s2Yobb+bkEkqfxg
ziJfg7DTbDc6whsacOjxuoTrpN7W6zP3YIp9CwWRyNf56M83x2ZFRRjpW6HgbGIpGWVck6DK527j
xhfK9Tn4hxAjfLGIiC518RrT9PJZlW31jt5lMLAlUOUtgAOgj0q3KSEVM+9tE0bYTG9tW9rdcPdX
8ApkG7v4scNc/IpwRlb9l1c6kXaRqlQUABQG2fYJNrFHhAPkkEkLUHuYoD8bNfZTng+MGC/Bz+8D
I63GnLJwpPbH3MJqoBeaIbfQCDh1HPvMcKcPkykAm3VxfZ+FIn3pEkXonEgGIoo8Ie+v32SMQaUs
eQrFqSGnFs0KiITzJPaCR94JLA+/xI2uY5TAq0Sbhy5nERdgSB52Y4WUKiTxT0GkvZ943G0DyBtW
kIKDrSAgv+kCRHyY/IwmKEeK/9Ba+nkzGHzA5TR+zbQq62KcxS5ORWTpO/EQ6PZkSiHBK3LPROjp
44WRjKpY3Ajl0uGpXY+ILBzD4C4hL0DDThBo2b7nVfN+YAM1fXryVFoxVZenkn2cuGpMcpHdMCtW
ZEwDCWeKrAk6cX5T5UcIGmS5KqYzBgMUc2P+R3PbFbI+g7kIAuDQgRzZN4G9wMYEUExcjuJrW1dy
WszvjMZsoVDqU31nNl88t2jDmKHP+cZTFIomLLkHIbOVRQEES5/x9dbxpnCyLWSqsOik4kjK55Qf
YVopWQHIFEITjxTC+cN6I/JUwRmsfOWLctGBD9g3nrFSm6otx07kBwcyGkYBIoqmNfnNwdeZrp67
1bbUHTMv5xO+/5aPWdlBRklLXe5rgIYJrFqSG8v0Ny9NgoqR6AbaOHxsRxiCkvMMADcRN1zamUfw
DBysoVTk9kHMolYbl8lEoD2wLnI5wTuXuwJ6VFVELXsl0UbsGOOvko5yGcqO9MZ5m4OVOBZB5ys2
CiUnjzocdCeZPs8IHL5lldwSKHgXcwlZTbPkzcGGoumVj5wvVRLSSUKuwoSGhZb5VrycbjjTBz/t
jBMQR9/CMnEHsz7h7iv1jYmdAN69TcPZMo+5jgU5DTiyLhanH0IbnrMjNwNaaLG+2+JBnU1KqGdL
FdrBs39xxIID5a6aI2PKzz9Y/te+GTNdLnC7TgD2UdTkEF74beiKl+TNQGmWlF+ZW7wDYnrHoEN+
07zBwRcDYhlxrfSXLyjgLosTLG9tmA/+K2p3/EZTodmq6oLCnDahmSYIqL9YZ4ZyDPlrp5jMRSNp
QrGhESOiVhHgIW8Zu/vgZQBuR7pt7t/iPaPk1KhXSx/RMfsYPELa2bme2QUr9ay+gHznILzqkATb
JVIOahewRYMU10wjYSvQz3U2QdQr0KRYZg9HNmOki02KJ3p0ITrh9cit0aq9T0v+yLlgrBeAY/ay
5B3j5XKnyDsZQJGrOW1I7l5iOit9Kx3DG0ix80K9t6PIxu9xr3XrNOUyymYhQ7S0++8lQE84+cNQ
x79hxtB3bSH7ofQoAQElLqe36x88vDTRuLGRhytEaDlxJDt276xs/7dZDwAHjjrYxGI2n1IHc09C
whGdERlYEyyn4Fh3fuIYozKaiQvguPo7VmYRVuyUPMH1/aqWwWuz1t6JnD8fGozotEw/f4qsh5jB
OavSSWvDOGl1IOg0sxDZ1VYlHf0HD2fviXexle1le25YiuEmX/DMb2QKrcVn/apK7xEom73QJoDS
jihC53G1AxtXP5EonGfis0axCEYELl5k1XQw8MC+8DSawc8+G26+HAGdH/ulsKFE7sno02z9H26e
kopDEan+P9BLRYyVURSnGcy4NKzt8HRYszstsb9PTCGAs0XOiTuLWIJgflKRdnMUZtCXTKkSwvKU
0OC9XpTZfvn63SEJkJJAGWdC1LEypSfVYXSxxzxKDs6y6qSQ0BffFHsrS3gFbz6EoUo9RHV+N9Zx
+5ax7YE7spXb3YIyjfKkLMS+9lUTQ4MXBFIkIzUFRcd9ixWmC41NGUiY0dTeHOWgUCoox6DN7A84
b9c936HGPery16QlclODryQdSOYkQxLkrWiDrdpHVvOW2dbvQtM/lZVKg+aQXpL56X1gLhlIh50h
JZ5vbrIjxiUhn5rUYYWJvKzbeDVPxz9bGAvWznsjCjAiaaozoj81BFYU6bZBSuSKhn7jN/C2poiZ
uraJpFt6CaAv3Ul3wrbo0TfbZw2eW2JAkiOYSzP+kVbUSM1YDp4acjjMG/DzUdpqIFHmmik2tpu0
RRD8jOgQOzdqkxcTN4lfYh6hEqkYtuQvfJm9gtWFuFyHkT/VfQ5aRBmDtwS42+jZ0FDCG6SupsGc
RZGy9qbugi6IsEsiMbJD4LO1Lk4yfwJMzm/sW+W5hq3PF3b7wqBbzNY9SDlZeB2cD3uVYljT4uMn
Xfg2LzzShlZEnzZd0HIvG17j9tu2LX4GiIwKFp7vvmZMNWTHJ/b0Z2qs+y14rwyjKWgcu7NyXcOD
0IiYNEpb8g3hsX7l/khLvDUcEYiU+bLOOZA3MeKzrSxsAfOaxAAfW1SGO4VXCLRkwrAQB8K1XpdA
YNJxj7Gmrpu0wHZZ6/Ak60fBXd0ta3UiDY0mjHFX7BkQEEjh9+Tr55htKJ/aX6ObsZ3UTtWHHoDM
cwmup6V2RHzIf2xizke+rT616+estyU4gNWc6G0lxPVPQ7z7VBtoTY3RtaCowpyAP9v3BOoMQkNl
cZ6ISsf0wGvfT1YCCeH98o0XM+34I1sSE/SkJ5q1K6Migc9To5/+yqxcsDnUKESZgD1EgUchYozI
IQmnSvSSaR+uErVdbk/bbk0evQlHT8dTbytv3xJr81KmwRj9/pCwCJFqfRvZrJ6bkADD0FIDxTcx
Q1qMDkHABt+bOKiQ97ztkMI3wF69WUx1rYGjiTRZM098HcnEbLA317poNKQooscUh8tEXZAXQsdq
WSmuNlaRDQnDKM76GH0m8rOcNLd1ejifBCJY24QoskSRad97Qtgo8OoFoJAK7Bejxag9DDy/JzTT
5DRKbjnnL1U2cS34QUWmpCdt6T4FFgqnXXgxVSSSnWLimqe+30Apw84SphCI3Tan8PBm7SuOmdV2
muk8Uqm8exyeeH2XBh0QtRc1BcLzextUNq2+gp9W7dbkwz9jNos6wKjbRh8uDpxJp9Nzcj8ILWvS
uWoTMcV9JZfzLncO/1C69OQZeM3l9hu4+/LFsCaK9x549NbnLo+YQa+xW/GCYrD7WMLm19Keczc4
gVKzRqJPAASLXCqLoM/7gu8nl1LcurnK5afb1TqhIBnLodV2RoygtebRBZQA7VcuQSZuqxxlOW/R
+6FNqJGcPl8nyh0pMIxDhCp07NwvijR9x/BtQ5rm/HM7QnZSYJ7d8FjPuTzA13u56oY8oIV1jWoO
mEitSID7lBdLH1wlpMZL8q+JuEId9MYEhJTF6nPH34nT/55YGKTCjrW01L6TAyNHKiA1eQuUM8ui
Jwx4YoZ3CODGjHDEVvEAkj9VVEHuZ0kT2ID07Oa7MFvaO2/qtQz3GREw8MwwRutSKefycfhWqclk
hDS0x6sU7o7XPkgZbARMiL5pqDi6fPrqXNbe0D6a3geoiZ18aVk2zlxMhpfuPWa9e691AyaNsC72
/yeINMdjJdMSpYo5R251vEF9U+jc1iYyowBJCNHVMSHgtYb2l3CW2BxbwCYqUDBHiO9qGpDgYoKC
e0HaCnlcnRaDEsJxU7iTfWHWKsQEPdfO0fNqg+beJrvEO8oeu0COIK01jdkKS9wwQ0TmpOJS53JF
LTBEkjZvuLV5y61vI/WqrHSuLYhOfDzUy7tMcytWL+gxru/kqgOwMD7+DkBNSA/lepFpXqVkxeGZ
FhWebbtK/Ee7leCMisabltNjqON/EBazNS5stCpo4Kq0Ox49iJamfLl/6WbLtuzQBCwdMb9yHg7L
eZvPkJKTXch2U+toF6XITNT04fWa2NdvRzArF/UdHsKQ/Uezen/0CyklATKE7IwN47MrQl5g+btI
00PAdLcJkqxK4y8acb5AQLZnBkQEFCvqmjunyoFUBb1wk2C0jBaNQF7sx0fIETFrNmVMhHp7GCCF
rD1EC9qDWQrhOV/PBmLimpRhbew3ykslaNtv8rjElR9pcX9HZ1YKJut6Vkdd6FZdUGnz7rTgBLIX
LhaaX5vafvPEm2++Ampwqp53K65G8PMImiap4eCSJ3+nh+B24MYEb5ChueuIyFhDIMuat4s4FQlz
wWqLpo6zpmjxUmuVxyUMUk8mwbla0JJ+cc3welw3F3E3yTH459CwlSGYAijSuHitLX9TmhVf3Qfx
UW7HSTmzu0RILJ2WsrDC40y/sJIJpy0ugKN7xrfhQi8equnc/UpeAb/CgbfgvSeeMjcL28Q3KU2k
J/y8rfKaHgFIssCTG+8gsHEGH4pqb7hYZK026+t+HJuvL1HGD6tmaIsQKQUWryXngLV8LBUmEjTA
G8FpB6V+AlnQbcMCyXhXSq3dwuHmT00h+X7pxOYBknY3iXGU1a9I3wXKuul9rWk7i3PVaGKfb+pN
FQItP9bk/AEbXMBj33Z2BDLSG+291lfkzV/zXsImCVh51U6iXnsYY4Zsvu+qLu59F0OXhWiPPXVf
RDiXmhnbIYuF8rEMvJR+Z4WO1Ndrhlf9IphBFBIWuMkEtvnpBjC8S2kUbUvGV/1DYDy8GfjkZVHP
bde8PMFE6dHmYWr5UciNyYiUumbh2zAlu3n2Wx1H7bYeIKUu/Wdh0dqwI2XcqlP12orOLIjjwfJi
OaNf2Q6eSzk69gRQWq5uzlsqE8RR/V2O1Rwi9mx/fOA/NPphlLsDgt2r/aiTOVHNgReeDNBpwQHd
4bMRL7WnmuWG7tCmn+Utj1lM0G5cKZcfOjYAhMFSIyWXnxgl3WezrE6K8bEbEMz0BOMMgc8wL4Ke
Dx7EzEaqisMA5het6tTWhiFRtiZ0RzuuDZ+D0XRPKl1T5glgEK9Yju5g4FAK8gyyOZGIC1M3j/X/
2XmD6asTTaKtvoekANvDNuxcNSWylBKNRhy6B+PeROTvKyk2D83lEpOxasLNCpEOP/klfHDiGnsX
uedvZOr88LqVqxTdbC9G1489GzCuzDq1MAkMoVF4ysZotGVoVDjRiisTELhltpzvZMNUEqnyYdzi
2pg0eHGPg7/CEoyYX2UeKDoGsMqu5hyjytjxX7z5eKWRAcBWOpUXE/mFxXh0hJe0uzId+wVLFfHc
wLHs2Coehqo8p7yhE4s46oHazDsJNlNihXuE9J8Q+FdLnruBTxLjyCQX0LgP2w6rQsdpAm9VT3kr
dFlKgtnIHOQ9793Mv6q5HrxCUXGuk+OJzTEhwiWKCbxttko0QdpRoAdIhhZScX1Y4tMZjF6quVzC
qvcHn4E/LBcgw5+xZib1gRzKovxVJfkoLrRE7mIgyB6x9xxbXBUhJWkR8S7zYjmasMyBkLmUW2pO
WV1kRkwj20/VsTR5xO9Gza6DeqpKmfN4jZgNlWYQBBbrK990z1Wc0w0fVDRqj0EJcjHofBWJXaDQ
hoCMffjNDKRviyry+YF6lyzQryd11keoEkhAa6Wf3Iyml89b3KL1nrVSUtc2X59S2l4fj7yDckFc
kdwaNeN8dRIlqc+HBG/R/nLWJMer94lmmIdvRmXVp+VESKvauFhcO45WaoMZFW1zsTg3kkYl/5Hc
OMcMMe7g06Yry8zBOdgRfIAO5egFKaagk14x5qdZrTElyKJU3yOUigfMzEXp4dgfEA7f/kksp8iB
ust8vQTUgR3AYQ5+HG/fPp7zL45in6G+FnnTr6ucbF7VZLQJtwv7G2Ehmw5pTlJ5uZm5I//msUkr
IKI0hZ6a1HGWtzhEvnbQdvTvX0rrQ2+PVeK3wDNTArZrfaCvyK0wHvW44OKZ1p5+hhsetceUhraG
1Zkno8X3W/7WGJtnTfCr/RPp5T1msHO6p8+dYJxvk95QvPLrAyG7QF2MjVxFzZ9ermICzqu7/3Lc
YwWm4jeDgTAWs1gjSU8i7fXDf/KYEYX+hpV2RsZkBedPmq2Z40cd/v8K0OTpKx7bDI6FrcrkmTgd
NYDzKE0U/tx/v4jqow7MFrKzlf/cPT87S07VRpkQLxmGvSggdzLdO7zIBcmXN6x5i1obBlCRwug6
HT7FlFYuKd/GSAwThWsS0gYGcVIk94ox8F0HrH6hYdn8muGXxxg2HoZvaEjdUQgJ5nXLkgg5nMCO
dAXGyRUF961b1hxFHi2xuJRFuRqHoKz28ax3bo4oh6tWAYN38BbdYamUC7ZN2FQBtwas7KUnlB2z
pOldfY8n/nkl6ayKTwmJG981bvnVBAi2qFOVnC+vuOf1AexZbKG+rZSLNQLOdjTFqiG5rD/uNKb0
iiutZyFADli9Hpc/znKrsYXDRA4b3Hjx0nn4vw9awqmN1m0kieQzSodWnBwID88ZsFx16z4whOSN
uM60LSdXbTM4k+q5xnRrLuvxVpmy1wYgH6PEsIlGo7mE0Y62VC/XGHTvuf/W8RDzxlcf6aOS+oll
FlRc+NxU6fHBojrXRmzTMyA1o7F3B7QfQ4XltOK57ncY35K3rNLp+UWuII/c2fDd3oliD/6LD/zD
XkZeDFzUsjJ3EPlCuLN7+/UuKcdIh5sk2W3bXWIWQBYnNwkW1E7BClUvckj7+pG+NfORC7l2Bn8L
5WDjWTjTYGSHALRhhpM0V+4lhU/K+/ROujOWQzFLlP/Qw6KlD/QZTW7ILQavLSCp1KHtbnwT1oke
Zcf8o4xL/vH86ITs9/sk5zyuLkj1/sh3HUzYJvNxpjlMd7j298yX7WJLDl04TwYGRkUX1DnXojaD
JjgdDgh9oP50xipl8jrLvLQgPV+MSgQo4JTNbrKbxK0tY12F9BZnXXHQaV3G8pRp5o3coIQKUX0S
w/iH1UDg+hYE6Ki7aLFt2o4PIRPU/BVH6EPTOzV6cskWf9u36k5UHcOkZIj1fkRrg4oJNjQnWI6y
pZ+9c7+NDq4k1CWgEnD39s9302sekB6DzPXGG/4Qr+CGm/OXh/0Ks+2ji5dFyi4B18qTkRrxd3xa
zQv0eOisexFto2iSus0yDD/AH+KXiB95eXULNPk7ty28FBg2qtugcvfN1jDJY76LR69UsUD88qh8
H1XuoLbHAGmZw+/tjpALwoUN7DNyyXi6U3gtwtVzBkQXqoKgn5a5FaNTnJuDxZdqKJiNR4mcUvZU
kUfKT+jSfrSyxr3P9bZD3Puy7GP+zJwiI+5mSdWu5bQaqh6Kc/57tFVuC8b/eZJO4Fxn4XtV9MDx
WVC6u3jyYYHjgmrciFpUB1KKHVsCIjTkkpX+LvVp/O4auTnuCTV8yL2X+GxmaoZBms6DMV8LlPyl
oljMw2bTTZluOJuElC2Wzv78520b9cgtbLHZmHdcDjZ5+cxkv7VRVXUp38J1TeWWI2uxjcRly5ku
fyYrZ27eShYKDL8mUf5BhCgNyf/P04BGE50jvvluF6YN+shFbj+Roi5eIwmZigQ28wLpM/4zXhLC
+Z331b7FH3Z8gC/d/kww9kx3AMZ4us8R+CW058VFrS3mEyENlZsq+gRRAqblz/+WxRiVVuns5udj
LdKbliiyJ9YTsTy/wbHTfeAOhiWqSBBlLjLtstTVwG7fkAO90fhk6YIU8qePVO15bL25a0bKu5/1
0NBxC3eBt2508tYYDhDbFEfRglzp9ndlFY0cYMAq1yX9bSkjmrvuWS9CObS3Xss3c5YF+PWkXO7V
5FrbvgNH+owdy3XMY8sfdDt/92tQhGEy75QYm+HbcTccd3L3dLvE+9xQKYOUoBGARoxNejuxS1FF
UadetxyYchVCi+xQtyZXFvdQD4hMu9osD38+6SrXnH3Ubc5Uu/3v/pxrgFS2Qct6Gs+Li+XLSiJK
QxQvnoTzjpCa0zI3jsGbN8zVjepCLEuc8Acx3fXQZ1lhQuP7SJugZX5dNs/GNSq0FMvwu5JISk0o
aCy0v8qPDxYkgYzqxA3dxtQds1wgErNa5Ri5hMjq0e/LYBV5u/f/dJbwt8kYzcHgJgNJKGsCgBAR
vbFi7WxwWUhaYv+EMkStZ31eD3x4JJgkb2CYY/3JT+LprcqNs4QGskkreRveTC3BhpZh8bldnYB7
PtL7opzcPBrTtb1DOJcmkZutW9Z2yV5pA61+qsJGAyNvSTZQxXKnpFnjBC4hQ5Cu+dChzrlBFRn2
XnUwOhm0F0p91adwhnK739j7HsOWtBIRu1fRpmgA8eNzhQvotcFOJJMW31YoIZXTcj4stx2naNXj
gL4IJHKB8tAENaYEzbi4eVfX8YqucTGVZ/n7xKRzErIK5Ciu8kdzZuxoHSlyz7lJH4mpMmSEekiT
NgdxTfgZXqfAlW8ejdh6c3Bq9fCU6kgZSz+4IavplIDNpkHPN3+hnj7MN6wjhOwOe499JNGWYFDq
aOAfUjimoa40KlEtAA20BLj0Qw7BWRLkasLtqaTiJ7Tw8v6A+AukDjf7oRatU7u1pg6ffeDEppke
UHdU9mV7synt2cgLsilck9xOVGQIOHMJjwWcSGqnisgk2LlCtCgoMuZoZcKqzMbP2XDeWfCJkI2R
rjcIKh05ks1XyiQpZfEapLfLGHi7kpeZ8FXDGUfUouCXgwwMWytWB5Fsp7mMTL/Qy1OXLMCIapCJ
+jCoqa4v+XMU4TEtCjKwlV/S0oUPCeXBiu6T7nGrg/Q48ZDT4UsN3LrVMO//+nuQSIlCiiIjVxhP
DMujKWQJCzFqPPYX3xd0bI48E9DRm9rZeSaJe7KsSjex/rO6kl5y+ICt+extGS4qWtent0zO6Xlp
GK87Od/UFv3PBJ0EEPFNT0SAmeOAE6sjcFlyylvttE8CYo6TJi+Fr+ZAqHwhriY1x+VT1zKMPaND
gVErRWh1LjSZzfovi8zDoxWhqa8cvj62KjwGd4X9MwiUsC+FarNg2QJGLDnOzDbh9J+cpEEYO5bF
WAtEOvFcTu7h6BJOn8J/dUMp2sbuTBKPpb9zS9sGzKKNGtTvyFD1rEb16jVNZmCaH92+6SLwDY3B
0/RT1HL3RF84C887hr27ltsMz002ifZJdbnjG5VSe3Rf9HIuxkNMLoqNgihRFjwmWWoOi+Nwj4DQ
UZEnKdBNWt6/t+QhMx8/Pft2EihD1tquH2KWwTHt3l/K4AmtjVx7T8sgk79cVUv2bzu4mjySrDN3
aR7D3GdfAQyDQyAFxuMNRVfwazk/YcuOTG5AZ90Sy5B/SrgK0dHKQdcEbJr1uw5VeupLgcYnLTJ/
G1jRnPk4CCny9pCS4SBAQdgpX4chFUFON2sT6wb69UUcW6wuSYI2KaYOBvboXUP4yy5rDdv73LWu
o9pOfj759+yCbgfTUHFaN1bTwq4EluCVuMWzm6TP7cc9yW/KmXgnHyux+LCzEhgkyQ89iVrEmp1o
tqzuZb71eDtQqNuvqT+uRgyqw8j6qDW/ThIqGMoxqlAkEYvpjwf8JDUj+coD5EDOYvmBNnZydXfw
nnG0eqSH6LZXkkR6zLK5p76/NMZi1ZyuT6er7ZWUkYFbtl87BkkZ5ucPkHamDkJeQdGK37Bzf+ib
IcDfbX4WAsAqqKJV9pnKnTkl8Fi+t7WUrgsvHQaicnVo1iex2NwT1UOKzQqBRfqgw2GjOQ/dReGQ
iFAWdF9bkCt93KhYfTGqyxwOIQUuHRh78E8sa1KERVbZXUXVXODes1MvCrAa7237CQHhnZ/+g3cf
XJ6JoJBrFxZsjgSSXQf+uUsZVCk7tIMqD+P+e1QcQsujwZY9Q4y653oWY69iiBTGFSzMzCkNXOq2
XJODhqQfuIFBYRZQ2N9lRUne6nDt8SfC0+la0BitGsPnkBRDeYgx1z0LDDj9F21Apjmsyhdd79jq
QoCwrMpLG9OwlNBc3NbfTv4HZz4DWJrdvk75yfmFv2ootibonmuFjqIJOMPGrRhqswFoLK36MCWP
OMlqZcb/FJrAryChWkuW69hJL5oSdXkajl4flUPFoDlpEoWDpl4NL8sKGLyDom/go5AE7JeCQ3H9
/1ZAMdnTp2O11iYxKqkhqu+SY2WW2bMZ9alHj6SXpFHJMnS8I22fvb8eJyZXTVrI98ToKCTeLSrh
Apzndtbj1szyRZQgTtP8bIiXTcuuMmSMRjwvYEy24P66/wSvVOYpwr+vNbu+9SWwYGzKJkfUjfOe
ESh7vSt+XGsm+UROTdxO/ZOTcl/3WtKiWuYA+SMQzHgQxv0OB09VaxSRhk67hSWxetxi1w34pvoK
nDpZgR0ByhUi/Mce1bHE8utrMluXRC4Vn09ZDOJrQz78SZqs95i7tTIiAELY0eon3nBQyOQiTWYs
ZrVoA11tdQh9X0+z8XmreoVQdUPv+fJz12nqCGd+5JNL5dciHtRZfzHB97dMXWuMXyd6DOlQdzz6
D90p+PpRbxAAlEBtAGAVdRYLsd15XD5Kk/r0LaGax5B1bpsYTenBhDq/LNyhErQ7b6OhUNCG3IY+
4e0iYpXZO0hqePzlN8+Rbi2NzWq/kG+CRMM0tlEfgpzOMw2zZWq1WI/2UZve/IW3RTe7I3Kcmgyo
yFA8fXizBFFAiyS8ter1RVmJD+DPFZopdzX1AHsGC28oNhHu40mG2M0VM7kJJdpP50/8dN79AkP0
tvxEBqV6Yv45Za6J9ewS3VPZPTHpwpW+vX+RYI0Sj5CzHjBz9EXBQkC9V8deo9BxK9Y3YPV5jirR
ZtIqZ6/S5vR5sGvQqkOMj+hUv8Wl6Od7to/Fl/ka/yqQFXb2DQP3TBhctW5j2ZDLrk0yJ7hu40/4
STt7IwZBN9gWRjmGs4g+vT8Y9SG8bwnfM0Zd6nxHQmcsU924c48nEqu7Srv2ONy3bsn3+E3Z5f1e
2YB5wtiGwxZfnr66wJV5AodiMKxXGgsX4Yu1SvmL9xSzaGFPqYW2F1p1zAQ7HofQfgt1zI5nwvAP
eej0/IOhozefOMvPa99BO50XWITk3Vom5qTB+X3WMlyPHYTfOzKFWrRXTUbl9+1LJ+K03586w7xV
JHw1Q8butqbdcKM5t/uViODxA8G7ixMdHmpagahNQPzm6WwNPxnu9X1Gzwic1VdE7gUNl4oMu0K2
JCYUWxeAlvbFOUsgN4FG9DdZr5U6Ok+hSe7+aGK9DaRxgPFhzYT0N1cAdJRFu381xoyMgBauDTIJ
U8dJwrV/fxRmDoZGt/FCVT//GNQPBL9/+7dDYItDxAoVjINHPP6WVzgIfBkKVWqkUv5FuCAiX2OE
4SNQWFb/j9MgGPZzq6kuFWysddxaSmmNHljaZmQ656lklLh76J5YnlbklULRIC+uJW7OPLYDSiQm
CZyzf+rLQ7I18YUppM8FFtgJMvsNzu5+eh2OhZ6DeHCt18yIqBHkn1okLs+SwD6RPjDRZ2fH5od8
nJyrnLcZVXfoSVrIlpg89g5tqsRM59fSftDx7/VKnpef8pMmPKMVqwluLfDwisYpY9+vVZgiEuUc
6MAyGKTei93uSqGeabFi5ajqiAkT8HATvbehq3F+BX4YtvYFo03ESf0sEpNtp383KEVnkfkGKlpk
/tPEv+pKTJsB/nfvIX36TaTBFPdTUVIMDjoTKTU0YJ3nZ+BX7sY5zb0B4hPvaETMs1hclHOGLKiP
JbGs2fJ1Q7cHXegxWj/wYgeXbCIU7zVILcXA8HJdHIxNQ0xqybajlueXtP3EZ3RSsPucOuCLu25o
5Qju/fBxUFCaexZevBOkhMq7b5H1bsQHrzjpVVIwQbOxWzZ/Ti5IwG58+A2lkrxvUuPdq+Bx9t/b
bAKvsK/muVwZqSH6UbkjEi/zr1R6hR0Z0ye/QJyzPbkWKqIotWB90den+N+oAAXbP2ESHZ0liHVZ
75H3d8UQvNk+ij5Iz1ODRkk0aZxmg/D7n7RX6R9WK1QiVeZABEM/JSVW6SzS2vEd6DaVcWsrgjdX
XGBdSwpe6rP7zJwZZ9yqefGi23ob3AMCqmYCHovj8XhKnGMzdL+O1gU1rFnBYAj7+J2mf6i2IKNX
yC07Fzbs0Ts+rXWTc/bZfILVTzU+7rdBc2QP9IMwdRHM6NGf/+7l6wYa5Qr++pvOGKxpHWUeXxZR
OEBjE70ivMQDMVreMLpQTIYi8YcsOQDCUH+O2oM5eFV2iJ978cK3JEwTPY9FiGlQSuhpc764Rsmr
Z4L/lVjVFKjv43PpN+HI9fyPUcCJNK7tSQmK6XGopYF8Cq9QDCjnNzo0TMO9ddAkzEKxB9a9PvD2
98eC6F8czlUhOkX1CRmZ5kp7y1kh3vrtUKp1RTDaQC5+l7ZCDJQdf5ZhBTmbINIrjBZlBF9XuJ89
Hq0DjF7Wbtpfytc4cYAOEB6t7MArGlabrxNLDNI2gFivQWK2Xst+qSt/gKGlkUR8Z+e6EtDnOzCz
7kVupL08kY//mbhk51AEmamjSPu8lX86KTufwPlDl3SO5axl47BOaDnbeaDdh+nlq9gjwqf7EWrn
EpP/+gBtVZh2IIkqPlga7H58zAVaAc8HZyFX/XS2T7Fp/CgHfGhVIGkHwOqV2xnS2L+sB6R0AV0a
jefqGEMh0bMEODnktB8M5ue460jwYv06wwvoBeG/2fy+DwcFwhosrP+ns8E1I5uCKCM4HVHOGPhE
NctYV5RjzjTiQsPz189fHdlpDZNcBhNoIIp+sg9viQhybQQmoRT0sSokJalIcS6BepdQt5BsVZ/7
ibj5bgKiGlE9e+glPsDhgOb+Hqyk64PwYWaFiKjZqyW2NtIT3Lzte3SxklyGNv3u8jWrdxqNku+j
q7oG+5yPftcR4xRJrhExkSO6aNig5ZLHeyKjJFEbHDBKcpDb0tAxEU8FTB5n20sCaTheZiI3r/W2
krjiit+VELWe90nwJ4lqOxfjyJ0ndAhZfJ/mnh3QFEBX2QFui8DsPj8WCRrTpNIL7TKkdmcMaQat
uuIzpXrTpifx6X+FyXbvhiJ4u+xgCFZE9XloroN8iQm+3jXu5HR1VTj9M9vJNc5uw0UrGOhmcYTY
8if0OkSjR73+IHsQ5OXDxGLf3TAsV1ty3NDn6QSUKeZ3pvQXW3DbPlkyZus0V2VWBptL7M5YiRiY
EMS1qHZE2hsxG14oXXgNTI13yaNeCevZYjtaEzU6W93Q5QmNx7ne4UTyTzWoWJUn6rb0WuNYRH20
wC/ZsBheeYn2II9VSVCZkAUCT7lDFE4US0OlM68eRZ6BjNFHybCXAS/+5pGEWoVT46Cz5+0V+SWG
yol5XQhrSXJD7B8c80h07Rtny8C0Z7SbbvXsbA1qZeNOvRIbNaYcd46yepyWm2Ag3vzcqm1dDExG
aFaaaaA9BI3e2BKuztHClRPws/qiWpL+raM8EEVXkqrMxbFS26Jwvfs3hNK8UE9U5+wTnXzNCUME
P4dQ5kEjhRsGmvwvCRwcZxGNb1k1gx1j6bOeCrEZn/DPOfjz8pOW0Z9KHiVlPjKVm3QsxEVdGBAK
etGdi/Aku8ncaLnalmbxXJg727P1oys7OEz6j/3+ZzFqDbzfB5Yt9VWtEykpttz6gGjqDPWj/hCJ
jRuGiZGTBLTK94TyUqoVGaU4Fv9o8Nf9pknFG/buPIWUg+QEWNFGQ8qdZoGAHuPBRz8d+KMRTfcK
GgPFVBVdmGEd5xA3k+AjczPzNq40vLgW61MDkYD34QKeY0A6z0LcM36Ehg8AcVsz9U2eWdr7jm+k
Cc5AEi/djSydJqKNgESGw30cTnn0MsbmlmzP3ebDzGNWwmHU+9oGxQKNzVR59/2dTp2uMa4gxSGY
RYbs+u2CDS1/Z6XfNtsiQEn0UyJmKLgdyfpYHcmPNd9vZ9a+BitKpEs/2vH2LFMqB1m7bl4sKNFN
F+zAPd3gYDDw/izddkVZ64VNHKi06lV8zl7sgNb1B/lwCwdE0RcDegN0FB7hKk+l4nOlC0XsFYbq
4tcINx8nVryy4vavCSj+/yk+1EyEymFiPIimUB/fHPTIoGaort6SEk6aYNAzSAnYhMgXdN8s39Is
O0XcK8AgTWQoVaV9o/1c6aOqNX456vxxZttm4AasB/dmDZLvzS2/DgAZjv4ujVV0U/zoS/vSfiWp
gw/Fi6u/Rd5D/jBZEBEGyOAs/UR7iHEcJq26wfvFmvIIkZ8e/xK6AI/KpYGX9znUA9fCMVG995Ku
+/kVBR6yk2YUJisAeWuN6/knLvwp/fbKFg7/YJRsyogYAjK5DI4+MjPmEAdoif7EtJOpDjX9tAJj
QU99MhhASczimd9tD9JYlQj9X99jahnADFZRNTDYCXhibw4L/4MERIIU9b2cmAlzePnSC8xCJwI+
k56LPAUJRugO/DNHI/HkQhGcI2uuc0aWzzjKhVhpJ6rFh+ZCVheQPS/wJ1m7txtYuU533Aq9pYRT
8/7mJnt5RkijNbveCocz9fd3+OH9C7DKJMzXGqkHEhAUcq7ZrC/vc2rxRPhsr8XAaZt9GOvdGAeB
R/i/AX+GQ1EZKPYdluBhmd3dcxtOKCq+eG3BVD4MogMu0gMQAUh2UB64yWDWAGoZd0c5dwCTexQi
i6JjlqLr2bDFYiRiLtudzVonHl0mzNZi/2+uIIsTqKJ+zaAj7odxqWtOjWn94CVNMTd9MJJiUmb+
d7rHDBuaTkDsihbgqgQu+bMxmj6WpPcxijotrbAdjeCSSmatqD2Bg5bv1bWvZELUeO4p+uZ06zXt
He1D5873e9OI0xbWlQrudTF3BbAzhF/JJK2jipzjfAsUbWJTvC2jzF+9hamSsV8RC1gh3J+2Dc9H
bpmfH9OenAtpIktzhkQ6TMqpxY9+z+LX9xu3M7UZ1ls2n4a03Q02zf9iAaIgTucaM2zyFxPOyjP8
11+PMohk+oI61IYIgX74u+9PEZXX1QRbUASLszdpJI7iuabvZ9SJUvFmrtFEDBd5517hTUpcXlN2
9WGV72Yt3XfnDZRwpQYQWjYepuI7R1gmZnxR/WllyFBLZncpCGRHndasxvyT2otU3ufKuxYE11uu
ip3L52AuHh3BEErMg/bO9n+9ymDgQfUtcJXIv+6PXxrecpIpZuzypocJSbmbhhxPqp4yJDt9k25q
FLqv8P5cfsiG8msh3w7gP+XKiG9Z1bKUfhWi5M2x/AzKIWMqqNZ/TGQjp+ecWY9X4Dgs9VILdEEI
lWwgOicEa0p3HoIsaPuZ7pCK0nl02K6y2pmZ/Ic15ON/jlDcGr8rMDmvBjnhNW9ME41tCZTCzGCP
H0LW9NLmE9tiY6a7b07BixbXom2GLiDu2Y2XuJVZgw5V3X5lUXTU5eTF2NuxH9l0lvjdhIZ8AOoy
rRfSbsj5KCcX7hnFKbtKcZWkzYQvGUIv+phQLPpi0Qe56IFzAYMrqlyHkd6LC6L7x8xqKAOmQ0KV
jDs69sPDCmOip/d8VoRN7eZbVV/9I7mddvgRid5D09l6/7WAbJZmULcqmp0trtCf+TjJTE0UpvOv
lduAxLBmXAJinYUvOgzzyBFIehQgLZo6XjvV1RS7sQCjDhqKOdEPIWCmT/Ow/M3nyOMuu6gb501X
FbMMJlnMoyfGtV258O06nN7qEqwt/MRA+HWMEtWTxU5BKmKtYZC75iqUV/q8SsL1ZitvD1O4WM43
I66d9FVhYcEHUta/3sxbbDanMBJys5f26BJoU6MyHFP7xyrHRzHeXbGxTHYeI/wj4ZloctF3lcYN
8CthN6O0c0nJsODIV9gG2qGXZFbYjHfXtVSAhTVMar3BLqzRm0eXIG6E7v8D+6zGqHh9ko+zs7cd
Pue9m/QQEi/AnkdH0JbtY2taCdjY6Dij6e51VB6D2rG9FMZBPo3BWWYfQYxpw5UzwDBCzAMelaz0
wg6VuJe4Ye4/UCLyyBjAib5TXjnn0VlrlWXmtlQstz4KfgotXjLIZ9FwfWR/Nql7eJCZOI3Z4cpu
BYKVUQmFViXlFCyRVpRchZZNXx515UM7YvbA5YiYRul0/qSftANv0IgnsFUguyI3T8+Vng/JdiAC
Ag99vmrXWeRUiJrZLlFWIemEFddUqWmgGqrSj7Db/fBY86mlFhODacE8UiSGJTcO8KyLlEEKRzUQ
hcooXzxYz9f5pMlslXzAsGPWr3YDTAoKSTjI/hMFFDIVFVqgO6PvJJ4+kHg5RHJL+bffoKhxOsTk
hPFV51tc/0KmRQHgrOXoBK6ojQNsIUeJyc+eDXlXPfPrSqI/6cRpi8IslEDtElkXD98bAKZGo68W
NFVxHs6wm+lBSPJjsdZS2XkgSps/YkQDI72jQRZ0m0FZEbqM5qCjGU7T4bQjhSExtoMHdn1SeINt
7GUK3E3weRiyEbWP8OBpTICeaJ7lXZu2KP7a5HyAHo7ZJfQaFwTdD5Z9JgJUoIBJfUIgz0z9UU82
tmBtVhs2reb6AxFAB+c+W6rcuhYRgfpC/7scDPEL90xZfOoN/Isi9bJw7r302rGfCbhk0rfcq0er
xFl8F2W16KLJr4fRn48okgxeLSf5/A4+/r197hptvqdeN7uSzMQvTg+mMYTZ5KOzSdNn7wQZM1ze
fFUcuxbcB1SxMIQbLlY0oVUt2W2O1p2GlDuMx4UZe5FvOiaU9MedD/uMbm+s+V0EodEX+x8XdcJb
SM0RBR+SxI/x0m34zs8rQ7vnPEc9f5bdf+MMlCEeO1PuLFFf3F2UfuaJsFQKbRG5CbmrFe+ZhnDA
GmONmvTb8QpaZLeXf8OQxpJn2aHE4VpRl/c0JXI12pracXDDiAZQI9muYHiVXvTb9rMJ3sp36DCf
Sz2Rr7qyzhWXIscsIwTwY/2b+zKSekp/0moNcclVT4ukzy3uML92o73fzQzmPGhOC/7M9hWsm1jT
KpWRodrKSQVSRXalGMKRggIBUfNj5CZ0cmdXRq89WnxAQz08C3pJBxF0gd0z3gxpQuco+CN/uReH
fdiauEubqTEOUHFo1d7ozf9YtnJ9WzFY2C7ZmMHtHdJppL1nRFIrfTJ7tBCWJJFJY2YnTYolur59
mi/az8o02ptKd6WfgXjKOlPbM1DrbLoWD5/n2JMFgbRyzQbZAcuXyYi3uayj/uYkUEcshzJcwWXK
RwcTdh3irLJeNFjlBFVsQSTXG07E5m6X8boillfMx/ynrKgx8Sr90FuI35emxodhrb3E/PX8U0It
/kOSunYfpJFLWVBS5J0zTI0Yd21WcSc8QQP8v+9t4skLm4IAhwszbzFRNUmYHswy1W9QPKU/9Io7
I5YTBeIFQMtfBDUlgpbl7C2LXLNSIzOU+PimkQnG/cLFHsrlRclKB6xkX2MVLtwu8HtI04TzseTK
REx28XfXMdnaA3aQUD2ujjFN/OEMM7jAtt9ugtEyh+tfP7HjQder2qDOlC1zoZ+NNMAF8uQv8hCS
egqvKN4el0aCyEvteB8H5D+8nsMGpl/Pluot4cRbt15g1a3pV5vemcAdNJ4a6cwtfJYRVeWcUn3u
kLrs5EH+jwOowIzQcePMrWNyODxbDPK2l06DSfHQrTVQPBtoZiAr5b+ayzaSu1AQF/ExiGnCAqp8
XDXxBcM9tT1hMxr/tUgZk4ykKA7AOnkzuZF9TMIxAVNk3LqDc4w8bFYovXIvl0pNDujWRGQYOdGW
d7hM7xWZIFhFljIKdiwow2T5FyNlDnooFiZ8lEoPXp1qQ/XEB580dWAgcRW+2+iwTtB00JGQXJIt
2aYiXe2azMvixj5K2ZAJNCYy9T+ygABYD41W7+5j+enMcsFKWkNNRZIzQCfRV2MGjYGeS2IOZ4Lh
zdrqSSSzvRpWXTqqTz+nLZBATc/Ubds3x/4bqgDfRgc4u+TxeNHzLVKPuqhe4U17m6SX1tN2ybHH
/Vnxs2S1uN4DIfSWETfvQcJ+yrtiwCqZgjrN7Ko34+w1Q168XYo15UBt1QzbZRIIa2psgzDYeZhr
OarKWisFiGyuxIOP00Ss0faVJyykvsqauD7PH6WTZqpVGyILJve0+Q0a/e7J3I0PVCTjlSX38Yde
MmX7N/LGjdcA6kAdLEHpncpcDExVwyGO2pwrFy3S/+rxExKDiWFdilZ2buvd+5GGSu4IoRqB/dbq
zBrNyr1Wxkg/6A+K0IWCiZly/7vLP3s1moyfykTzEe0dI66G9ZWMiRjsCMFCGlY//NaqC9W9IYfg
5wmR3039pTzrDTSkhcguRp05sgcFQdy+8LNeYQQG0xVjyF+sImOey5plz4PcVH1Dqj9/+ljdDfdb
r4+vV6eQtBdxZbnwrF7ttc8ANwnMblNSJ4t6emqSnNWwI/15KIu6byes/l9+tGTv2RuLxC7bzmdJ
1t6rKVphQ9FSIPdpdOeHQlz1u+rUSwNVB+fKKhGP03/SDuagH5QE148nzNPd8IPqr+qrnQloceB4
jo/QKY5ukywCArM33eF35e1hKkpWZ2+sO1h51+yP3HKolXioJbVVC2o25PGnQhPX755lae5ZBMru
+Fs6nJg21/UIzf/CfiYsq93qQJwdDOZYP99iMzwVjKC9wrwVP/NL//tNvlumHRmOqA/BPRsbBV69
JPd9PsF2A4m9qN2n5z5g3Uj7501AHxo5lvL0JFy0sJ19Lz/FqEw04Kk9l+BXI0dXDROlQwA6H34A
SOaHDXrEpPqhAe/jZg7yWwWYc4NEZunQglEOYysolnqoMTlze39OM50iKjtNrBKoicZFOcsryXQR
Py5kWnk8C66LWW4l+MX6Dz8GeRhq4/MNDPKzKB/ugHFumeAhHSXSeBw0j9kf0iAfGEvfa3CtSGue
gCC7UFpfG9fcZijAP9XRGAaI9iIkvHFfioQdmn0BUK00QYRvdgAR+DhO7vwTS0f0nWzzJMVa8jCb
zL5Q8Iwozoky13n3xfUQt41LKPDGj1AEcJIIPTSxlokcF3u+fNOPkKNhopwq+56JHtEccDHLEtia
cRZPkVwjHRf/Iw2Nu0Msjmu6tM44LUIX46P7KVCuJXajWcjB57CcdBPXHQjDXPiM98/ef8CAspWR
TJ8UO7pn9TcOC3hbTcTU//iVEE5RDaPh5XT64KgH5eg9njCKmbrZuk1gkN7zbrcX6bcVvrlpe9m8
7Wk7rdqUAidzUrTiSwMKg9Vl7+8nSKV+F55OO9VYlcXC83hK1uxdd68OrrmbYgdVHan4xY3WCR+0
U/lwFyGVBAjOVTDB+gPqSBLkLkmnJzMSAe3i4sHaAnTpXpxpKvcyQnq8F7cCSgwzrnsqOE3GD0Xl
pbkvJZ1VBJItdAWg2AUhnsXaremEuXef7wJyW1lOScj6efHW5Fbl2+3oWgrL8y5Aw5ZdYDsFQgda
1PnI7vFtcILE81b++4wuo2vuIoGrmen5M/4+Qb7izhlUAXmWZ6c+jZkhS/jSDP+bsHXm2Mfb6g7y
gFkLYGrgfwTZc4jsULkL5mFB2RZNo/rjC6N7FcX1des35hihMcSIcH3Mxhvj2CSEfH4/Fbb2/024
t5OmWM8MJUbcZSTPUTpsSBLxzL8waSq8oY+8oU6QpatV9iuuryKvc+qptuACfYmcgvQuchjgu0As
Jhn5eJud6eo7mY0KEmuN5D5rkCiYN8V2f3ZsxeI0plscvVml7gAbQPZ7sPdzJeudFX4VeWXvqMw8
zIu7xwPXTKliYZyLcABehA6Ul9FcIogZX2KLFAEg1uWeyjEkXQ0vhJp4PL99kRBi+Ag4nKQDy5Xk
iQQ7svomWgX407+BHRkXMArZGPvc5pAqlmPfjYI9qzhv56iujVF0AQmIhLeyazioWNJu7foMsqA2
hR/zFHl9qoCvdrF+4Uwt5gQaSfuZoG9o8s7BPOJ3+9MXFnUlk4qWBGvddAjQf8n7flST39FOuLkw
WkwAR88FFuuJiAkpN4DWb1+XDDEA0nvmHfNUKPDHsrrXUOWbS+W6uyFVyXAKdYzgw1HSpC0P7Z5n
djb5fSWTYtS0N9Zc7eg85k7xMLNRvhyktGr0sZzquT+P/FQije8MQ9DnhpkG8TSmb2Toe0uGlIRk
P15FOluwVM24kzGoVYf7fdyzpm3HYcsa4eo30nb1ZPFO8DYgAO0/WqXYZOd2f8gB+QIBtZagIW+j
QnCQrt6yEenUdhwaoXoPpBt+lh76ycJpMycdX/RixAbvffe3aFKY0HOBgTyBU3gJvqSqTn1krIEG
1/Q8yQFQHEcvezwmS79cue3azwcMZ+EazDiyvEBFIl6AOR+4rmA6mnzc2tR372cID8mAsRCnpG0l
WbbBKw42XGTCj85Eg6DqR0mHhHNERZug+ZP2J2RqPyOuv372UXhVfGXb2iov+u10Untsxp/JPCSH
8givEThSi2iG3kxM6bmAxXbMkeN/p4R3GXmMbs99r4N0s6klsq2xYZTrvjtBWsM2h72oJqrVCNLL
G+qUYeO3oBXsayI9JEAE9LEVRi6CuDjFCnLk5YoeynF0AzYdv/7VMHf6OCNJyl3rX039UaPri85e
ssDD0wF3M3EQcbVNcfF77bQevp9UaI6VBbSfYAbi8FCSYPR7HzM3h5lq/Z/ZSZI3JZhiF7ww1FZT
E/W4GpldfxUyprC4dzmcRFO3HuHKlSes2fjcwI8xcEdWrQtWei62Pdc2GlSG/zELK/hzHTKzjbuS
wlq6ZQmTcf9N5qi9PjQx0spmshheWIX/zlkYpgKC4hppN8TBRYJAF3UiVUl9ByaEUWwqev9YSxod
vf39fHODDFE4y7cnrOUlwrRfH4a6L7SZlhT7MRpgQowblgw6H999TwTptLagdY8CIiUI3URyrWn3
JBejjFEBiw5zVycn7Dr8s4YdxU50mI+lNPj1g7j2vjB+ziD7uQJFvBTxVC6S2P70LYj2lW8zB4Q6
77cytHOfXBy85VJuzDjNQWNlVjCuR0hCtbEnm8HIK1AygNa8v8E7lVSoz8/kk+QVKQ58/NVo5Ztv
pxhfZSSa2z3lyHT2YgDdXlQI8km0lR9v1GTWO58cowLR17CFKuc4VCbW6Y2Wn2Cxn3B4tlvxLqOS
7bmVyOSfCr08LoRTQ9n3trhS3YhQxnrmnLzxcnFHB49uyxK73ULhs00AsPnNfthcz2BKkwOo5R+N
KRkI2Sov6XndIsg6GM2XfW/4ysrNhbv1ic2ykZSyi8JjOf61N8dipOXq0tq0qdXpNGsdaN+csioi
MopDnuxXQzsCyL3RRQ3KSU2f70x5qrKUt3P4rPoxjIOOSMIbkrgOBN978Ly0Uh6TnnFjGVt/Na/r
EpOipsQPWtWrVQVD3tvdLZ/3omAFE9xzdL+gttG6f1GbCtryW9fbsdv7OmX/H0qsa3OsJlfGtyTs
RXPU8mog7JMZSFKE3uP989WqEbVQpiBuVAoIWn0qWBDWE1eg3paZKFZLYPZ7gb717wtniDY4uVji
uXskOIl9rEhDJgFn3BBgBwfvX18iC+miWtdbKcfrGHHl57s23dhfpM0a76D/9E1SXxfzY1YsVSmv
ld6+ankyueU7HOhGUg6OvTHoGtyMWKIl1ZP+9+0A1/2btYrzRPHvzPP86a1v+NnaGHlv1KXNGr+y
9oFmdXawnzjo66dzVRAWN8SdTmqboGPAI1MbA2LhJLEGRNBaNEuQ6zZAV0DYx0IY0ZOeqzga47AZ
69/sSK3SFH30keSM+abQgsGPbxRG1ZSnlEaLYaqaoVq/oxj4JldHTIOiwhavF6feF1aDIUSSu5X6
ugFc1MsjPb31jxMrgIaEqjJ8BvMUx9eDB1VxNLQgnT8EmMrMQQ94IwY0VRj5SZzWaAGqv90B5yFk
BXKr7qR6vmJFBY0orwoF8FaUEMWWImSAz0D67ZToYu6ruY3HxiYZdc7ZXXEJBFgAk4yFKapSz46W
cGTEvWlt2QfXJ3jXSmgQ2TMC4AqnqEsuap2qZZAn+ReyPA6URdaBcWK6JUHk4PxGJ6KMyOaWYSh0
K6mMniVQAJbSdYoJIH9GTKTRBX5ibeIBYZ8EObhv8EhOewDKhtt2/QNGgxBKxzPCZeEUqBKBuiBR
Hl6wuZ36Deo2m/WAXlUgzf5JDqNVBkZD2Vx05DcwJ599xb97Fo978grEdM2L1JdB8kCLGni7kYv7
Nx5QyVUX2Ry6Pr6DVE9r0mCTpyzVy88YbjWpR2b5q8oU6unQ98wDympkt0vyZBlI/dNBUnVKn6lU
V8EPS7CQh+J5pbv0qTFavhMSGfE5/h7PToCD0qQbC6uBPml6QORiH/yZznQldEcLmyDKJ7lM8TUi
BQKS0WYwL5CdnnVIWfWV7gB5MgrMj2JdWelJngESXO8z31Eo6ZZBNwQ70nrk+EmfaB0LoSxPeYC6
Oy1qcw7Xu71xr8Wn+7qst+2fnMaaOlWJmCKxNbqD7ybhxc/tVtNY5MjkKGlJIV6LtIiTzrgEJIoj
piQr9+6ACa28QMLcIxow97Rs9tRP07mT3r5/BPV+fY/LSxN6GDRLEVEo87AXO1yT0Srlj9xcSuJ3
o5mqIP/O3YmMdYrHHyYep0pw8RqIEhT3z+REI5vFmuAw6rXNEdH9Px6XT05b8oXHvSRwvouZZ4Un
wSDGcB7rbAO+F7VZdFkXb3bWMaov3d5Jm/uzyhwAG4nVH4FmgV32M7cCNm+YebyoP8Uml2bAtxdH
yPeP3gjKq5w86dIKe01rbNrCQQune41VxfgkdVmjKAWiqDs3ryUTXRGZuCG8Tj5v5qwz8uhz8m1M
W12WzivsFvfEnDfyiS0JyBbbvG1iEZJMwU9VOMagE9iOi7qa1m7K016H35Q0+wgJNoCBs68iRXSH
S2OhCLO+hi2U8XGp8BhL38Fi4Eb72vxtwK2MaIGUcN26rG+70AYwcESArIlWSG1HrsFap8LexUk3
CK17xmfYN4RGy8fr3ZsT4rE92xgUgflsRHVyerSDiNDyT16OYB0N+0LTT8c6iWm9Af2nOUBopCrM
W75GrytB9ZZ8NHW9LX8G/wGr/gwwfCRyWkuagAQzWxeoHHELj6cnwoqDvQsppouWRKYRQsUoFjQJ
H64V5Wh98f4188hbzxywKLOnragJkukaE/UXzQVr3Yv3udU5IEKoTpFHz0myyY8xJ5NTTbAagrOK
1a+7jUrS7XIIETI+MmNwKazkwKZym/Z7COt0kGY/9FHA8JciRzzzfO2oCt+lY80s/Jhka5Ia6+0y
LZxKh21VimlKg7Hzh2KVuopaPlfb96081jqOs+ExLAgVyl3G5V85Azxz7Yd0Bo+ZUXE1fCeZNt+7
L789+78eXt9fvUL81BRWiwsVMion8Hx9wdf6Ou6ALgBh2YkvRV4SPpsTv/RzyGDuYuPP2RjSUpoQ
cSYt4b0puztG/ntma+0pxF24saPF+JJamjuzV8FxDledYzOE+HKxJz0GhweveRy4F/htgdp91Y3/
KteuT9OKhVq4LJpC+vD96Wrw9x7pIQhDaPLolTNCutP+HJp69t100/n1Px4K9YW8y4JS8IFK2Q4n
9HB3+sfYW+yTTuy+PKHri970u6o3kvAtAJBVK+mNy5QLJczOckxlOETpVhd+rIQRplARoXxOdzQF
Meav3VkBLUVrCjPmdSoOFQPuZ7N0AAVk5uXzn7TxwS9XYngSh0Mz0uT8c1rMSkAQMO4JX/4Hbf7g
NSIashFQPtg4tvGiJk5rGedBU3lIYk0at/2GrsY6IjbZrcGD82gdjarYtmTGo5X3uOiBWla0B44g
zeXs7n65CUzUhuJSyRKdCzK4DnhBjeQGE4yzBG1FmIqCSpuCRoH38oNRgA4KZOFj47N4U5MUbQqS
d8aav7h5Ros34/9wYF+dL9HHZxLvidJoArvI9qv08rr8FCHhf385bOgPigVxPAclNpxyENXXazlE
3JF62J8qdyxRU8GxkotQBYbByCC0qvinlS4XpbfmO6swUmY/BidY4Ll4umyYdnZ5vpK31ERWT+6Z
8UHcH79v6g21Wp21swOGd3TQ5Bpa36Bczeahj+u0vJyiy35Y3R8+3X3cWZxKVMJ4CHnFdjj+6rip
5+XYtFW4LA5FTgZwSZzhlB4h2lQnLspBWHfpAbuEZW/0WHCnV7y/kJYn1i35OULqx6wuR2cWaKWn
9US8+lg7clBpKZh48QgBywKInAM9CK6TqJkUwVqwN0LqqDiuJJkdOnNbpVe5mpJDft5AnSd6CW3y
6yaAeinvsL/WZ6YUPf6vxakPH0FNx4v9sYAnK3xx/skyesxgqnSzmV5qGh6hSwTik4PfI6zZfAxU
cdgEoDQnfSJl1cqdLsJj031ZgE01OvAR7pSguTwaFUFMQJR1nv59ue/RtJsxRsXGVVxUqnWxvHx8
crbrOmmvkia6oQlZnv5uunerp+hr047OQXBKDTssYJmPOGIXWQJdeSbiRE1syhtnecKWwiXPH6r/
C1dWqgBzp8OTLdRP2QwuCKG7rmlWLUehNybAh0XuXriBFwv63M6881wks+FhWnMzEDyLYRKlo6gC
7iOGNo3oZRzQg5B2Xhj1pTdxdEqVtxMjSUGsv4V72sEBtyfGIWKW3ucZslaWmR6a2NPpqda+i690
zwcuDL5F3ibM18KFVVrgE7DOAwcYgHjikizVi3t/Cu1TnP0iIR5xeCEroamSvZF/y0T61fNG7EwW
h+3P607kZyV/LFUcWOxT9n0otdZe/bO5RHi8Fvo8BwZG3zjxPW072wGnJGWfqwAljdlsQi0+3qlU
D7WQbEeGKHVB4A4AaeBE19qsMA7gLY1HOcxYc9/zxit09udW69NArJdCcEavA496bTlBZZum2APl
VcJKe6klcu51T3+kALkCkRmgymH1o+t9WwLY5vZfBVLTPrcvd+5ghqGaSTloXBANNlUBy49OhHOf
Ug2PrWlb8gbz81UNamQFs48p2ZMWX5rUi5b41k+jC3wCvbRYPvGEzmYF9JW8hwmzQt2G7IqcmGHO
mTszWztXZDM19xipKh+AzOFOXuyd/pP10VTkEHp1AUg5ej1ZwiSrvpfgj/I5oFM1A47P/k/K6DvG
NWS47lrSKps35iEugPYIvDxG7Dl4/l92XRiPEUsD2Gx+LO/98XC0g0SENpKRlgp2mttaRCvsrkea
njBYWFDJHaYKrbG4Oisr5o8FVoT87Dq1KDhMPaLcssshrekDTSJ1xz0n1naiRsVjP3jfJbTo+9KY
37d0582K8fTAZHeA2MfdOlItcNDkhY29Ks1mmBNnBAIxmAK9sEct5ik0clQXpt5DNAqpp3KHGObb
83riUqqANq8XJowj7VbrRGiWLuljdciYG8E/acDcrU09RH14avNkvzZC49D8UEhugZzRANw+hguG
8xdPQaYJUdksX4sWaXdezb0x4vgDRT5PFiVvY/3JiiGqJRpajPxD9O0agPkwbqTTX7KJK5srlpND
orJmDYt7nQMkkZ/XZal77S898jlDskZ1ozEBzx1/JUi4aRLrbC4Kh2bsyPBG0XTqCFi/jyBn0Ili
9702JMcFz/mtJTXFHACTihN+g4NbR1N9ZLldBFVHnj6kXwADsL3XwrW9OvXsYPQKXl4y/XpEtqP1
5aEyzJYbKiOMPRJCcCRCay6A4gU7l+yY5vjlyHHTv+qenKOx93HOlaqRo5U8PvWSBkXOLpaLpdld
cbJ3cUQUEmy9zGbj5bDMaFATkPrHD0FaO90PhgOawLpMHdlOYLDo4hasjZYuhPSneWBPooBjvNKC
kqIVtVW0xvG3msg1nYS3hCnYqlg43umoA6kak6jinZ6g1L4p2JG+rtasEDbBRXGZicAjzsKOBbQX
I3glDX9GjKrMTGs+Ryj1O2jWNlesQxf1Ye6VZ9MuvKAYFQbplHuiZJtvVeS98fG+CbPBhZbSRJdi
V5pcUIGEuVr2LjmPetd6ZAZ4voAehQTR7Dzbd287QJUpGSraeKzrgoYxhlSmZGDQ3rB9izIyADvL
tP9kGw5mHq9gSb5dq9UC8G59Bh4QIpZeBY0Qx0EmJrRPuhiilQ4I6T9AXsNRuH/ygKPRCT33DtFP
caBG/59fOijTcfawqSH1OVxXUDlpAgBlElm/MzQkJe1iJKUCxmfx3HFxwc50sU6icQWqjb5p0rM3
37xXi1G3JnAidVU41/zFHMEHl1MuNBOLaJpVWJO4dMaCtrBU48qPzFBtnhhfqMSYJ2CfsqWOPYn6
P0xv7AACW2Bg2i9l+oCoFog5aoIOHcPRSGJ/M/H/GkJsEaGr3GeMZimu52YMHO45s854qu5ijZ8s
lKkgjc2qafzhq4Fg6JH+22TKaCB1/VBwmN82Vueue40Rh43sdBbTXYFl4RG4/62XBX091jZ7TZKs
cmUaSwWYHJp/a2KDLza6AXoSksIMahMM0tjk4J6ltIeJyIOmKIwIgEUf9HoHBKPEYQxJMGMB8LXv
mSaHE/JAiOTFXOFnLptEBAFGfVB1bDLQAgRzoGJbPzkdyom+a/g9Q/igkUzVqLR+VbvY4xhCagHS
Ut9TU5f3Z9ae1UcN/07eoej3s8Cw6FSriycGUwYYr7cBKAU/74nNRJc4Oju1gJ0fAbD66SENJwJ/
tNrueiV+XFPuUuv+i7P/nEZrhLUhJOOS8LKAPB8bKRQKeBE+0sVCewEK/EmennKtQnaOn3zsJa29
4BNUzcWzOLL689x0H/ss7fUipQqfw8lYTNp+isJBmzD5LFWtKj0/hmlF7bULSXiVtj+8lKUUJGUm
XT9tqqGUqrJfzR206l0Dz2r+2R5pg6iu1MSQDcqkmdP7O35eaMktRmgNmetJuituVfw6G3FB5Izr
pusEjuzqiEV2I6TmukxLsiELrbzDgzt8vHSNuzYhaQgDNp03bTzTpU83lflm/MDJzWmXYP7sq12E
2hxByq0enD9BSwvLCUbj/KQeCLxTWfft28gARdygDrtoQTKoPqRlXilb8kvO6NEVmbcH7QcB1NLj
o07942gdFDwd1lhVFrcPARy3mdAkPOqkjhfaJR2Ry8MQC7XsFfEJ1q5341Wv0maci5kJRV4ILy89
UTmwo5zusUlHV78HgfXH0XxMUXtaat6kgaVzdAUVKUJ8sTp2nACeyEJahHKbdpO/jfSu1M+hppHk
wpMzInrg+rOWO3xtTItxM4yeE6vLyJyBRTMKXerMlFf61/rWQsO4mzrkxUVCuCPT4CGhiNpqV7Uu
b4dM91qzh7q/7uX6y/bzpmVFtQ1jijivx0SiE1Pxq5AfbRJRplReOMUoHH/Q9K/6CNTU4Ya0w4iv
7wbdf1m32Yp0l0KZqYsslMLyKsAIEH/amNw1NbqDidXCjJh2WYWa1aqHsNd32RU/D3a6psWbfoX5
9a3U2URUtfut39gNTEHdKyHhTbwo+Oa/Sef3GfuSUSk+BuUOuplQU7/x03CbTU00Jgq1vJsFUGnH
ihuKGfaz1ab9Qqym5XUolfybtrcWcaAamBNF+0+yCk7m+NNJKLALTthLng1oEJtDpv2A4v398xqc
uzXV8v+5IcJeTHy6IfpVYHpJQeUk4UpZv2Ljqw0KMFleahcrTh0BQtT3Yw+Wkye1Qwo6dEua6BOf
O3IEf5v6/+PSBZXqLw7OjDaBe0kXlPQBujc9utWMKt/PutkkfN7UgPfR5lHW5IFmFV0hENTPn8wU
6FRiXY6asruF1gU8J6ANhY5kMqwW5hkEULbGl4jE9oW+4VaMkOYdObBspJvsRQLKGOhlLl8HMhcH
hrua9uE1irCXk3ve4I30jjeY/9ZajCIN7M5d29pLoXJhkaWMrt1YWEodnOh6WgOqdDAQ3dfkCy9b
Jr12aoNXjza/mCF7OwQC5WJx+oNLkVChplHxEmBV8RArtTXQ0vVhKtKeHbruUNktndozpqFets7O
6cpAZmNmvHXKK5EgmN7D2jQx+xy5v2qkmNZ2YfVfX/TiRHv9jmQzRLqeQuTQCFgq37kqwQhSMlfa
hPZzmHfRhE0UhmpV1PH8EnRcDYwIMjXW/KanhWlGe725zGVXLc5wvVHcnEA+7wSO4fWKDbCzexnd
4AS1O5qk7uercihVAJ4XbBvx+7uleazypZ8Evyqsx1IilTqgtHf4OONpdP/ILHLkCeIBCMQa/4DT
Y2LeD+wRRIMh+7/V11tA3vIwwWhrBj4w8Mj10OXGoDAXmxM/SoJteWWI+tqhnrjN5oCoRJgZ9zeY
cGADFzzc8GR0FwbAWl0YjZ11JT6ko8A2JBxhE63bcOAnCRDO/BYyVuWByqOHGoGAHZCgSzWUJF2U
3lBsqMDZc39KfgpwhfCb8/kemWHLaRaZwHwO6yQ8e2Xji1AXemPbTzAoJenjMDEzp1gWlxz5aGke
Wr0JolkMfBEopuASHbZ4Z+i//BQoD4KWKJmHtgLj02bYuTL/0H9N4FXIcwz4sNsX7bCrWgRVWvki
/DjM4vWVAlFgOg9ZMSnrGfwq3jU8CR2gvSsFxWMgiOgt3fN2UC/0toLalqC0OOKk/iRivAXQLdZZ
K5voMuoZveYrrf+gDptVnANWFTiWvr5aIFiG2nH0zlvhsT8lX+dLnT9Ymr9zmgImLDSuPJPSXEzp
ff5FIxDB18sjjQQE5rwsEG1o6oud3fmUBik3WQpgAzFL97qr8khXrj6SAwALybbvRrV0HJ8IO67R
ebEP0Go4l/kqgfHoKYzm57e3Jg/zf0FEQUKoIYB/WYBRbmCERZNEyr7gixDcMAOwKBbxh2omFM0a
MIz/ZNZVswtKTBIsJXjeLpkvi8kl2Oxi5C6wAOQ3Io+gDvkOB4obWkRzIHDJ6mEZjYCQg23B37/f
HR19+o2hWaIhXZN6IDg1WpJGksiP8SX/O3YPHbKG7U07QIdrolHnGeCAMoXf+BlPdrAZDnjMzwv5
l0Pp8on+sLlJa3/JnHg+dLqCIBN9Wuxm5eztgjYYSg1wJwZ3W6oxCuSPQLul8rk9rz2u2IiJhzyL
g6A+bXP/kbPtAXvgFpNI1zEI3sdvvojmVAT7z2w6sR9Mbrcejo+rzpU5Cxkwk4GqibLmf/UW06CM
44n90ZMISqAK9ByehcaB10UowD+YFgSd75lSnBK4BQ06sCi1wr1uS2hzM+h0jWmuJGOZ8EIC5L18
8+5ctXtCaEvpx88eAhGeeIoxBNghsWYReUbXUhSv857RKLR5IFhNiKt7PmHcGaojVtw9wUcmjl+j
CXWs9UX6KEr1RJXmFlammLT+icTsUTPqiCTPD5uYnR2EyyaSIz/1WwZsJC4rFb+qpLWDovMa0hAC
YvtQ7gD3nrsw/NxBbRF+kx4Bhp0dL0P6seJsPwHSM2AG4I8ySa/YqMe6YrCn47hCJWX6vjNSpyBm
LOjIxO3oDFBMMy+oint0Q98RKue/x4UyNOi/RfB1+Y+ket7LO6c8GYxnBKn5mmcT5h2penKkylEa
sr+kWAMOKbUkvJhJ1Q7HV0vqcYPYAukrXNAp5mJXXztXaLLcVL+fd0w+v+ZOidC3tJD/i/iPuQCQ
JjGx+xMopCrdUtS/zwC1u51ni+y/y0aoU+yASVV31tkp6iWTTYwKEDVLmkhbN+QeIQFdDemE/+6w
jrRphfvOrV4rgBmGC6V2uekrx7/mgPR0rqMDOvuf7RSKaY+4tUoPZaXr3qcs6szPOqXtiYlKvuS0
fPLSE9ElrlOtVJe6J+4N5vkYamrMnQt3cbefy2ptgW534IkD4WPQisdCp8z5J+2+SHs25tU6LcYt
bq6OAu2frxxX+6/5TV05KwZfMDg2iU+Cp472QmDmyJvhYnMql3Z5rwCWvNfx3raadwCgC6ZYWjnI
ZiHxI8708a2Bc8/9NfNqPjvjFblF3Xo8y1VEizw1bTgcVGDueXftGvfYnwxHyW6nbEWj+X6oqND1
PPDweKKQQusON6NDQsSa/nHmkzXEQUihomkL5yr6B/BFkwLvVYcOrrAXBXrj67TLBDzrT8cbYARo
1VXsH1ANXKUcfSPrdwFKovk/b852jKKslYPTwEvjdiYTxmPlEFbnhG/SVy9esCFIUXiwr7W8UhqO
3c3c5+hHG3axyN6YAX+ylfaiUTy3RRjYyPQvPbb44eI2JBA9lAn5l80gtjPN1Yd4uZfOEr1g2Rre
D8QshG3xzU9DdKwYZZKs6abr/Stm/VBVuGH8SUWg2DraZPOvU7EtKwO5XUgbyVUpRViu5Dtr6EDg
CvzwISWQ4TsSJ7LqfJ5pVolzfEzwI3qvx4qxDRhZBqxKBLwrDUDZ7uBsk44ES5pFGtL+oF289fGh
ISfEpW36RwBvNRN0xyBHD27otHn00soRKaCCOWbP8Lt0TcXJ0IZu2XIgpXWX4O0HfT1Wvd0t4I/0
bdUHENYtFGEHNNrHqUozqMwDGWG8xOBQZYb90Ra55KqUvJufHXiZvfEpGCjhp0ncHl08TPHgw6sW
PrGzExU34gSWc5ibJHJqrWFV1JXqS2lBNprAYvZov4QdvojFJFfwGXngBil96XORQr9VKNWFyuGa
SF++/YRy0aWH5gM9pGH7SlfzCfjh37Gp8V4QTmvMEd5j2X+pBCJZ7IUIBCKaQViEpnnEDMoYfvtF
A1V5b6ILChEnLlLEqkkm+6zEj2acdI4/ztacL2ZfAW5ceC90KvVLEfQc/fvliXjFE7z/a+/ee0Zj
uXARwMs7/ZJUPmeVFp/jjs1vZEf739MMDf0xh5SdyWINlcxu+v5NbyqeZLAIO2WiXYxsXdJ5uIYZ
zKm82LHMHIMkX2t169k3kXZj7aRGoT4xZkEXypvzrgXDE/hS1eoWzpewmdtXu/u/b7FYCHBvO16n
h+R7i2P2eXXA5HdgYCXgStZg52q/AjWRaT75Ji00ZAg8GIbxW+QvbRSnTWDbCz44lE8pBrxelE8c
A+5Tx9SU2Dff4hN/XKvlH3NJVTYdym+xWmWlk932uzSqKTNz8N+BE7RY74Oce7kOb4b/R6kzUocg
nQ21EFfzCWy/LQVOWCaZoQhI6pzgxJckLCv2Wd8vWVM23RNpg5JoW44CgIoEmSvD+Q2vb7Q3CBDJ
08n86N3TEj2fLZyKHKiUV0r7mSI4qaWETFifrz4yRTFYvzcndC+U0KPFvrnTFGF9UW4UE0v2GeFk
rBPGGd/Qzu+qSC6LyMw0Jr4i69XbgV4o36HUz29Z2+gAy9mxsreSDWCs83d6XX6uXn3fxvDUK3CM
P6Kzci2kqyOdn22f3DXr47YNSmzxzKHo7qddJ9mxCKX0//FTq/AhiHR9hpdt08gc7U8dHKnoBGd+
YQZw4FygwAdgAZn/Krt5oe4ylTVIRnM0sApDNvg8+qm0Wnc6yHw7cXAiP4d1jvX8EaOMec6MFm78
xALm3NX8+1OjbCrXwTT2OzB30L6/gxdlSopVw8G3E01ZPaeDLOUcpUB1tfNhzLZkJkao0xLnzu8t
iWLPkseeS1xVqf1azosFf+SkGdXvXo3xTTbpsCYPP6oWToWmY7BwrlsK+Op3WlTPN+lcrqzm551k
3b+LpVZuGC26ouR+vECILW52XGWe9k+51r/tpXA11bw94/gbCNVt797xAk9txMhvH/UIh8DVkj9I
2sA2AvXi1zCEn+cOJD+m7/WhPWu6URw4oFCnKL0U5YYPLM3dLVpjcy3u7dTTi4ayYP8NgZZuG2gq
vDZnc1n2/LnTTITLSYQ3U/wpbmZmRKgKUWiaBEHj08/zl5WesaRzJRhBnLYmoKgo4AUPFrxn9Ski
A/gl5cnpcxlxggzfToxT8BYfEcep0DZyiggYvLog7hsCpCMHy0y5nQTuLlazc/PwPY7rhE/ZcOvz
G+0PL+IOrDfFkHqRcrPiO32UzpQLHm9iCBoY4UcKqz36xWB8UYXMouaY2kjVFMz4lWla91z70BD2
/eTpxgF7tFyPC89COCvBrQUb0J/pl0wsRYryPy5132HgN574KLbcTHNzVjKOxuNd5BRwstPuBQQu
9KNElXsy3Dft4CzhCTEAVAtrPJIBlKRzAKQDzA48e643GCKHWVsiLb3meDxJ2UCQve7eMeQ/4lmT
rrsnnweFzkH4mUpySdNIXQEdMjvepFRbvmLYBwjP+BnuNC+R4BUMlcfSorfjzpdyVn+rqa8AT375
Pd1xQwzchlzavM4aiKX6i3hxqLIpXfZ4+SxB//IUn7ZfU9psjlneN1ibFRx8ibyEKRXOKfguENut
TlQ5hSHYMwvfTyNDWyHw0DeIDulGQxBWlk8TW/B/4ZZxqhELfH1CqfOwmLOAnWodAj6a9817R+W3
6zcYRwxGHq66AKucoG+t2XhLHcqs885VxZXTbwwJ7JouSUIvnUUVE+9hMaPcyntn1ZwSI0dcTI3l
f9P5oNchI8lI4Jl/NiXIWGL8GKxXY2Od1yfi3FEQnJzrhBXSoHe2d2oowzlq2m/abZORZkw6rklP
wa9mEw42n7KOVEDPndK9ya5AKDiZw1XHvUXScJXYG3h3KKig3BplfkcCS4kplmbEPcUNscR49Lkp
V0fZgzErlgIPJrE5x/4rIiGsnEkfJ0eipvJqrOcR5vAk/GHcTtrDjzAqDRKfwuRtFG5lgpujdwcg
FbHTcQY5HE79TN3qbUn+DQc6qNdKDPZ0Zk8fNVxZM0H+7Durk6FT6beBdrxChWrPXshmpjuNIiGR
GvVJrcGTtpQCw13s3/ShpJCUsdC+VD0Zo58toBlxe+P9dI/onmuBQzxrLtZWMiq3WoG5syQUndVb
hXOYU7lPWPXe/dxnc4kDtf6CjgKbdL6GdW1kB8wjsVEEs3JzfyY0B4qtBqDiZXQwBgmxU8vjqYfT
eO1wIPSWILiFS77QBvCMEB84Yx6q4+3egFDdzeeV5cAI/Dw63IOv0fLLO155Dmia82VfuqBhl8Nb
kyY4NF84uybasiRVjFx1X/rEzuUbWCp9b7JJ7rAmSxvdZaIMmyoeA1XTShKU41JSME9KSNyqgZjd
OJ5xt5bms76Pye2cSOnbv/1RoGJjSSwGSqAaVpBDNextBC+d8TxdwOTAP0GUdnld3zjQ6aWQjM9L
tuGRIYZiXDWBIwd6nfSjEBqTbFes/Z5Ya4qGwGfwbDHyiOLcsRGo+VrU29gvjaPdZASrJlm/3jMB
EMJW2QA2tRaWtiOjmPxAhzo9gPFK0HmWyufQ3xt1BuDqt+ZxjdTip49EvdmCQBhKiZUjj9V7ZSU7
Va64TDsE5bmPAuOdiu1CPOJB2wT4Yizal+xmi5weNIuJVKVT1hJGo9vNSjNPwnPvkwyXx4wAMnY/
W31SrnocbVWIpnWz6q0fpp3dnrX54SJh1u9ia2DnU2+qQ8zDRzGb3H4mhkiHdbhWEHB3N3FNNQmM
T1OhZKiT8nJyZpj5lw4dVwV0CeWRdc/QjGpCgUwvMa2yqnvih0JvZSckLdLe1GwzsycBggRtSbRk
0+hpGXeJTLaq2Yfi+JA/kCCubuCeHllDXV/b35XhmX/90Pt42/r+FZORrFp7vcT/UDwDPotkMwcj
9TTAd2MNovAQikJihy6gWzNJsLOE6y3RgBhJyP/cx/Rl2VEQLCcp9xBoj0KB2HxCvI6rkUbSnuBr
K+A2Rb98XSZ0dy0E9WxCS1aip/evfGOdz5gmlfBqLjUJKgYOMuDck8pI1CGTXg9Ml53FKCotaeyw
Td9VGwQMY0XAHLEsuzzVuHk6HgIUSGHjvKWDmjXJnoK6/oPvMiCCctu2N8InG6nqGTRzZP5MnmfI
ZmV0zzcOknvvQJeoLBzar9fE6b7OteriTRQ1Tclifkn1e5AxHnxRi7WN2vJGzeBH7bzOEBVEis75
CYVsRdFI+8a3lHEcyH3/zFFGGDyZjhaX+XADf/nqQ7HtdsC74WC1YjffPjf9Y3ds4FummfNL3BwO
D3uO8S7mnX1pLVjBlMHJrhs7azM6DVbnLRNszZR8ETgGz4niIRc/r1qALWd3G8XtO1vp7pHAdItR
RmFe4Q2iNibSs+SUEMx+p7bZOdSw7q0P1moVaSgHcLkzRSutnxXN/o/J8JxB2gbeygz92gGOU3iO
Onn0a34c9UmwcKJXVNKzQeiBRiTfwmBeN+FwnDzG9DHQfFVhW5tkJWZsNt/wGmHzIW1w6u/0xOGc
p7JFTG00ip0AEsZjE/YoRy43uAkbJ63Umj/gp6xzUZo6RL3mvfIeYzlXUfQm0Tr5A6vmjizVhgug
ZJRARIpvzGUrv6QtpXp/7eqQkZoRuilFmGHqqL+GKBmGtFDxsoITIIZmOIVcpvGJT/BFmtNLH5Lf
Oixpcnh58mhC6RA651+zoMIdxc46FBQZ/W1bYsQwZpvy2QMJebIQQImqDab18by357gvL2jovi9v
OEpp64XYEXwcYe0ad4i2Nkm3ysQNUGURgK7km9EuNPK0UDn8cH+BgHy67DE9pSFdTzcOrMRsx89S
BX8B3pTBb3DYRjIh3zSchS//VRj7818ZPTVkO80oJnlGJGNNx1147Aohx8cf+8VBI4kxaGPvya9d
SylLBjpAxOSDvTcaG25VOffP3RlkdsaI1pmkUQ84EiNYXZYehag/H6FpN9p7FvNk30qpuiXRasIA
FSwegyNFyaT3nvrHfw2opzIrdLO0nSZp+sDowu3utbdOTsi7LuDjme8rW7iYt2KtP3ZBvB9MeFfG
NW3iyAVWSQe7Ow/7XPAE7OdNXI50IqPNxtCbSGUITcd6ELEkUP7EpE/zCB9XT4tUn8FyJeFo8sTP
YZT+h161grvfsM2bsWtOcfbmKgG6aQRen5hl0/wdt2SA1wv9NdzD2TKDBwOPqv3/vMAcAHi6d2lG
w3VJZMg+9baC0DqjX6ii/DbWy7+YdLQFe9VdYZ4hqwLjPUk9jA+OlBqpv3MeE/LmXtR350lrpuCY
T2OmYVd2WnKpwvaXqsCehRukHHdAiD9nGYOZmgSMVZkzcm2FLbMWf5oZi/YvPeNLAUtPgr7u23xy
bw3cLtm+HZAfYRxupGT9xqhGw4aSTPjnlc271maNNpOmUKwgpUs/1R56xi3jZdhfZURIWyNb/3PF
x4vG2kcA0GpFFwl6eDH1As3uBPrsFNNixK0lEPPsHib1Xj4dOBrt9/hAnc3cksoP/zqFHaLyl2lT
8foS5OJG9mHsrXW9y1nI7GX1+baTEnGKjvfapAaPIoSiwS3GyMgQqeMdG2SXrJMmoCqlVzoP2G+t
i4SO3qZpFm3NXSo4GmJEow5GTMA/f004biJydfRTENTCIOAZ9NQVyWUyBFBvUvbmnLxRdquot0yV
+ptjl87TCAelkBdSGxN1NP9fOgYN9NjJtKEg6wRTjbMCwPcgem9WCrTtqbt2oZhe8dHZVe3gk37i
TXz1H3FdBZ88fd79dEg6TG5VN8L+vey5j5eWZyv813v/f3jeB8ZNK60jVVVYSy/7M5CeOWPAva9R
SS47pRkhrzMfGnAAjwN7XS8FCwDctMrNGZY7RsOH4DUiRLW/qha2h38Mx6u/8Q3ZZ3gkFqvn52NX
n1vdsMYhGQfVNeh6DZ0cG9lLDhRm1FZluKxkCko7sN+TFYRLELhAbYpysqCfIZ5yrGEuaxTSU0Ls
UsMW2Ep5/PQ8iynsiFbr4GOSv78d96pil6TcNaXOrf9TWtNKBt2X7wiZngyP7a9pc3LxG/QqASsR
4UfppjT/2S3kT6ibjle/42z0XWbxI6SwCsMeJyKCPu2kXdPYnP9HYuXmcUj0bOSgb6QzM5FIHYm4
Q2st2fgke2iIA/QGHHAhlP9J4aC/6F1biP0iH/VG2ZAxN9E5EjMgEDyF2vQeF47Hlb1MeocbBtfC
X19sapuRHLC6CmTzhBWemOKV/27PW7/AItJGQyVoL/ubpvSLUOHS9S98GAp8JQwblf1V3lYYMcuF
uaHcypD94Vclii2Df4QQi9Y2JvCKjFLF1XXerBZBRXvwDa2n8XDF/+Gek34ZbjytE/PBqGk9d687
A8EwFIvWZ0WSS2rguMVlmLgkVCt7hwmITkFBCSHTQdXpK6EJLaAIzF8PQWF/CUlLC5cjiNoLPSNj
NP4Qxq+4h7XBSn6feR/gsm3QuEmrgy7smXJ+bX6ZCk+fxw9kE2ew2yQ9yvE3iPYtcyNn/eKntoE7
mGzdIVj0G3A0nSQ+daJIkU3ixRdqWN/qlbZqGKiwUG/m5B0MOAHPh2nllU7UoQnXVtCveKwrtGSV
O/tvhEWnn7qzlcXu+5RLHYGAqUlPK+Tlhs/G+s3ip6mdUP5wzzDxbx6Um6Q12RkcdbFFPjHbiXWU
eMmX5vXqxPVFJTzbHDnCoR3QrS8jIG4CDH2W85Kh46BVV//RdZ3D/Xpk2QShI4A38J/fgcRPQvq4
kVKhvScsL8H2KbD5GHMnx4657NWee2sqYKtA1vzh6P9YhLh9YJHyHhH5AhI1Z8NGqso66llK9ddv
bPuQgXS5Q8tNiLGl5/sgvzuIwUQHND6BOUarj7CPm+MP3mESKbpuAMFPq6FoovrO3jFhCYIftUFv
gcpTvWeWbw0l66k2FQHwQDV6Y9n1KVlqAavAAoFsUtPqkMX8IvMIHlhCfiOX2NGfBUzDl1xsD5P8
gZMUw69zVlkYNti+60frM+D7qHAlORzqKIaV6gRaw0LXsf/OpXz7guGRyHmBiMqOblTWXekrosCv
mNsGfNYaus4CC30i+E8ICjEwWTVFwBHyhbh+lEvVfVZWimI7RE/ngtldj9hfm1ok6tZvCBUUs7TF
LggGnxNjt+ETWlcr9Qtd7YJUO3n3iybKQ2ryghqSi8NbiQGvMLDDphkV2Qd4vK4NVr+OjMiDvR4F
bQnYRK1GXSEyAwLafwCjDsTo3ydZQeYl6+k2L5iCFh+DEf0rQK67mybdFW9GLaJ14t2CjpclHR1b
Qk9FCP3tBiiyn8vKo+vzjbLQeMaW1VfyduXYioQ0b9I9y3ZFSIECDHHCX7+Mfbgm1ZXkSia56oQ+
Tkhr+7zQWEUvlRz8DoGtO+loYGTPoTSVfugLHqEBkQ3EIWi3HQuPj4Z98RVqWN4N33wL1NKtHK1C
/QbkC3k3pEeYiMq2rpe7ExmOARwDSMDIm4teqMBZhjAIDGvcSC4unHGTl3jzUeT3h35o2pTh+mDn
GcaFMMY4+YzjL2vY5Gx01U3ad0nTgtjX4kV2Q0ldsR3Y/82Huy82Idyf0sDw3HFiWNlcL+Kjkchj
RD+2hj+51+SbffJoTzXnAsvFvX1JikiZ5fw4Xv2VfH491Mb6I2cZFF41lTflzvISse8CEOxnARLJ
CI+XPbOSWTZmqeIYYdXXmbvPPrfPswWxbPd6LtHEn9XsIh3qge3WOHmbzfim1vwL9pa1Rkey5uJ7
kOS7Z44jpZsHxlpqdHcGtLrFG7dhRiXBGHOUki3U6yd3aqjmH7jWvdgwH785NdtHdoKLxS05tgoc
1Zr1ORuKmtfbDuo0n6OoAc6G4TcaJsPas3fsx1ec/hKU35GuGTYWxRmama9MuBpE3uaV51EzPdAx
gevXcId8dFsF8Lj31CQXdqL6pgkDSqaarWTKrlGwrKBZqViDncuopaqJLmiroj4pnbudRz6wSeYx
L9mOm2HsTjz/QpRPwi3+aNYwu0lsmU6EwJduGIep/dJAkbVByC2/kolP74Ja3SAytepTp4Kwu7cr
jVXp4WUyOhW8uPggszmAyJB8DknMHAOGLSRDXoDhToCJBJhIFherobr9sT1ss6JTVLbcc5awziPN
LopylYQSSKCuyPs9MevH00zhfe1o/10hgJC/zsCI7wchBmUgvmgy3gxs/gOSeBGXq1+H2t/iA97F
o333vAE28Graz89yV/NcbcJQrNQ4m87QYjy2EkW5ZrtmzV03r/X3Qfxy23xweQoiBZ0VAHLClAPH
8Z40eHwjhj5S4nbjSMcqinNLaiL3cZlgine9/j7T1G3wRqDrvd47HSqzZ/aJbd2fWeJOF2zeuk3G
dwgLhfJCLaB5y/Zm1HoMhXgPg8AcF1oK31Il4KZmDF8k8ufwD4ON9Lj2KveR0z/C6WEE+Ab/3iub
1mjIhOGR/9Jdgdh97QPePi79dlHFdWRy6HvVZ8TPUTOuJOMK7HVl/AV5HtkCbBPRxW/nnNsnGuvn
SrxSEz1gC0kIQ0yZXnRH4lzzNhAXeWih4M0gpFDALC7X+DVqWh8XruLFeBdyZXOhOnIumecQLYAS
PSfEWp+mHV3BmkrM8quLBo7X+T3RO8/cQQwjuZ04lxgYeBuLNyNsxbpLroSewmyxhnV8XQ/auJnx
VxjZ+rk+LmJdgokSMDXGOGaESiYpQ8N9YsR2kepPEvRD41sCerNSYQFSPnh28v+PNLPS4v5xrNou
N/Wb6925zkwa08TfuRd6FPYLeeWxlOLd+p//q1mYGx1vLuxaumc5RRXnwRLAB4UoTtS9F0EBDr57
6DtoazqukIxdKyyCFjni0BKHcGZ50pvd/QXJPwqGPsIQ8BTkHkZz9XD3LhEin9H8MrFidyMCvwaX
9FEoSTIC2U9Mt0lhGOVxhIKHX5oPI6p1tGV47VgUPR82sxV0aFzZ1c46wvvDbT1C/tzukmUU2kbK
6jEN4beEoSEX3lLEhzKFv34/vgHcmApb6qYxqSkhao7iCYYD6ipjaq46ceTJNaOVNpkdn3ktUabT
JcUmhUVgexbUULuUeTSDBWVAJ36AIQNagFjze8YpbXgtBLxT6ma3yF6xx5oiQkwjyMHJ3q+c0pEJ
gbYgP2p+L/YlX6FsT5FXPEkjOMeXK1Fyei5CtCeUAw/K+57gmAU1YHO+okFKVICLN7IXUNdk8n16
B83+YUBIF+58VGBvxRRed+CCf5PzPEmesniropH/TfQmaso4YC1A3clCdH+0hvtO4uZe2SMjL1mx
Q1/zfRJ7nA6sfwfqu5VOXNHq7A2wWrIU6lbxiQqKOteO3WNfl5q5HjGtIgYjZgb6pcNj7WKXbvHT
eigAb4G3PLGcDuBw6o89PAWaV4ZCU164oGD0Go2Zw2UM6QVS4G6RjpWxPx+e5P5GsJhZvjhoNhI/
bkrVYtrLza2QipX0YJHEMh9urd0+VNxQDzHwqGX9/caoMGAi0+MSvom9EiF+wG5glSevjg0zq83s
7F/btYIDVx6UbC0qeXfW6CtRcTGF3k7gyobx3tFh/UAbhwTKxZ8OjzW299U1s2mt48epcz1EOqXj
yhH2avghPKpN7PtEh1KYTsmDgdpBl/AJreucs8nM5JRIi6Ptqi5iL+eGBRASmUuaVaX1xCkX0Vge
yCVkPBAR+V1YKR50u+cOq1C9zUJvmfDvUKni9D/NwgCjcQ0HiQnThGFmXnns0IvoSpnLdtyxOE03
lfzqD6CmDrdAT+4B8ygjDxFQrzvNParTjfeyB5K6V81eeGzz8J2fGDitKt62OeOVZYedstIXKbtI
0oAc/Z4Iq195ihNubBvKhJKvvvlcbApJ0MS/K50kNW18kfzeYgPr8fNkzEHOpqW717z9s0BJ/fzd
jZ197cV48RI/PoPJYJqXHkyh4E1UBwvQ6i82vDjHVie1MGCW5cdPEc7T0ff8DF+jxWdaYw5H2gCz
i6FDFez5P6A2Ik/csxPA45+HaF84oivAkkkGM1aTn8HWG7sOOvU5PnegsSl7qErr9KlGkUKS3J9w
Lxkhoi07ecDZo1XuNM7fw9PDeing4YV66VjrBuI//j0HSBGvfqNg7q2HFtBbcIhbHjQQRJ71vTBw
JX974jfYArIRmsknnxfc7pqf/DkbySGhNIj4VKCQCRmiBx1854Y49JkBponeIgVXyG5qP4LY5qtE
fcC2rht2qtAE30hTsPoAyqy4YGWYjo/8Y4KZWS2xqt758ffsOG/m+wRDhbAlBkTK1sOocZBBv9Lb
HmVl+o32P3q7gOBcF42p02VtUO9PKL3GWhLIyLvjDLWiX5EYmk7WyVMP266nKOHyXQ4odykw0Oi9
/rjnUC0MMF8HYulZ29C1Do69PgWlOSKoP1lW5O6eSyLUa9tY//bpkWrjWUROOQ07SO5wZwy9iyfb
39xV1pDuNpXzuc2oZPz9l2Y320HucljcipH8sSo7KPbstKAXr5NXHconuPNdW2eLbegY0FehhcY8
6edPLMI7q7ycx6k/g1k3el2eFLuXuhboP9KmmgDJqCuiLKQrsOpoHiccW/j+D71zg+loB4DV7tPW
VUkWVm+S1189cya5A4S6WvadL/iTIfFp41yRDyfkJpmyLKxp/ZYDND2fr39xGvWJpqawS4Wh7Zn5
Gf6Q79KQ4Am3CRvR1mgAKgXZgHPLkcy58+s+mcf+EJ/oibI0X6DHzWqfNiPjOj2cDaDox/aAVahj
GMjdiR5K/WOG1jJOsq9X3DCNnHZ2QsexDOfpdZ4E3IijkJY9Z6Olqb9G0FxccIXjBQMKvmXCea7I
js7/WDRYUopI46cooLspUg2os/3Dj+FdyX54sMGAmGgrBs8ldrMmdNHaJAmxChQEzC0DxwRZnkAu
nqUf8iLjXmJIB/4aLzQzHqZXiaw4VTfLSnOcfw3+VyNqkIHWp7ytmBvAhuxL2d0cPzPcJ4jQazwA
ZwmUpQ3REUfAbQPbGy5+dNxx94+O+CGAL+2fV/8PImGn8r47Nuzr3V0imGlotRffyqBXfNwjRBqd
tOxbRwB9YA+2yLLWBKneWbHlRsZaJ6qH6sqB0LMngGLNMNGIZkKKZhzDa7COvBgIYL57SD4S9757
1VOPfKqGlgLT3ydc4aW3NzFf1Ncgb64Q1GkEVKW2IgIfM1PsyiB+t7eMYwtPSs8rzJIOjp8zq4MJ
z0zehRmPvHMAW3B51ts+EJsOA7KHe+rOLI8l5fGfn6xH1UA1GgDiPQ4ENlelxA6zPKYTlqEDP85T
ulamcfNkQZ803QtufORj6c4pxlKvcBZXpdde3k7UHfTBrNmvYSBJU11wP9RwDKoAHmnMY8Q1bsWB
UN21W0biGfUGhnSdQLGbZDrhG4ZLRPw4rEtxvXl/Sg0wzp2jGsMoNr4st5ZFHsgw6iRvijXLPDT4
fzoRmDhDT6M2clr6MOGy+g36tRXMuH2aNfJi8zjXjnCVmw2hPzoVUtm7bjY7apmoE6CZS0VXI2x0
nhkYfh6MW7cwNtazMaOZELWfo0iRNBJNot+6vZSPsjcbYXcsKfab1sUhcpeMFzNdBMRPqRLl5oRi
cms3IuXVLJxuCUAmme0PyAyHY9JjamWU73T1z191JHYcTI3fjirnnN8SSThS67zgSEfJvFj/Icm0
PzYL1XdgrRQdeeqrNkadVQgNKlc9fp0Rxr+K1XaP6XIGV8yHHOVfuZ/Dzm735XDBap0whirjCu42
kaDL5lsyrPpqj9PK/qf6y2pT+fMj7XJEO2YHEMFXdiWxfTKWRvT0tjAJ7XU7zxoY+a2yKZzRkzEL
hIAscWEqzmKcZjckdLmQFghrzmAZmc95DbIzg9ii1/7YwDnv89asRedGRej2JXM3Jyewzme0FfEH
dL86smdsk8BQJgjDB7qE2E1sHQo8MMHRkfxUTzOBDU5Ap/cuoPFSs6NLXptpTnUeDdjft3Y/YEym
op0GGbVRwNrI+wLoqb4WDXmO6fHAmZralDPf7kq4dcbN3rOPghdSN9ofSgRYKrwzigeIMeaeckBa
34GQOKyZVb7BF5TBMJCPO0PSSLJhbkT2ZFiGzQ0Q9uPfkypisjkWRUHLygRzatXBA2dTWZpMYZ9T
9teiKFO2d0W8EffGmWrblNvn6ipraAJpXCzV2N1z4BXCpzAhTX+PqBdZLtBFlzuuBV1SJ2Xx6teo
miC3TDHIgFvrNy/szJvDdgV39eVFaz81oihuio8HAN1j6DjJXgF50J6Tj0bgNzQgW53saQF3IV+K
M0LEOVkQj+dCncPEN3U2ftggXJbMHymy4ASPjsuNAudQCneD6h0paMb6USPFs1Dy26J9ODVRA7A4
n1bf8OBMjGNcTsz76aEyHLKicpWjzm/Ad1+mgVuVwYrNctVx3wSW/5zcjIfYIjVDYgyrXUkwT7kw
ohyhbVB+aKMlCmiDLrErFTDywSOas91+mtLfVWKqyw7EtvJ38AHlPQGqF3sJgpS2BMWyFbCZkaO0
h3daXELKmY5tFh96hske4vpNnigu/hKEtvvGYQGt04PH2Ps/LxZS2/WLpETvxDHt12Tjtn6PJMAK
M/d0FsNVZMvbRepL5kOHjG+EArxROSWkMEjN68WVDVLFLSwW7Lt5ZjYOLVlIixPXa8Z+x8poNTsP
yjDwragFkPy9pSEiFocJF6J1b3x0HVxbFJ8dn1Sz5x07UPImJ+DJOFVgWZoXL7JIQSwXoH9p7sVr
ZFVcPYRHNmpk+q/vWhjxPezbENRORA8kiivCBqLbbCuqxkw2Y9qqUsHbp+4joJfHG7iItF0+C6pC
UERx6FpI609YjJ5BegSyxrkBZX0t+VVy79NbQ6s/FQTxaGsJo2of89e3fRfqqHpR0qiUnuYz95G7
+buRZFQoP623PyewsEgHfjTVcWJfaDIYCqCtN5WmKcDh83QWiWBn1TRs/ibZRelySrI66uRhr8Fc
xYN8zEXiEx8P1xpyiwThtDbsTpUn53G0ahrownc8RMYVcsvIavKyeBYRAn8nkWaaFZCOwJ7VItQa
LxvijAHugo0hlOLxP4V2HLjYQl2k2Z41ahjyhEfz6hvKrp/HOXYLYOdWfDbiD/eiSMfoptvcYegK
7Tt3TFrcwjwYhZdUfkdKJGhQF/6JGm4CJF/pvVY/FFA9YcvlBZvJZbyCAI9JlwzM5n4j2Eu8moLa
t8tl5X+46QoVcGLcJGndHCnmMrxQpBdbKhZ9tFlwmmYYKAW7yzBd4vsZe6fTZDOHWOQUzM9+mCt7
5zFdAwBwKeXj+NdokbKxlVR6OzJ7oDyQ5YGBTqOrSmSQ+S2sfoYY+gka4ycWd6GzDzLVw5glFVky
HweBb13KoAWJVPzs6FatGdeFTUhf5+2PBsxQkQYzDdRhMZky13jbUZiNKafRLOvzKx6ONRn4ZhL1
iCw0MRaeIYxiFXFTiYMD6Zpeu6sd5VZaPRvSAjc5YOf/2AXFfhxSp1LI0RLwPZaigoLhvActUyOU
N/OP5fsuF+4Ew2Eid+r7dIm7gGsI2Mj1ZXKly7CPRuwGdDRmpkZDLD+VdAGNAxdxE+qg9pyw4O9F
zNouky/H7SxvlkC22/QADTQMIktSFOIxd//yEMjUevUR4DqpBBP0fhaFYKdL2yHw4gR5wfovz2Ek
rn5fCPo7MIrq1YjJzAWFxeap3iJfSx1prGeRW6QSOexB4iAh+KCd4QyX/xIMQacl5GmTFgAN2kPE
GnhnQov2Rnm5yYBkjKbLi6MlMzQYQM1wvTVSkzadF3KO6xJUFcpCyn06i4R2JqhTSTAD39M+UfBQ
k8iwegtoC4uKXhSnXNJs7llGX45c6qYa9fGyJwDuR51N5G8GpEVpmHE+bluozNII14tihwL24VYW
7Pmc1KtxCM/CRfldfRJ5pAps0+ulgI30HazHp4/so/Gc9Nt5SzBm8V5Rh+8H0o2kcu3DNf9YHrUy
rucRV6QHCfsETpJYOEsFAGJmm2sL7SADB6+EdCP0kt7m9Rnx+lN/B62pcrPv2/T1utarUKFFryvs
Tee1DL+Ae9Y5FzCfZ80qyWtj6yIuckL3RIbqFLFB9RT30JyYuQxInqxdZp2M3UXcAboTeReAPIVH
Ik4Cv4xp64FHqm+ociJ8ioLOZMh/xp44efH+BDXEry+QLTXf8h4SM5hlWT6HDZLMRMFfWsnwHoHk
nsw9zSFTF/YbtGktGT1bDaNz4qYlun2As3NgFZVEJY982wDTic41e+ex7EQSj71fMZfBFUi9EZfY
X6RZg+NX/VtMLBFnkcqnWxqXPDf8yqwA5NBhF3KyvMuSRXmzm/83Ki81Dfcl3JnZrLGeHxMSWIJS
HR7f61g/pB8UEuq76BZPGB2cRd1fH6gpSzPeSSWOPAcuXOOi3eUjTYCDiHvrU1J68cebj2zG9V+Z
2Qz+OZ8oyFpcOnMxTjG3LweT6IIz6W5IJvRvzWA+f9aOAoQwNity3k0Jskf3JGO/r9+ZgJwH2mcT
C/FKv1yUgkH6YWPu74wPdTjvDV89f2TRBS5s3ZsIgosmlTf6FGBqVsK90V9mpv/gk8N9ZASuzM21
PPLN6ABvuiJ2TFJaswl3xgv2umnaKUWFwUCcWI+CAV/fTu+7RFlVIY0gEAqihvAscyIquyfXYiCX
NG+h3O/4tjeZaYobcuaNAiDzQtjKN+qS1vVN4dpZl1t2XThJqtyTWqSmeUXs1o+JhdQDovYEQ6ea
eOCF1Vmts+A7tC1hvgnNPDrEuStYLP2WurCQge1AaxHpLYx88TiY9I0ZEDyqSCot3jKK80bpeZ98
HK9sy2L0UYpCnwITNSagDlkzfm47efjuCYDpr47CpSt1b8FQNZGX4UByIeiC8gMWqy/Oxg+dVF/A
AO5xhH+ZYBd5Cf8TnweKMBNpR5S4OkOp2Bevmc0IMT8dnVhyIjjXQSCJtZoG9En52MZIdbKXh6TR
D0aKtvjjq6jPz6cypUSGOoX238ye8rYaUsxtoSk67VHibf7r/h1F7uUOVG9ba408r4w7EQtHq4ij
SbyUh9Cx/P+Wi0chhi47ulpO2DbFdabWfpldAedgBEcVVlqSNU0Rats1riFylC3agg0ueispITKg
Z9R5YWNhVNuzLwzspMihu5ptWQgBkUuPPBK6GF92u55ZSqBUwpf3eJcM/hS6g9Zi1CgSimVeOTtO
3E3VQEHQ0hjWDvr6Mo++PlzbWJ7F309M+JlAWZFrKUj3u0Ge50Zc5uc49AoM/HUUzAlQQmw3jrii
gp8OK892iwXrOcZIJ5WkEjSYu7D+VOvv2g6AXllIq6fymaO9O/ab/DM5ZZ0SN0OhZZwFY1qRhQQk
cq3+Sfl5dVc4ejorj7j6NIHOJ4FtHHliViLZ8dZMnoNMo9qkm/weRC+U19S90OKHs10tuETVK7yf
M9v4ytCg4+vItA4/FmnoAoDpKSlWbkvrmXYvd4X75nNdBhpf1bZ7OIPffz3K9pgGHmv5ewZo0WPa
S4Ct6twAPTvyj6Nm/ldyogIg/Iz7P9MJyughU9S8vNqKU86Vk31a1x1sj9tU4TzuVqYYtb3hICsV
EpbcIBMGwIKv6uP+016XbDypMzk1qUd/mWsAg1xziZsBpW01Nkxrei7aHrK4XOL4AuqyZTE/KcJe
VdbHYBQC/qJy7GRqJAedP+wGD3k+OMcEBdAhhcq7SK3O8EWxw8aDKlTfp5vGzRkeugTAAlxoB3Ne
HkyPPzd+cvwhHZ94CMPP+rGz8gYxsEXhkKgWrnu2t4L8z+S+P2JCvX5nD4VVNn+ZZPyWZdA/bCNc
fe4Fd/FLKfE6nKIbQUvvYoYgPQWXGDZBxVtGAEhE+Ns8UaTnGJZalycZfmHvV2MTHb75OvSywmPL
hGbcd7RQRcSpPKWuvwMdo6lhb9pg1heuMb4t4AGqQ6vYevTD1H4fbNaRUaNon/8b386ZUkviSV5o
QqssalFj7pzxUTrdrI5E8ILf+fqKzOdi+60Z+zaCLC3breXJ/Ye+R/6idGzvCcLEHQRa1BpSR7l8
bMBYdNK3bv2W8xye1WzQAx9WOI0L1P7D1xblCmN6z2/s6gzyW+sbYwPz1D/UA+/GHPH5A32BbIDh
3afFaGV73ebEAma+WtS5GcV7Az2a18NSZebhcCDeuqaSBEpUOljYG+caP4co41ppaAMRDa6HNLo7
iopTe99cJts9LB/tq3sImldBSwqqVekcUdKcnbjvTyBNkUr4aT9Tuo6XoUus3gneVXAdhRxTZkSm
rEOlJMvwUmhITJcdl6OdWoArklb35WgivfOdecm+BOXzGpvJK9ncEiTq56cmweKaDhI7shR0UtNh
See91p566jbKnofKoYmLNlyY3GTuZMY/Z/1VYR/GUCTt83wh2oAi2T4HbZ5NGr0yc4EHjyJYg33m
lCUkr+xN1pmi3ajyG+n/xEo8yX27vm/FaUdsoAExyq+hKvr6rDlEifEphkX24tA/rVVCTdwdSwiE
n36ATs2LHaTD3BSGPBX8QRnFNMmMea0vsnSRLSICKo0Kang1pzxMc+RQ22Zn4GWzHFM3R8ujeENC
VNOM+7VVpMuhDmG3EZ1r95DYQ2H05A97M+BWfNMUMOdzhuJna2LsyyCUXPkNr2N+/b0mgWNr5BGQ
QXS1rk57cUcC2sNaPlDnbZRxeoSC5jnOYOZamv7cswQ2BPRb4fIr6Y8HKJAaIuszQk8GGl/7ntJh
4WVMfYTA5XGthJuZSnu8S4U4viDebJNDkxTEZuU9sIxAzg5bJ3ErNMbciN6TAxSU3Fk0n2VXY6r7
fmL8YL46LA++Uz1s8Nw+3LkNlEAWOLUY+2z8vJIIzfMxMz99QMzTN3mASzRExc0x+NBO/3/GHDBw
RNd83yoJT/xdQHOCBSKS63tKcDAtZbZ6e62u5Vk5Z+Lxs8BmQVFQToxGTphur4v54Ui9YUXWFXXQ
/ZNbjxXUuWu3B0GL4bhHA5gF+oC5uMnOvZ4DhH/0i1DU3actRooQclUyAi3zeefozIZ5U+cvyjLy
iHedYkWLFaARE/pcUIkwc9BbCqJRBHWJtzZYSP0DoVpFo07tS2cAFeGBa8ShIPKBruztTI1p3PP1
Xecu8p+nZlrZSVy9aSjFuUwzO9MeR+TXjak/vnk3luLYJ+xdKunCU1ygV6RNngyisMRe7b/ycOHz
Cn2AGE+k1ZhCwaKhagqxzB/wMmgj6qU8oItPY+R5rk9ivgn7CKOOPsWMD04dY1x4pVZ8+EL5JEj0
A2nG+wNJzvFR7P0VSLC0h6QFCfzvBuTkwq8crJwfR/fC5OwPw4gGK+GHUeRkNKVFAfI7cXTIdwjH
x2xgOa7bXRlNwr17AATYfPa7iItSDVxVHwzGcer4nWaxlVa+j7VLU3RedjW2wg4qCV2QD6AFXoiu
eLjqVhFvuW4VjSQaC/i/P+3Dr+9NfmsoJByBi2BCyD4mxDHxjHXoXLGFgdtFBSFpkdpA0mhCMWwt
yHP1h7vVlIQeTWGYJ07mb+lF5nbC4uEcO8srDJZINkqW9wqNpsQLnoaP2d2IP3QbMwTEvH7pNy8t
kHpB4PQBOmoTDfWcvRSxQqGVSFIv/W4+rbgCNWAOB2RvWSnO15a2oiz+2diYo6+0hBYr3ZkaDCmw
+DB1FDxaUtIwc8CUwgaQTcQkRohrhzdUdlroDAyHg5V9gNsrv6SCeliZgCF2gBCG8y/0rYMq6q5b
re+WYJI6Hd8/bF2So60/2ut1By27TUwSxykZ4MMwwMkTNr3rP5bYh5apWzTu9m+pkGbErXvy6xLx
ol75ajgv8b654iO97zUSkhBhuPEnH4yMXrOJrT13VBrZizkMIFbKcltwIAwrCvjV4YTDcViO+UHi
BRoHtx8tt90dRlLk+xt3bAGK2bQAVoTunlVzj1fCsLsmU5B2thlEAprqhg3a3aJgVa7RzUeGVyJ5
88nTv1oSKGj1GcHwlFKo201jwxLVsM+JWX/gT3EcNhiQA9YcdzzUYL4256DEM0O3gtdZwI8pNBw5
xExlHK8nujkRl1/0exvu9pYp0AO7deJscZG4+ynoM7ocCRL5OCAyekS0VPPpZumAdbec1EUyFeJE
ddD9V8WLdwOMW071EyIxRwENB4TdnE0olhN1ZhBZyuopaBg5OZDXS+8dZGNxaGtcNCvuECu4hmFJ
K0ldyELFf/rweciKvBN9Q6KJjZfUD8h+wHgX1i+zKJjshMoqcynbRpx5itutxhREpcjX2QcO1V59
YbV8dRCFeLeZOLOTMh6jKH3qCusdT1Czxf+XjG9OZI6ru7qcVsyI8ZeJ7oXF9VhybfgTe27nUy4n
xKEPbzRMtx7tQX8Z8u+yg5kwJlEsg9FrTC5NDV0k13BQpjyXr4Ygf7hWfm5WcCfYWOj5dG9091I7
kZ2j3GhjlQkT8N3Qk8+IOfZFzq/3nfO1RwFmCwDH6wbUoZMCeOTQu6v7DVl89XqczUkxk1pAtNhK
dZEU8U1aNn9RTB267hJFwr6uh/RpcBO5zDMmTpcoA45XBmdzs/y+uTYWBp0V0j1NTOD40wDaOVzs
UcXGPNnjfFjJBiWwahCxIyNMac8VNhW7GkZ/WfLT1yicvUgY23w5Tx5jF8tDoxHZWhkGOSx+Y2vp
229rZmg/XB+PC5JptZodjsFotiHj1aUlKDs23/e5j8bdLgvuLiLg6jlecMlXN1yKszqnsIJUKjwT
bx5FEVaThSc/8J96t1v4irYgukOKOCwFIZaURekJGD33/CcsSmQNh1Dg0Xyo7Oz79BX2fMgEmhxT
zNDH5aToKFc4xX5JiRaraiCqL4+qrMEBS0HhzoG55k/MBL9LSCYEY3J7VriVApvJ417GgIc01bHV
kXCtO0AztJePODTvkmkdB6zTpEKmGxCHyayjuEnnUTABEr2KwPPdj3ZxGyp7YqQPD18UAcoI/Ot5
6gSnyicVGSaTzUVwJO2eOmWpPKdSZ64Aa1cppqqq4k7fqW8j9492U62lGedUqDIF1J64LO5xvRNg
YHoK4O6jeTFNKn15zEdhXDktKt7Is9SVumco5EQECDvYt/i+8Wqk9TfyRbqoT8Llc8NzFM0fpqkK
799+uvgmrPp2scK5ZkVA7+u4VmoCyrZYFiiVvWZwnlIL+kHQ0qr1mLlTEBKoR6V7vA8d8H3pPr1r
rVuyQvOEA6KfgmZX/+I97HPYTRy//hB7TqLkK6BMBEQ0mIjCOkVIo42WHywbyKQGn7Wb481Sq8Jx
Ul4AOAjZa0b6XOfkhv1UxvyjIAm7Wutr+T6ntYxGUaD5U006g5DllyywGNc8GNDrXqYitAZZ7hkk
uEEcKWoXflnghaakV2UEhfjO6BbsvD5ZAQf/3ZJRYZ+PkKwf3k88t7eTTH0v2D+Z7J+JV9Ky/jYQ
N2XEgxug3fMXvlJNOyUErsTnyYl9NyYDoWfPqTQyX3R9UxxJelxtXVvHHFz32MRe+Un8XO4fjRJK
L4dWt7tv+kIjj1eCpQ/bJiVO1F3HQZ3OHPs4UVcp4vmdQviEvgcq9Fi6Ic98v6/rQd7ouxAqzra4
bQFvbLSso2f/KwMZt+SMTItV/8MjzWRblpsneJI61KEraqz+M1YQSlT8Fn9KGErdUrPonCrDTC8o
1RljebLgcRe3Kfuhp6pvkbZtnNpmr5XuFZMC/6mvhPUryONNyRsZ9dF31532Ma/zJtVfVMIwH17F
FljsUAV94Mhbv36mLwB7q6jScnjbOhuqUwbVq6FgWk3L5S41QmcRWwn71aTaw/mmUXT496jTpXyM
6mXy3s/XaG08RhbrRLuAcucFDI7sdr/ER/M6lgZ07zPEE0Yu+1DKyyPbHlK81UMyN6LtB3O2tTO9
L70S7hw2fZm0Rsnl0zSjRitwf8SS2vNo8hf7UDItGSapvHICRg/SnCyeX2xeqmOvoalGVOWPtSF2
k7SWIT84IxmEY73d40E4oTW5if+1oFrz9cbEBGMlCK28nieYcaiQxKcJAXHz57PsaGZnRBKDjvq7
eGRkbpLn6HJmOLoGFOgEie49vm7QObDv99W0IvSRZ3hx/Bigv6lAJMiVVmIxv/ip5mjXrTL0oZ9w
9D/iaC6EladN/qIZ91yt2w2oJnPHMtFqQTlrKrnhTQL68BapAF2Mkr3cpJRPkeuI4oakZeq2rHCo
Q/neI6IKBDlI2Le6/Lx1ZdV9aDqYBZnnMUgLMkjSiQBfrWzpq+CAOU3hR9IjcAphoiuyQBB7JDmS
5uV2XZgXUpZ4az37EaTiMFsxxQNsWFfaQKYQw5qlDWk/P/zf3G1uKsI8eL6icuH7M5G4V2KTjUkv
+tsGsHpNfonfjWv2VBb0raaZzdX4Jc2jJBlYj5C20p1DUSuIdAnkHW0XTxnzharaTR9MCIMpS4pb
0kng921piMJtQ/k9145fxjOW/J/EqeFJfSjZEbor4RTcbnCudV01a+MLqjoCHs5tFmtKDO0MeOXs
txaqlMw3OQVTzQ08yU60vuI1SXRlCs03TBavP+AIlQfLMKgqcUuU/3qmm2aii8IIf0j3RGDQQqAT
E0BlKPzruQP0R1Qm2IrEEX4TlfhRcWBpvjfwK4VoaTuiOGG2wt+5HcXjB8nZ5oeZ9Di1VFaEpfMF
OJo2g69KLy2My5Jtvu/rspB6/UAzMJFYv3F4irqCIupZ1Ev2A4FW2NGOcoMOPwOBXFCz6yoEh4fW
Gr+RdOC6tHqsIy9MnLBomp2RVABzZUU+eeukvKb0NM0+ygy6cLULhJgqkp3R798fj6fRnsPyQqjm
KmUNScgL7X+TKSxpXc+AjqkI3217JjoGAk+hTU/MlHMQR98dLchcKsCK4RTzbYJLqo9nYEYpydDM
ln9apHSmBZaEx+fc89xhWRWcpb6i6QbeUd2TBXuWjUGnXmHlGSQoDA/ql+ZfZ1y00z+4Ml2yNe7J
KyxHvaq5qsfqlk2jPUN9s8jmH6aGNfWYWBGlF245zZ+HaPH3f5qqYuPfB9QOKkY2mDbRNnlQhPRr
GKFHkC6rr+khhOf2ue1uBfi5NVBMdgRN83dRPjBb0TDeyH6IqiqcuaYjid2hrlCIFvZXx63VZNbK
/HjpyIlV5hSvWK4faphlSdLbjy3VeXslTRH5UpBwYTMskudxHzbaSAWmO5y+6eGIlMTu3UCGHTt8
AwrI4cMqL3uTkypuFX9+DixckS8SAaPOmnEi9FC60x+7EuyVWTiKGeU9PLekVEdV0ikDCV4V1Nmx
9QvB1Ax/5V5I0CzO3OijgSbJKx4LicrxtI2uBkgCwNb96VAFovxu1kUjGR17vuGU+MKOXGuoTLvJ
ijdRxFtH/cniQtk8Sux4cKzNO5PA5gmqGSsNWxrwGfihxDA9KJs4qWARM636/3xR6dxA1sggWoTH
qFA2LdkNHViaiBnVV38ZX46vpNdm0ttuK1ja9sE2O+Hej+yZmbfAgQ/c2WVtfSfIT3p+LGeCuQ3a
B7/5XbUF8eFAydP43de6gr8GBSOi+fUQrOMd+elbXXkm+t/shZXsdYzBOc6/40ZDAwCWO4Mf2+gH
MTnszkFBVmqMcMZWs5IvUBfVBtDcyGoQ3gWLZ4KFUSB4LRHQ8xmegmqdObD1y1++YJndRUBliahd
tAqt4jSiL7E3ObD3gO44AyozhcoPKCwupihoATc3qsNMvSkjNKb2NVoskCw7sDMn0lqN9R7nG4K9
hp383UKw6hlle692J2NSqlf04AoPmoXjizq2YJCg3p1z6SGoVbK2IxAaXg1KgWnCtUpHRqVvhXX6
EdMK0qsuUU1rIP1CtnqwLsEwwh106c8ZUeQZjpIapyoOF11lmEQ1dY5pD5O359ZQ8uFwU5I9aRWJ
Lak27/IYkyZeEw5xc/FQxdvZifTifnEZ1gQQYbr5DS6b6WgMkEELzOMONnvZXJsA6ZQ92hPwXdwv
ykLsz7JWx/xISP9XK6w3fRIe3Y0fdGwZqInVPzkE1uf3CJD/2V5x1D9tSOjku3oXIe3QhFnu+mq7
0oIf51f8YOZJmxdLvwju/7+5rEECfcfcWJwhk8GgSZXiKNa7lK81CHUnyd45Bw7FVIEJnXp15alY
grS32UH6pFQnuZ7cCtiJh6mI3KPLF7i0vAhhI+jnrNsplpmW7JuS/vyv8KW2Oiex5wwyWpUOl/Gv
dJWAmnzRtzpQrHOY5ttlaAm6im/VyC+bQvaROtDbrvv6SOcqg0Z4CPEd2g/gWQ6YEAjDWX4j6ZJd
93pRgx6atfGHB26AMRJbmIIELYPhLVsIhSpOT+8KM2xYtlEpcIcYhGchuABf3x+aAw4ppZMoT24m
HwYZ4ZMcfLEVVLp/4jbIz7WBEjiPv7FI3RgqK/5ylUHL3/R5ToRQ+p1L1c1j3D9SCWyyM80sTN3z
DQRMm2ts4komahRrxDbd4gFaxHuSkR6RhdvT0F4UFnTLKDcRojQ7f3IBV3w5pqlULPPECxUb8x0Y
xgieI+gvZtNdTsYWpZF+l23b7L6GOc7kp2zF9T2apJiWdIHa06l4OkuIgTvzRlrpIhx7HFWgbZyO
OS9UrpWSLIKlv6M34W1DpN0JxBeE2ehdY81piKVJoqz5Xx2VrG8lRrEIRLvyjZTP6585sPiQNiAt
ri6qwNcUO+QER+S2LdO2/bN7/jlLHst0yGasvxIrYDknQuKIDeJlkpiAIKautWErXyBHAg4I0FRs
kctEQVcuZTpEcVbpo871bre3ClLNA87I8UZMBfk1bDw+nj+IxqzydfAcuvS+1UO/DcHNU5+v9vGG
97v8I19Six25OqJQvOAhXizYelsVRMsJxvcSCcELJ7mcHVZSYsHnOe967fFTHFIswH+NFpBzMhWa
wHb0MxaZDEWFQ6bgm/aOvOrOq/fx9Zni3gnO8bzyiwG9umzAChtgl6XJnP9yJYuCw6GDWHQti56a
hSMzMxDNTS0Om5ajvovNDVGVzdC+0MVFZ+s1WyzPDH8qHbwa7S1ZlnLlsEDQHlPpI6pCpwAwHwzQ
EZbGRTL8n8YA2cvhSHO8MxZRWUDT1qiQD7iPHe3Qga/YnTg+hf5KoLDOIEIc9P0uPwJ8R4MQTMNH
S2zHX0wuk5TIwFAluGAfKb57xkaliG6vRavbSak7U87+ilWBj1uEWQ6ad4FINgBvh6nrOkLszFJm
hpxkrChZPUbBaajE+Fq8jx1FrBuUb0Q+74pD+UjuZqafTAeqd0v6+F3NLRdFUHIUUV8HFpWe0PWc
bZcud8Uajs8EXp5R0o+0hDz9ne/2rOUxYOiMBAz4QhOgwkFCAqNuVGtqL29CVzElE1d9nfbcqPu8
dPJEzzd0aQNOBQruunWb5M+1t3lJKp52IHqrUlAUbKOeQil0Kud3/gYE5RqfXTBn+bBFc5n2lJoh
nUJ2+I15ox6OcZzr/TcU50cWaU7HZA0l3+uQiQwFyIO3M0RAOKq89myb9zvkpy3u9Ga25ID0i/lN
F4GaNHoElYYQKRlodJhkVUzWbjIacp34aUXF+6OyPOSDBu7NE4zRCczsN8f6K9uE29KX5O0ctIdc
cVfdV9HJrWwmmttHaV+nZj6GGyCDDSCh8XBcaSomLDpHns0SbUrae+xh+naFasZMmM1iooa+u4aq
zbQv+jJZQTKpb1io7y+BCtyei8pnpdqp1TB7+theAVCwxHW4RiVcSB7XMHMld2NuNq3dzzXY0Wbf
Mzwng1X6xnsGEPuDZjS9+bEWcAN1k6zlG9zrAj+QBGkhMYlmMYRk8Z53CndBguHTmTZSxk1t5ZQt
3cNHa+si/dRtOazGk2v5HWb6W/eF96ZgykaGdXMCjTHK2HmS3+q8tA2BFwYCCCrpg7mlKrhHL4zH
jnj9oDjpRkgmyLEJJPENd07isfXknGyAb9jX/Vu7AE4KnIzAcxp1KLmNFQ1BUQl5spbtd8+Twk3I
bqPpyu6WX/xafEdjHxFv3ZKpladZBaYcsuU/4yKSI2yMxwChi2vAG8dwIkgfX/IH0Lor67v1UTUA
k3nZt1lXlUJoHLbGLh4nY0UC/76SX5aEBjxjZ/qNEA3pEXfQoNz04LWqUYQRcHHNG7tMNI8L3tsU
qbAlj94hFGUTa3DFpIbbveiZXLWDpFkw07K3srGn36AujYmM63BgbyC8gWeljs2VA/semKX8cw6m
jIbOymnto77NaSaQ13DEjGlBtkw3/nGj2LJmSKRNv1JVskvr5URksF+8Q8PD/1/1YsbYDq4zaSJU
Uc2kfgBg/k+SnUqPppjSPyv18eF91OtJvlvukXTfm9mHdg9hFa+arLYvA4GppFSbHZOFqre32m8V
/FCQ5Q+XAxseh31aoyK3fKq82T7X9LH9uy3gS8TPXZVIb5zebG75BfedHmWA6Vy7Nj607ufoS0l6
++J4WDdJ04Ned0iAwKHDieaxdPvS2KNbm8pWg+/UZPd3QckUce6emJBbKcWv8bIF9HmG9Pf8blCG
E17tLQODAhJFfotVUpiN/pNkAMMWjH2j+omATqkSVGFC536u6Wa0WKMshgPPgplSGTA1FjBafzWy
H05nYAfz4GSVCADyrexIk/uxJYOC8pb82p3j/rGBnDg63a1eZb8AKLn7OXLXsywSlONRyUTC9QOX
ZlEdr7jg+bCFTRKPjcLX7VG9LohQlxjzd/rS68dmdWKI/No5eVOAjXgTnSW2asLGEeHZh1GyVcb7
6y0oSWsSbp/EN2YfJs2QFaLq5iMU94VWvE7fPndUOusMmx8Bd3gZ09cSbwUYYBpv1/ObKAsto/Bu
5a6g4xn9GGZOY/d4jgTAvwTw4umlVPQ/PgGVa3ovp5GvobBp2Ro7nEVwwZvVT73VZ/83691CZBxj
62cXl0iGx8AkW4e98PVgeY8zEFPJTNN+T/x7OxY6Yv/+vmIFib9SfOyKnbff+K9cYR6oIvOBAy+x
pyML1nC4YnFDN3Buf2Znn7OiPiKeX1yBAXH8fSRdgQeDfH4ikqjpG22/DLPgrgUxHYljzBRvSLqY
z4Zm9IeIlWRkN5YWJX/+WWd6Z6xWbAbmIAPFqD5vL0LkB+VYItiP1g3AnjJvYG2NLA1VRBeKlNju
D7KbzK5QlU8i3KtLeYcT6tnN/wKxLe+ruCTWdqEivElXG1Jioypdi4tFyEMBJ3QxYhOywdCS0xvZ
NtZoS51Y6oQvfYhtI1Px1I4YvQYlAGja/4xJHjYcFTQWZF8mDj2Hrre4Af8V9CRWEWOLVPdfc2N+
VbPJyGGmoWQM5+BLpuW1syDPmYYrrZkmZBt8iBncrnHFUVev8vvZ8vQr7y3Y/cbYSdNSSJh2VWBa
R+L7D9L6jK7pEQ08+MvC8MsiHCxevJacqPUC2bW23WWyqm22nRJlIYaVORWC1SSbwug9NjMqtPxM
Lz1bOtOJG7lbNNPC2PBg4nyEz/0RNDjMbzMiRlvYvGs1yVrQaSRBlOH/yD6kns/zZyf6etFIXm1N
bdFzHn2hvEWJTTrL6M8ohAwDFgoD4+WCuyRfpIyFuq0KkbDQj46JWiFWgykguJa1tWgD68xZIVwr
j8VOjxBVp0LxYCrIXGyOleLrtm6KtaA8FrE118KiPZcdspejiOnBu7kAzZwCY7r545/rqkQ2DEvS
en+YTXZO1UYrWW0j3ZpyulnJWPzMcG0D7L0MAkiLuMHBYESsu58mcqbXe09XWtASL2FZUTxwLPD2
oKrJcUe7S/lHljw+LehrdnuZBgrrUz/1/0WB7gwtHHc/w6Ik5muIMM8XKQ2ocDIZsJF2sQMtkId3
+V0WsBPOmW6IOp2FN83i3S9neL8la43PfnEeLBuJXTRGylQJufpc8OwC421gvE1x8jR46F+v+k5S
9jRTirSJFw4u+EtYACA7KU3TonzrAzdN4xUFO93yErPHHpQ/ffftvsQ7CGB4pa/V1QYl+J0FtD7x
auFM3A/WphAqcbFuoE8lpn62E1gOpmgk1DO6W337REhaDYPqfsrPKIO8IMih1eOxYIsG3gduSoXP
cmdoMgyrLLc3fm1rhxC3grfhE/TUJ+u8E3QH5i8EYZ8HNkyOFiJNb0kL2q0hVPRDYBkJSpEqdIKy
GJ/g9X5nDc/OFy1hbemC5GGG0EqSqIPfEGzURrcncIE93PdNj2xIFkIEbV3kNaV8orYokC1hP9Xu
jiO7/tuEJN4u0S8khVsOupoEpRmzPShl2Cw5/75P4yT518CLc2xLu7voa0F9cDI5dIJZFdftFxiP
91k9af2iMGDlJGDL4ozhwbqCBmvxOsBhZSYHk3FlMzvrO6emeXcEK/TDssDfVihg43cvSFs6uViD
Y1px61Dx6sb7Z732cXENoq5KZPksM1lbgxm7et/ud5kCIshj4Y0PCKWpI3Qh4lYiDdRzkFPLoV9K
QPMPV5M3/yqmdcDv7wk57k62vpZoVhRTqLmeMdoEbefv9nj28PF+J/cHQPLxEIrrwCbEAEW9JuEU
D4pVmS1U6QoqLUGLMCelyAkelwH0Ot0i1lO7J/6T/BglhUE6NPmIOWx9VZZYVhM7ciukKLBBMZNK
WNAPg+V7qaw/NMgiexnPI4otouBd91etb1LYFBGOWhH+gP3idDkmLV0kamlERbWRRZyhJw5wn6dT
+qYbdtnlA3vqBDnufj/BJT+b3UOVdaDPodKjr6FBZvdX630fM15eLHNj4Pyv+Kj6rQGTyaYX4hvA
kqcuOSmDUsDVjlelLqNie8kac/I2ejpEIT+jwHduyhT3EVG9C8og6j+I8WHvpiGKjSmEG7pj7dwZ
bt2++CUTnww9MliKc2YfJPahZGUZOnLD2ukUw//0YM4SxfIRYNLoAaLywRhBQc7S/gRT3cA8P+kw
2vmbn7uVXUpTfFkEjr6SsoncDYYuv++dZ/rMGJHo46X3SGPOxVHQ6BX3LK7igcN63eXbExGT6gGa
2Ci0t+D3hAN8yzCBHSK4irKZTQKuQjS/FkEC0Bn0Mlqu23qUjPNPkzmqbS7ZnSnVmaqbL99VzIzh
EgSZZAnEAm7CtZ9BVrcGB5g1QfeHQc7LFR/dUZCVwnJpPcoPWIAMDqzSGsIi66SVJkCETCNO3FZk
AOkf4r+2B3SBhAZCSMf1FSCHK9MMCYBIOh3NUkVXj2yAJHA6etuk7L1NCFy4lnEZ3IM3xmyyV/1U
0/XMjHa9weelqfTE/X80q51nUwg3h8op2IUAehVF6MfKM36BKh8Cg7xYLHfI1tzyAIuhM+vzFCfD
aR884XqS413/ez1u1YdfM9P2/KYG8CFXHZgFcv+OOnK8y/9m50jUEZqmo8ZEmlLgPCgZiZh4V/j3
WVzo2P7VCnEGACXYBpaK7cNJjoYf70K1ysOS8acUE4rO9mApjxBwiYkwRZUSFmzo1oiEGck0gzlO
+oJQIDruX1TpSnxDGSaBMukboi9TfPkyEA6FA9obDj6vQeMljRImVcYsCL6pR2HGedQE1wJan4CC
BKvYFIi7Z4FIcgIhwewrAVTbR9Y5eok7IHkNEZ1s8/3XYvxy6UrmlG1AqMxEi7qOHkVeZGCWM4OU
3yW2Lf58+cnvKl0/pLLx1Pypyb3gtcgRFuh2lnGRsVXq+8sxF5j+BIbbgB2G5Ph0cJZ214HzVZA7
Ibsb/eARSnT2x5UFqwGwjaDYLBhTQkZs+k/Canwnyvj8y+gcTSFYcytrGWiUP4krZaWke8K9NMBW
bABL8t+zUWWsMz+zzxVryTNWpmnh68TNkDtn4UVQQJm+uJnLj5f4si58VAOconwwhcNWKzaUlxOb
4CEDNlZz3acvhp/3r2/MsJHcfSwsYDa2VuYd66UU+DFaWtpE/c96ait9QSQR475HS0fPZoZ1mQzu
XbYnfuBOPAwfgdi680GijqqFpTp5jxVkJOoBD50TyOhBC83gocHdC9pcPjc0ZrXs1c8pEVpwNO1E
9cXVPgcOfB0K8picF+1Ig9/0hF447I4I0Fo3PmXiVwzG6xVShqQVadsBrDztenJyZ/1vFNmtNRc6
/Tazksy9YTZvLlz0W9B0CUzQ6h71xUIgOkkO2eL3MK/x3TnlrMxlJiO20eT3eQXzlD+yT68Zf4sK
NJsQjq1inDMpvTEu0/nf+v1kIR/PKHGM0uMV2t4bDB2QyYr/WKUULfsMWfLcdPRmFHRS6NFB5fFj
XGjPql4m9NKB+7sen72Y93hm5udTTjrQISNZJCPJhCMYUHXkaK0D4euNEpAkfRu4ClBdEzefda7x
ubKsfngdHxjjPxA/4WXHUCjJKiLdjSHTteFaPv6kJ8WsNWZRxRz7MxmcBFU+EDS/2d6IMD7jVBRr
5MB0OpwwxhiyTQE99BnHoxpec5sgXOMBlmWolZLYiCs6yzLFbjlXe0kMDgmtHqRRGkKsxz+kksUf
oULobOKnF8a3ILWj2hfJyqarkRYuLPhmtyPHrfzOYxt2T8kB6F8J0w7F7+7Ct1aadIh7x+gTNx+J
i5AYoLTyKd9i5xATXcS+ztnjelqz8vIPm39Jo0wTbBBIMlys3ChLRqjOjXw98OlY+PH0QLOXIv1/
ZHze5A==
`pragma protect end_protected
