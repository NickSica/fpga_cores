module tcp();





endmodule tcp;
