    .INIT_00(256'h022ffc2bebb1d000022ffc2b10a0b016022ffc2b6c92f03a022ffc2092b11001),
    .INIT_01(256'h022ffc207a21f000022ffc250000b018022ffc2092b1f000022ffc2b08e0b017),
    .INIT_02(256'h022ffc207a21f000022ffc2084c0b01a022ffc208df1f000022ffc01ccc0b019),
    .INIT_03(256'h022ffc2bdfb1f000022ffc2b10a0b01c022ffc2b6491f000022ffc207b50b01b),
    .INIT_04(256'h022ffc2b10a2006d022ffc2b6c93602a022ffc2092b1f000022ffc2b08e0b01d),
    .INIT_05(256'h022ffc2500032193022ffc2092b1d002022ffc2b08e0b002022ffc2bebb20076),
    .INIT_06(256'h022ffc2084c32193022ffc208df1d003022ffc01cd80b002022ffc207a22007f),
    .INIT_07(256'h022ffc2084c0b032022ffc208df2085e022ffc01ccc20703022ffc207a220088),
    .INIT_08(256'h022ffc2b10a325bc022ffc2b6491d002022ffc207b532544022ffc207a21d001),
    .INIT_09(256'h022ffc2b6c90bd10022ffc2092b2f01e022ffc2b08e01001022ffc2bdfb2200a),
    .INIT_0A(256'h022ffc2092b13e00022ffc2b08e11d01022ffc2bebb0bf12022ffc2b10a0be11),
    .INIT_0B(256'h022ffc208df03f03022ffc01ce42fe11022ffc207a22fd10022ffc2500013f00),
    .INIT_0C(256'h022ffc208df03007022ffc01cd80b00f022ffc207a220bb8022ffc2084c2ff12),
    .INIT_0D(256'h022ffc208df0be0e022ffc01ccc030fc022ffc207a20b03b022ffc2084c2f00f),
    .INIT_0E(256'h022ffc2b6490b001022ffc207b53626c022ffc207a21c0e0022ffc2084c03efc),
    .INIT_0F(256'h022ffc2092b32248022ffc2b08e1d001022ffc2bdfb32244022ffc2b10a1d000),
    .INIT_10(256'h022ffc2b08e32250022ffc2bebb1d003022ffc2b10a3224c022ffc2b6c91d002),
    .INIT_11(256'h022ffc2b22a22253022ffc2b1c92093f022ffc25000207d0022ffc2092b208eb),
    .INIT_12(256'h022ffc2500022253022ffc2092b2093f022ffc2b08e207d7022ffc2b47b208ee),
    .INIT_13(256'h022ffc2b08e22253022ffc2b57b2093f022ffc2b22a207e1022ffc2b489208f1),
    .INIT_14(256'h022ffc2b66a0b016022ffc2b5c92093f022ffc25000207ed022ffc2092b208f4),
    .INIT_15(256'h022ffc250000b018022ffc2092b1f000022ffc2b08e0b017022ffc2b6bb1d000),
    .INIT_16(256'h022ffc2b08e0b01a022ffc2b7bb1f000022ffc2b66a0b019022ffc2b6c91f000),
    .INIT_17(256'h022ffc208580b01c022ffc207a21f000022ffc250000b01b022ffc2092b1f000),
    .INIT_18(256'h022ffc208ba36265022ffc011011f000022ffc010800b01d022ffc207a21f000),
    .INIT_19(256'h022ffc01c0e20661022ffc207a220716022ffc25000206e4022ffc207c42226c),
    .INIT_1A(256'h022ffc207a92200a022ffc207a2206d5022ffc2084c01004022ffc208df20727),
    .INIT_1B(256'h022ffc208df1d002022ffc01c1e0b002022ffc207a220076022ffc250002006d),
    .INIT_1C(256'h022ffc01c0e1d003022ffc207a90b002022ffc207a22007f022ffc2084c32276),
    .INIT_1D(256'h022ffc207a92085e022ffc207a220703022ffc2084c20088022ffc208df32276),
    .INIT_1E(256'h022ffc208df2d010022ffc01c2e01080022ffc207a22b10f022ffc250002b80f),
    .INIT_1F(256'h022ffc01c1e206d5022ffc207a901002022ffc207a22d010022ffc2084c01010),
    .INIT_20(256'h022ffc207a92f032022ffc207a201000022ffc2084c2200a022ffc208df20716),
    .INIT_21(256'h022ffc207a209017022ffc2084c322b5022ffc208df0d004022ffc01c0e0900e),
    .INIT_22(256'h022ffc1d00209019022ffc0b0022f008022ffc2500009018022ffc207a92f007),
    .INIT_23(256'h022ffc1d0040901b022ffc328932f00a022ffc1d0030901a022ffc328912f009),
    .INIT_24(256'h022ffc2086d2b04e022ffc228962f033022ffc2086609016022ffc328952f00b),
    .INIT_25(256'h022ffc2500009002022ffc0b0023629b022ffc208791d00a022ffc228960300f),
    .INIT_26(256'h022ffc2084c1d00e022ffc208df22494022ffc01c0e32493022ffc207a20d002),
    .INIT_27(256'h022ffc01c1a362a8022ffc207a21d00b022ffc2500022493022ffc207a23629e),
    .INIT_28(256'h022ffc01c0e206a3022ffc207a22dc01022ffc2084c03c0f022ffc208df0bc07),
    .INIT_29(256'h022ffc2500022003022ffc207a220661022ffc2084c2063b022ffc208df20663),
    .INIT_2A(256'h022ffc2084c224ba022ffc208df206a9022ffc01c26362ac022ffc207a21d00d),
    .INIT_2B(256'h022ffc2084c224a5022ffc208df20687022ffc01c1a362b0022ffc207a21d00f),
    .INIT_2C(256'h022ffc2084c324c0022ffc208df0d008022ffc01c0e324c0022ffc207a21d00c),
    .INIT_2D(256'h022ffc1900136493022ffc010190d020022ffc250000900d022ffc207a222491),
    .INIT_2E(256'h022ffc2b41909002022ffc2b00a362bf022ffc250001d04f022ffc3e8b709006),
    .INIT_2F(256'h022ffc2b2591d053022ffc2b00a22494022ffc2d10832493022ffc2d0080d002),
    .INIT_30(256'h022ffc2b00a0b202022ffc2500020661022ffc2d108206a5022ffc2d008362cb),
    .INIT_31(256'h022ffc2de0811301022ffc2dd082072e022ffc2dc082071f022ffc2b28901300),
    .INIT_32(256'h022ffc2b2891d052022ffc2b00a22492022ffc25000362c5022ffc2df081c320),
    .INIT_33(256'h022ffc09f0809006022ffc09e08206b8022ffc09d08206a3022ffc09c08362e2),
    .INIT_34(256'h022ffc2dc08206b8022ffc2d00920663022ffc2d10a36491022ffc250001d020),
    .INIT_35(256'h022ffc250002066d022ffc2df0836491022ffc2de081d030022ffc2dd0809006),
    .INIT_36(256'h022ffc09d083a491022ffc09c082062e022ffc2d00909006022ffc2d10a206b8),
    .INIT_37(256'h022ffc01050206b5022ffc250002064c022ffc09f0800100022ffc09e082d001),
    .INIT_38(256'h022ffc2dc08362e6022ffc2d0091d055022ffc2d10a22003022ffc0110220661),
    .INIT_39(256'h022ffc25000362ea022ffc208ca1d044022ffc207c4224ba022ffc25000206a9),
    .INIT_3A(256'h022ffc207a236311022ffc250001d04e022ffc207ca224a5022ffc208c320687),
    .INIT_3B(256'h022ffc208f71d020022ffc2089809006022ffc25000206b8022ffc208f72069b),
    .INIT_3C(256'h022ffc2500020651022ffc208f70120a022ffc2089e20663022ffc2500036491),
    .INIT_3D(256'h022ffc010202fc0a022ffc250002fb09022ffc208f72fa08022ffc208a83a491),
    .INIT_3E(256'h022ffc0be0e20651022ffc0bf0f01201022ffc208ba2fe33022ffc011002fd0b),
    .INIT_3F(256'h022ffc2500014a06022ffc208e814a06022ffc0bc0c14a06022ffc0bd0d3a491),
    .INIT_40(256'h022ffc208ba0bd0a022ffc011010bc09022ffc010800bb08022ffc208eb14a06),
    .INIT_41(256'h022ffc208e820627022ffc208d820627022ffc011000bf33022ffc010000be0b),
    .INIT_42(256'h022ffc208982fb08022ffc208ee2fa07022ffc2500020627022ffc207fb20627),
    .INIT_43(256'h022ffc010042ff33022ffc208ba2fe0b022ffc011012fd0a022ffc010802fc09),
    .INIT_44(256'h022ffc20807206a7022ffc208e83637e022ffc208d81d054022ffc01100224d1),
    .INIT_45(256'h022ffc0108036491022ffc2089e1d020022ffc208f109006022ffc25000206b8),
    .INIT_46(256'h022ffc011003a491022ffc0100820651022ffc208ba0120a022ffc0110120663),
    .INIT_47(256'h022ffc250002fd0b022ffc208182fc0a022ffc208e82fb09022ffc208d82fa08),
    .INIT_48(256'h022ffc011013a491022ffc0108020651022ffc208a801201022ffc208f42fe33),
    .INIT_49(256'h022ffc208d814a06022ffc0110014a06022ffc0100c14a06022ffc208ba3a491),
    .INIT_4A(256'h022ffc0900e0bb08022ffc250000ba07022ffc2082d2fa07022ffc208e814a06),
    .INIT_4B(256'h022ffc0900e0bf33022ffc250000be0b022ffc3692b0bd0a022ffc0d0080bc09),
    .INIT_4C(256'h022ffc0900f20627022ffc2500020627022ffc3292f20627022ffc0d00220627),
    .INIT_4D(256'h022ffc090102fd0a022ffc250002fc09022ffc329332fb08022ffc0d0022fa07),
    .INIT_4E(256'h022ffc090112fb3f022ffc250002fa3e022ffc329372ff33022ffc0d0022fe0b),
    .INIT_4F(256'h022ffc3700132341022ffc250000df08022ffc3293b32360022ffc0d0021df0c),
    .INIT_50(256'h022ffc2f11820620022ffc2f1172fa13022ffc2f1160ba33022ffc0110022491),
    .INIT_51(256'h022ffc2f11c2fc0c022ffc2f11b20620022ffc2f11a20620022ffc2f11920620),
    .INIT_52(256'h022ffc2b00a20aa3022ffc2b6c92ff0f022ffc010a22fe0e022ffc2f11d2fd0d),
    .INIT_53(256'h022ffc2095a0bf12022ffc209550be11022ffc110010bd10022ffc2b00b20661),
    .INIT_54(256'h022ffc370002063b022ffc3694d00cf0022ffc1d0ff2066d022ffc209b420685),
    .INIT_55(256'h022ffc09e082063b022ffc09d0800cd0022ffc09c082063b022ffc2500000ce0),
    .INIT_56(256'h022ffc329702064c022ffc1d0d020642022ffc2500020642022ffc09f080bc3f),
    .INIT_57(256'h022ffc209a322491022ffc001f02063b022ffc329850bc3e022ffc1d0d1206b5),
    .INIT_58(256'h022ffc209a320620022ffc001d02fe13022ffc209a320620022ffc001e020620),
    .INIT_59(256'h022ffc2f1282fd11022ffc011002fc10022ffc209a303e03022ffc001c020620),
    .INIT_5A(256'h022ffc2f1290bf0c022ffc2f12e20661022ffc2f12c20bb8022ffc2f12a2fe12),
    .INIT_5B(256'h022ffc250002063b022ffc2f12f0bc0f022ffc2f12d0bd0e022ffc2f12b0be0d),
    .INIT_5C(256'h022ffc209a32063b022ffc001e000ce0022ffc209a32063b022ffc001f000cd0),
    .INIT_5D(256'h022ffc209a320642022ffc001c00bc3f022ffc209a32063b022ffc001d000cf0),
    .INIT_5E(256'h022ffc2f42e0bc3e022ffc2f52c206b5022ffc2f62a2064c022ffc2f72820642),
    .INIT_5F(256'h022ffc017003639c022ffc016001d058022ffc0150022491022ffc014002063b),
    .INIT_60(256'h022ffc2f42f206af022ffc2f52d3e39c022ffc2f62b0d004022ffc2f72909002),
    .INIT_61(256'h022ffc001e036491022ffc209a31d020022ffc001f009006022ffc2296f206b8),
    .INIT_62(256'h022ffc001c03a491022ffc209a320651022ffc001d001208022ffc209a320663),
    .INIT_63(256'h022ffc2f1292fc36022ffc0310f2fb35022ffc001702fa34022ffc209a320661),
    .INIT_64(256'h022ffc2f12b0be36022ffc0310f0bd35022ffc001600bc34022ffc037f02fd3b),
    .INIT_65(256'h022ffc2f12d205f8022ffc0310f01b00022ffc0015001a01022ffc036f00bf3b),
    .INIT_66(256'h022ffc2f12f22491022ffc0310f2063b022ffc0014009c07022ffc035f0205f0),
    .INIT_67(256'h022ffc2f12a206b8022ffc2f128206a1022ffc0110036410022ffc034f01d051),
    .INIT_68(256'h022ffc1410020663022ffc2296f36491022ffc2f12e1d020022ffc2f12c09006),
    .INIT_69(256'h022ffc141002fa08022ffc145003a491022ffc1410020651022ffc144000120a),
    .INIT_6A(256'h022ffc141002fe33022ffc147002fd0b022ffc141002fc0a022ffc146002fb09),
    .INIT_6B(256'h022ffc1410014a06022ffc145003a491022ffc1410020651022ffc1440001201),
    .INIT_6C(256'h022ffc250000bb08022ffc1470014a06022ffc1410014a06022ffc1460014a06),
    .INIT_6D(256'h022ffc20a550bf33022ffc0b9290be0b022ffc0b8280bd0a022ffc001700bc09),
    .INIT_6E(256'h022ffc0ba2520627022ffc01b0020627022ffc20a7f20627022ffc20a6120627),
    .INIT_6F(256'h022ffc14a002fd0a022ffc0ba262fc09022ffc14b002fb08022ffc14a0e2fa07),
    .INIT_70(256'h022ffc14a00323d1022ffc14b001df0c022ffc14a002ff33022ffc14b002fe0b),
    .INIT_71(256'h022ffc2f2172ff13022ffc062b022491022ffc0b217323c7022ffc14b000df08),
    .INIT_72(256'h022ffc14b0020620022ffc14a0020620022ffc14b0020620022ffc14a0020620),
    .INIT_73(256'h022ffc14b002ff0f022ffc14a002fe0e022ffc14b002fd0d022ffc14a002fc0c),
    .INIT_74(256'h022ffc14a002fe13022ffc0ba2720620022ffc14b0020620022ffc14a00223e7),
    .INIT_75(256'h022ffc14a002fc10022ffc14b0003e03022ffc14a0020620022ffc14b0020620),
    .INIT_76(256'h022ffc2fb160b004022ffc06b2020b8b022ffc0b2162fe12022ffc14b002fd11),
    .INIT_77(256'h022ffc20a551ad10022ffc0b92b18c00022ffc0b82a0b206022ffc001600b105),
    .INIT_78(256'h022ffc0ba250b40f022ffc01b0020bb8022ffc20a7f3e491022ffc20a611ae20),
    .INIT_79(256'h022ffc14a002088a022ffc0ba26223e7022ffc14b002f40f022ffc14a0e03407),
    .INIT_7A(256'h022ffc14a001d001022ffc14b00323f1022ffc14a001d000022ffc14b000b013),
    .INIT_7B(256'h022ffc2f2191d003022ffc062b0323f7022ffc0b2191d002022ffc14b00323f4),
    .INIT_7C(256'h022ffc14b00223fc022ffc14a00207d0022ffc14b00208eb022ffc14a00323fa),
    .INIT_7D(256'h022ffc14b00208f1022ffc14a00223fc022ffc14b00207d7022ffc14a00208ee),
    .INIT_7E(256'h022ffc14a00207ed022ffc0ba27208f4022ffc14b00223fc022ffc14a00207e1),
    .INIT_7F(256'h022ffc14a000125d02d00314b002b6c90010ff14a002b00a02bff014b0020661),
    .INITP_00(256'hcee1cd4240624346c85c56fbcef4ca5857464e4148437749484ecada62c4ecdb),
    .INITP_01(256'h4cc150df4f55c448e154c8cc6041d35afbdf53de5b53e254f4c65647c4d8c0d8),
    .INITP_02(256'hc24848cad8745fec4ecada44d8f240d8494ad7fe5a53d2e94cd741d65964cc7a),
    .INITP_03(256'hcb5553c76c49d741c243c0f64b53464be1c7c2404443c8705ccfc9ed557eec48),
    .INITP_04(256'hc35a5c57dde956c85644dce9d57dc853ea57f4cae8d85d55d0caf4cb53ccdaf0),
    .INITP_05(256'h6271de75c1f9ddc640d1d1d34675d2dad47b4ddcdaf54559d64ac8f05e47c46b),
    .INITP_06(256'hf2c86f46487d7dc5c16842477e6854dbe6dfd0657c72de794056f5efe640d56d),
    .INITP_07(256'h4a634fe679485bf745d5ec5243fd4b5b6cd9caf1515e7564d37161c0e67bd9fd),
    .INITP_08(256'hd1f4fcf3fcdbc7f9fc55e0caf174fdf4c25f6efe5f7248fa61e0fed4dc66f2e2),
    .INITP_09(256'h545d51507e5b4f4fe359de416748dfd5edd1f3c160dff063e26cce57e6e4c3e0),
    .INITP_0A(256'h6e43f5e260fccc6c55d6f1474355ee7f6368eef7f1f7f476e2ebf1706a71e2ff),
    .INITP_0B(256'h7250da607bd2d26e7bd8f7d2f7daf74740e7f27065e4e667f972744a7f407f55),
    .INITP_0C(256'h72e4725a67ce6dece7da6471725b645fe4d978f758f4d372c66cd3577bc0c1ee),
    .INITP_0D(256'hf0c4d76454ec64e0edcb72fb55c849eb49fc404ed5535c7458fc404fc6c67fef),
    .INITP_0E(256'hebc875f77c41e55bf6426a49fe4f49fcd87553fe496a496a747de2dcea4c7953),
    .INITP_0F(256'heac4a2c7e2d75763d47440f957e3df616865ee467043f3cefec34a62d47d6276),
