`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7568)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5GM7KY5OzTepBA5ST1wPhsbsE53bQSTPPtVbyJZ4osyoYQznwVaCpmZb
begJCB2Ccgtpt2GM78iDCocaIMDiF21pgFG0kpRlwG7e8YiL39f0Y8byMc9SX/0gxoO1EOdS/7MS
QSnQnqmtqtcSHagA90wC4Dtbt0rxNoIyQbIAEKomXLRR8H5UIOtS29pI/BJH4ExfffoFvNvWOFTJ
TAwMXmKpkFu8TAObI+8ExGQphn1UxQnwTXgS1QTlweqmcA27Hnp1U23R8pRxM1zrpH+hDGx2Q3gw
d3FmJKbgPjc3qxPSBXS47NDn6x/XnusKSm+pezugdSdctUYYeAvuxDwGAIMbkkxbAGdX3HAzT7hc
mZNhhtH9wmo34dx8TsJXsJploqjYAY59urPE/yXsrovF3q332YkdqMj1FWnuXJ26mFoqFLt/WzKC
zViq+Dr1Oorla9AU2ZJIfr/Mv/kLzVwzdIOB5ChHNb0Dk4QPQyxZa7TnJrvhvr4aqKzj2q87oamV
7JxQu/PTenK8/JfbrtYKdeS3cjkiQzj64ASC0jBteQxq6Q9/TXHWTnYB4GSRZ6r9Ey/fWbiESDNi
Oqamw8jKedfryhFxsvN/v3/4qFzomR9eUP0nzlGWBiUS8Sx/73j2OWwATWOZcUoWi/l3SL5ReaLt
/fJplX+bDEx1yh0J1byvHK38F1VJ7o2uOW7d6cJQ2A6aJmSxB+rjbFlc6eU4M/8fIINsAxvQtQL0
ROsRL2IQxwygAkMn3Nn8UGyjb9wN9w3zfwC2qdfZmvs3CSMJjYQyM600vgDDXduXBX6jjJO0Fywt
56xJGiPH68JMD5K+3esQeCB2JAiKdqcT9rJ8Ws/sQyr1wooSHPPxuTUWISTuQ4yOhzi/G0XXUnXj
uiI47t6jmTndO3CdxQQejiytqp8jDj8jtgFD+QWItSI9A9tugXDo4mVHszfucPs5a0j84tCapGfM
WmA1GYSz6xNeNH/jKvFEnyzmAQcNMFGpfyPSjPy3uNi/75n5NDkZfY1IrhPjFqb8ArS74zeenAxo
zqhWk/OB4xk0+fzG/kVFLH1X7ALnQXye+9vQStGhGep+2GuRzX/38Xizt8UDs5Uxw/LivUQP5j7H
7bbrH01yXZ8Ltqi9jukzlQBxgs46LQLda25bnmVUd94qqA7X4L3EhCwhWy3e2I1iiHK0G9TcvfEC
uV7gMvcCL7NpR8uyj/CGhXO7rnFRD3YY7JqqUsRLuK9km11Cl64UWDb7+VbenrEtUpjkYgPEX4AZ
tGUM21gFItGDmU8TE9WjCpB4ZC+GxzbhVfiRd0kYQbdcevtpv0aVwUtPjSDeWfn+R/SXlslk9r8j
d9D/d38jBGoixiGHWTXNoJ7BBxNocpqjR4wJ3Wo2T8z7jOieX5pXu/JXXVlOE0q6WDimq3xHfnPz
F9JcJKUJjE/Dbzd1hK1uvuXURKAAygIl0lg48A0UHDAmzDxdmcpukEoGWR19qU1OSymsB5t4Yp5P
ZRZ2Ke68WTqJ/4H3OI0V5feUzEI1ylFkSvrLX9OWanvo2ZNGJyas2575bRYGIy0LyBjKRTrnr4sg
rHFpq6UXvEl6fPdAwk2rxTCMt0y+3iyJcyfmBfwoNUcigSppk91dKbOnf0LPvJEHHj/U+iC+dmJP
GzVZsaJrfMERVYnvkTvnqEPJk/TbanEHDD9akxFXpgkDxhCvZhID8V8+C7xXjXO8Cp1hWpO8HmwT
+e3qqEAp/JdT6xpdBctoXYReEfk4cyT5grmq5DDJyjrQIKXYIpS1O5aLNj8lAsSquLEUG1tPwlg0
YD5golfk9wJ4GCnRCXzWI1/6rw14FR6agsufPOxRyM39lWr4N+Wyz+po90CPveLlEQMklb9yfH4i
zTBJL489xvGwv8WpOucUtXpYn0D/Q0rSVaWgfuNTEAamWhgK2kIFUp27qoprjhBYnFvdHSfY3qTY
iqF39HwIq5blFQjuAv49uWigHnJn0dvg/qkqTvPWhxcBkA0dwjDYMhKIaoJxwAWJJfpFoR1DBXPw
YsH+JM1mE0haFB3ne1A+m7SXRGVa8nh9Vzlc/cWNaFt8vLMDNJ67iht10a6nZV+PLN6dBTqIM/R3
+uKC14OJH6uIqKlBBF3KI6TSy1ZsrVsNIru1wgZYpY6tDyJyTzwqf+Si04VxJayFGIx3b6uXsFwo
kBJiQZjaeMu9xFFLkBZa2RAke+wgUT2on3BAll0S1Z+FSTq2d3T16HuYAsm2fKppvVv0s1izfIIl
MkoifMLeERz11xrHpsLDJGWo0jOC9zkSUZ3walHKMfOR/Y/nj0dTSgBdmPuxYxK2OOfVU6Ki0uI/
paMGBgcZoXxhOeWXTyg0w0W0EHitKVCFC5znjDGbXkXkZOdNMe9TjmHZqFMUfWtLOdUcIsG9GnQr
I20TzT1Jfr6AQGGH2ByUmnfqb4/RF1+7Q98AGduT2R8PA8C9FUQf2S/v5mh2fA3iEcQGPlCWN18J
Hg96XAOCX3yrz+qaJDagGW4uEV0/pl5BLvwdYzm2KZgg8L5ukesxE3+HHZ22XIX8tGhwQjIC0Dht
ex3IY5HBHFAsnbRpf7WcmAEldT/bP4o13xodCNwR/0W3SqA37vfUdeMH11LdGApDoXHm5A2v1ysV
JiacLL2yOGUEYOpE3O0258xhDOTguTWa8/LtpAdd+5C318g2h1Kd4hGbVDLC6OTTXMA3RD1AvjLA
mqP2Fl/7Yi+Fv4UDMVSISt9kGc3I8WZmMKfX9BLQEpoE0x+BzrGH4SnQN4luKgYLndvb2F5ri7C9
/Ri9+GqpQ9Yr9WdZLBrVj/gwNp8s+shhe625kM/pKWp3f7Y/XR4Apr+UQKDHIfL1DtzyoqBaQcE3
8PDEF2SfmfQ1H6grj9Z/yEQAZDHF3wXEIZpA7fr5lnoqyRJGniR6J48/0b4j9VYPjKn8e5X7JQDU
J3/QPDzIJP0E+zx0APz6HbWyPF4JY3RsI9sidDF04/Z0oIEs/hETQsL9b5LE7YJhBgu4SUNFMtqY
YiVDTXulSLxpcxTvAHRB8wco9/sZGpFJcyqQRnq53NdhPbhzd7Kb9CD2ssfh4NZ4sf71XxaQFheL
0cNWeCy49nuTYYnN8S2A2/tzFg+qrBjwzR2iQvRjRdzE2OdSrTR3qKC32JWgdxKp5CjSLP2gVWV4
NuJ1qN8X1N0AJD2BPkITsX1d18j5z8fw9MJbuRfqPIxAt/JBvCYNG6Lby7+1dTfrmZInliYivdQ7
ChQYOsYyPV4LJFNEGH6UHGHI5B9HO6Fk8ilWwN6+1UVzTdn4ozksNH/8Nk9dqqBa6nneW5TAynXh
2BfcCcazuLzQu5mjTv3IK72XVfvqUpBfuyp31ie2HSS92lmHYSwC7k68y1UqGbfKN3TTYS9SeVG8
hFMkbDDtLj8h4FDARy5pcB85jP+xGPLVeZYdDUaXA5HYdCrtklUIoU1ef7NqHgnlk1smHdSgxCcL
iBHx0zSVhe0JGXUziEOVxAt25zZLBhzTpzwplLvx7BxhWrYQ56ebQYcBul2R95TUfjmLCpwBKpaR
HZ0+xf4r58xzkD3TLsyPK5URIZE+1mkzssWfwX2BrasHkhMwRL3zGKuBt8Zydxf8llyFBNrtR8UT
QVVOUFsvDHdXHMr8MKlP4oLZl8s/Ql213srxeFTGa2iiW3WjFQqQV/a7ARXfIfzygamAmL7Zk2WD
8/yvBo+iRZIqhztRoWNZCa+cjinhGZrJj0TLq2+/GajdzuAYustQWpqgAG6tlc7BiINgyg2S4s2V
hiYSS91Wo81gKxvTa3Oiy0XHjWSz7+wXJSq2P5eZ4SV41lNZLVgP+XwOkgZJQG+FqnEPmX/T+4IO
AT1TSLrQ9Z7MixbyEpQH95QA0JPJwnLVZseEsbzzLG3CmWZcP0MK5N45AF8bFhaiSoXwNSRJ+4CS
ETEqmuOB66KBBMSzwgXxV07Cfr+KaiXjFspvNoZbmyZHsmnUVBD3pt4XE/jjjHk92dEdJJEfRiOP
rWZ50qQBrKYZKsLQfZzdSfmJpnGoMTSFZdOsLe++FlDSBjMNUW8SXnpTkPYR+B0hXSY2uNUTXdVB
Baem+rnmUT6xOIFmailN3fmffVH8r2p7xJzDsNbohWl7eOS0JOO7Nh4Xs3cadMJcin+WbQL6D9ww
LdlC30UXUtyNykp8vwILjXjdLUCrukFvr+G8lASMTq8bR6NlEDMSHlIs6sGR8Nt/q9lbY9PE+NEY
tz83PSMgoZeA/FZN3zoeGMmpx/lVJ8y6Oj8Q/gLGmswOyc0WlqmxLUxVENUiYCmDW9HjnZPV2xid
p7LsFvEZVMm6D2rxO437ZT3DFn7xiHHmVK7hTh+t6pj5b27IniEubEGEo/hyDF7TyWMM3IrWuzwy
eNRgVGQkuiVWBK8wyZ8YUOAPIcQ6/N8pSH6rcPvnYffuFYjrZGE07pA6rzd7NqGlq0K16W2DFlNh
5iZYxBErtZr/hofXB54/i2SYQJpy7Yqmn/oP1nmiCLtGNi1VD+6JYsM2rJGNazOuvXYZjywY/AUM
O7tBoSE821T4Zo0NxEXBts/mfULV02vCbQYTdpEaieumzQ3E2iSxbla2b53YHUiwAwYrmaYwr7cj
MWHQ8JoWFgHFAxY0CeHk7MnDHOqzuj4dW+nd5yvGNi1feL2e3b5Y1eS12Y8H2NCQs9pWSAmgzGuy
T5VQI1M6ZAOyhtNwgk0UW7jxLDRkP9bsIzS/TNrI54fBRncfJygp6M95KSc3w4OWEIUtE6Qld/sN
DIvevj0a6P2ImP1s3TuaMSONI5qbmlOnN0CJbPSHxhERydFv2keG+pyoe5E6OHRxRUofBGbc+69y
N+dDb1s0PC4ZRmHAXo+uNtfSdikrFqTVJS5HCe+JpssZPeJV3NM/oCsrzDSq1CA/nU8odub5uNss
xNbBFD24t4pBYaTLYjwO8xX9udppk9MqKqt7GvEZMB22eYfhnxZPHP2Qc8PPsVaOb5dSNvyq5yQl
I+cBgMTKRvFQNticQQFXSZhbPEDL1FUlcySnGjeZnv+y+S9iFiORvWU0g7t+YLWY2wXFJjfzwX1l
APG6hlQ83t7DN7K6hHJ8X5JVi+V97AqubJf0RNYsRqPV6dDK63btMP0he14t9ijmu60kra3nqvaR
9gr74Pcx8O/wOkc2S0J/UXVGTIMYph2EEh3fGAz56wLqUOPT+ADMhbLK+jG2GHsxZ/SIIMltg5Lh
RkdRs5Q6z7Xn8k5P+cMZAgi/Gvas4DAqiqO4WPr6TpnCUtdrE6o1byNyJYwbUO4T9ODN6QkyIWwS
fTsJYnO/aaXNsoNlHZ6P4q7mnAB0B3wpuE/85DaDhf02ggqHjZ+w1grSDxVVpwYElPQjFwkRvuH7
tvhTu9pG7hB2o8ZRawM1W6+T2wFxFwmuj6wSf6gZowtjy5t/H7M/BRZIre9W2jZDkHGL1GbjoFf2
uPX8uwBdBQ/vVj33upB1PhBIJnHhqh+A06CbsKTYgYQm1GkBfU4q/FrwFApwW8LNu/NtzNYSLx9u
UHbhBt7JO0XtFbDUbf+txmRYjm39PYcK8Apm3GJrByIxL3jOKBPc6EWWoFV7pbc+n8/ofylsNbR6
N55D6qN8C4FchRQ2x5XNbaYic9U9B2mxM2B3Fj6LJDpUII1YT/pJebBVE7QUkI2rsRQiryKPQLta
TmAG4Q6aCY1sPJMdLsMeqySHUpWeeDVVsQbxVu7LU/IEmzpegQaa8z2hMorV2IipKztqqniy+4Oy
jYkwcEezQXGhcw6cQnQ0T4H6nAWD4OL/UIcwXQHsd2o4q1OQYAJ/aqC1sviYjFedcLHTdrCrjyNX
mdf2ABZJ5q/B3ZIPVC5vRGHENFaSempQ8Z5qlBZr77zsF9QezaEGBR97OHJbe1b2MTKluHYClnSc
+iwtqbsfRddCeMXyfd+yRdNer4lGBpALkljtrx7w4HdEFJhGctlwVtl7/IxdfvFEqtBgaiHWnV1+
5sjMnkkuBejiDU1TKuGrUob26xirXpQvZt9WXDCTTAwiZ1B74KeNZ8tm/B3cK1II+PTzCEGSOSyz
F8QsLr5KmMBqdg1DlcIjEWLt0DyWk1cOMpmw/35c69osC501b3AYU0qpfjGnTSswdhqgxFwECRr0
gocsqLHiVMfvkHlJgGnKmr9V5wwwifEgDXTQnShOcUlQ7KZUWLO6dNeNppZ/HPWvdi22tbhp+ZCC
bpB03/iblZgFzXTAKikEr4Brhz4XKIcGRbN7+vEcxJ9KptXrROYPFl3C3XnQvSJewFbGlYKdQBd+
T+3XkC4bmkRe8SKCK3IZz3sJvD56vGxXqkq01OfEwP8ecbCwYQIMYFcgIgtj+pm+P/LY0lSlYLSt
0pJV9bxtzWKpZvhNku+l96VpF4H632axp3q4/Fi86qFe7LCfh6yaTVXPn3N+1f3zAG0OpSVeqac6
apuDVAS0S2kJl7IR3K2Js0/UYPGY4DESsPxSFrqB+6lJED5fR/X9eY7l5/+c5mu61ekJpdYsjAri
UXA5WaAzC4hCMERIOuXD+KfuIbQOeN4CirTx0FbbxM6NRvu9tbJrfMsGvBpIE2UMRPmoegyTZKT0
zbIrFEDsT9G/6aYKL76iKCWuQMEnmi8RhbbIJg/WNWW1d3/gxEkSEZMmQWai/f5IwJ04ZrkFLhPA
Mjc3lbwCrTZvX3vUyRDrzhekzH6ovTD6ctgqjx4dCbaNcVq0XIVV5YaXsn5+x3bG8nL/UjnYt0EH
cTer0F9uoYTmJqL8445jbiaFobUYpJyERBuAWvu11trCIovjMTE19A2bakzeBDEhGXX+QS+aJcZ+
uSwqV1tnbnY9LksPJs6ddVkwzCU6DjNzKgw9PBYJ2Neu3LddyIjDm3P7ZiBp6/b98XxWvEHfNuqg
B5ac+VMg2rzVCPS3oRWUmzRS6NG97AnptqifJg+ZwF9L/kEhQ7uxekEow+YiS2Ou4HbeYcSsriAy
NYp1Csipj+p16J1dzC701+KZQBnW8pnFNk0Xyn/UP36goCAl+1vLCxuCVECeQeHDdWcI91+wQyml
roO+cUz4m9ervPS7IGZjx2a1tl5uRq5RGMdsu7doM23QdD0yEThiG0u7LQrlIjMlSvdy4t0wLL+6
O9Mh0Db4D+nE9NQMeG8LuTr2GYC2KHU0aWvlHeP37fbSnfDs/4a41d5D+F+5g0u8L7fi+iWhWpPJ
fiL3Ags6GvTylNU4w8JN26dTaCctGhjvg2AcCCSIZIYJDxp0j/2JTEwaNTzv4xX9LfkTnSeDYyJX
WeBoTiC6XojuEUP2QFsDkNF9+UjuRPc/syXVFdlnUSf8fz3vC5iAAUfIeY6uRzEbllBNC6IjyFhv
e14BMT3XPJxT8Z+IBQdbRIbxj7irjkMKKtX3PAUiNh9Z8nkXpk2TZkC7S0lRaEvibAkbEbkDNdkC
uwYtUq7LEutnbFCsSftiDNaazwq/4bhV9TE5jN6WpkKT/U0UBjtyseEvpSr+heZcZb7leThsrVBk
NnUVSyJMjGM7OSmGtoeYDEKFPwAl3puO45Dsg+MRzCSXk1LCh4fqlBUkhuCCURC5hSQ91w68eoo6
LW/JOxmgmZr+FUO9vuioDhnXYYyo5j2ZG84UShcBKMK4d9w2T2Jp0RTPFoZfViIDDRJDon6bwgPb
tPnRZgN5Dk+tHcZXZP3Iy9q62jQoQvDzKJyZtl/Y0hv3MXCWWrtgoS+zUcyEs0gEqVuxWU0g/oi5
hyYMZS94KgzxZhwJLJoo+j0Qmn3/9Z9cg4+aWoubo8NkFwY4pArq2ixNSakLZKWMPNPMPaRo231/
Dp8Z5wARSAluDmbOe+873nquMy3eCm5hEj3e5SPzx/aS1SiMqITy/VvIIttGDKQwS7PRz0hxhjd2
nKm4Xl/IqJ18tcgZ1bUUP4wo6ysJrjg8b9V68Y5nHnainIYzm+qb8x8y7imRArY511C1fbbYZQYb
KgM+z++HrbIsXtrNZekTfkgbeBT0apV7ctOk7KvVoY1vnGTlQ8rGY39SzBJhsaEsO/7XsOJUGwrx
PBxZ+JG9CkqEO1ePNnw/QUfr+/Sah4s4+zVSxxgWCwc+qHuYN2oOCXqDU9qqa0EVVyu7tEzhy9XC
/+A/nvdsy6ZTwW3Mf3yCyu/2rdNExAA69PCZVp4XRaPyaRhEVESvcutypK2WbPTB5o3sMDTvEQ/N
4y59671WEQJ59statByBhwCbyDy+2UTSGnw647T/q7vP9Wg1WV1QvUFR6r+3N/WaeEozhToz6MBq
e8/J5BEYb52Avr7Ih/ACOwRcQedBSgqNP1lgBnoNTEN1oz74MHzrpiFdx4Lj4mSFNeftNO763VhK
z5k9vHIoVZrNdjXR/GyhQ4JQobO+9Led8D4XflQAziBpp66qtkNoUZx43p4+mL9HGR2DqrZYHGGs
1ozE+b25ipHdU2XVoZ38+Zi0OI5H5PRr5K/ieuU+tLpXpxH1WVcEaRl32BP8RxKaR80beksVklmg
mPatdlZvJg3iEtZqniP3ApH+HWBoNexdrBJtCgIsPm75nQ7EAJcSf4PIIZ98HOROX3DgyehO+31b
mspixGhPSTwPkMeMTZj8IE9XoihrBTtOEHWRa/zAKNtw6ytvDpCnV6bmIYE/Hrk1vKNWPg6P5IkC
Qieu1rcN+TAqJQCAwYwNos2PiwdLmpTI+HZZQONc+Gm+UTroqLdWza8V0Z04X0UpVZSgZ+WuLF+A
yAFWWAJDf6g3oYs1l6sNqLzoznrQCdtZI6bCMgwR2lG0MFomVh5yh9dVfBAc6GdUMPU2pimOS+Pc
CIlev3BhRZRyHHRiMFlv79T4AoO3XTNEvgQGAlIDD6iBSThf28FsK/SUdktmXbKAx5jCRv9RNZSu
+lrszHiCP3Rd4m0UZQSldheAHP4c6+Rh/Ce6mXts/smXPspZerJcxTYZJbTqPJGPHmJXQh8v+e7k
dOKSZ7ObNR8enuaxgEg5oJtVlzHaZzxG4NFOQAi029cz7PBPiQxonR7Rj7NpPi/lE9a8PRrUUgQd
OdvRdBEYr9hKWiXHQ1ifO+3FYZhZIPtA63QAvSNBT+w48tDzJCd3W/K8OAV1XFSxgRY5dDEvSo0G
ent6IBn6mPnepZrjkmCjHczrGlM/UXDshlUZTqQkZf1tAzVE8pqKZN4M6VXnNEvKy0fgaJ14dmCt
XSgXufhde/5iCWTakF/KWTnf2jqrXzUtKslYw5ts64G6kCt0wBN2ca4hqSI1FWZxx5+Mf3xUNykV
+SfI8HPW9+5mbp+eUWoiNrxOGhZaD+z5TdGhB3ZH3Nsf1WqHpQRajXRE1rf2Qkn21Ocxk8EgLBm+
xojbNnY5kStjHhCA4HxavwPiZwXNcqzfliBP2NI6KIj3ZxlN5hS62656qolKLU4coRzhMWC2ykdt
X4Y7w/srRCFLC36C1NV9oWduSXqmPLHkEHQcaN8OMxvQ6BuFMYnQAnZEbmuyBZyUz2/UvBCiL/2S
YrpXbfqqGkn+mFi3WIsK7/tiyR9ukh+5Qa4ucHn0XkLlNxtKIdeL+RwmRzkjaKs+vIdFOtDF7u1I
6ERo0Y1E8t3FiXqAi8V/wzGoghIxX2Vf8Xf6/u4DqlabFc6b3Uu7p4jetxY3eIBm/AiXXSuNdlW6
d+I5UJQ+cJCJjJaeINjiTO+o+k3hLLJeTRqcYRDcBAidZ5+WizLc0/V33ZPlfWtw0V66tt8d8CzW
TBML5St+2fFpj4VEJTZ+54eBo5t/mtBdn5wKAArAzbtAgnO88LSpyg2HD7gVKa+SfBS3wpKMpm/3
BvCVcalSMKSX0L/IPzJFTSAuEjEnnyvzM4UpvD8d1jjdjPB6LS7Gx6N3vo7bICs8U0DQ7EU08cLp
fs7R/20kWE0rUC3UD5LUvbwR3qAjB6aruK55uDPFYNUpOjvGxG9zde9LxZ24RM73V2dgEh3/PkbZ
geTSAGsf7/mjwzl/Aw+A/Zbo3+iQU6tgZNubx/CncAR2e7ce0XWlH0ezggSsDHOfZ+ep+6SqBAPq
7yP8929RRGeoM483kB2Ww37JvI8kowoW2k+TjlGoTZhETCv9NXF9c63BaBo=
`pragma protect end_protected
