package cache_pkg;    
    typedef enum { IDLE, SHIFT, REPLACE } lookup_state_t;
endpackage: cache_pkg
