`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
V82h/mp8FbHcv3//3zVZ5VW10Mue/LSt5dvjsUkiSGtG5WaH8H9Fv7j37k+xy+3/pQvfXcpqBF/k
iaz4/vETUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n4WSOWV3uUjyMD/l4IGcKD1bHONRRplCKgax9lu4YRYlORLHEpckVBvOD9geZHtnlLIjTLNUcuHS
rc4oO2K5x66eEf5+m+hNzaPYWCrVKWQI7/tyX0imMAsD4JQXzU2CP3ATsQoldRyYOQZmggmbIMiB
stLQ3uoRuVc4t0kXI7U=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zgo3FUzRcS1G0FRTCr4C/JBs44dp3dv5CUvkYU2vM2fDyGtu9ekJcjDXnFGi3Qx2X0BV1gEyWxsJ
xqQkFlu/f/1mutspkUjOMtKZNCgPGDHkGfwBEPN/xT22fOBwQJUR+Oj5KSeDWe2U4t5UJ4XXcGMb
ZV9syPFreDWYOTWkkl85cAKcf/WXC6oz+tOUowqV4nSLA1PaSrK4ohf8oaOGNVX+4Ji/w6ViTIJJ
OqmPJQ151npm7Kbt4RW80tp1OmABkNI+o6h4rwtTS1IHzM6bJ1Krrp0V+2aEmmqoZkuKINjX5Pw3
P4Vi6iUmJI0uMpdsCPr3MEC8HH4v95WCnjh0Qg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A45QQ9IEoKpoNXpmniz3AuFZmGAAZIhtA2hP4/pi+Iwurx8nPI4ZkKpYXPnn4DfH42bSsec35aiS
Ve+A8f1Q00bmFgtclspinRe4YgFesk40ftn1mzy6g6sLCNXhUm/IIjCSNk+ie6jVQS7STfOdio+z
cvSm8QQePoJjzlJz/jkNhsD110PhDAevJWb+C5fforY6kT0k7ZmJmE7btahod6wU3o7t2HM6+XGU
DDNZ5E+RLS+IiJYVCOwsdqQFDuRaWwS0k8Mk4UuDiVWtU0+QLFZ/8UGJhy2ZDSYlL/8TrrsWcD/1
Vku2N+fkWCj38RSMWEEe5TmUHSSzP7uBI6QwVQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b+wEsHDGMmVXUM545W/2toIjDItLsHFsIOyFDid8Fv6KhzBePVZlc9t2c1LfdAa6UEpdqcx5kgIr
+oVEglJG3R/fb6dRp2mvlu6+x0AYh7FK0My5t84q7uKZ6EPBxHnDds9FLGQdMDUFv8E10WtGrG31
lkto5q+L5WLAzYgiD3//MgdbP+aqLc/75XWIRhw/PfRn4OqyBU7xSBeoK9TDxBwOscUv0cQ+dauJ
dUQ0W2ZCXwF6cP5c47k76Ikfu69J0/IO+FTLKMkjAB7Wzsyqbpl6RMVdJ/iYscNROh1xxo2k+52w
4l9VnVKN7wTWZdW75B3V/MsNTrKb2I6dBdveDg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyn/owx08GdB/M0CwlYM5XwpK1DLRGgNdNGvCa53fvz5ftb1LM2R7yhWTTXlm8iqXlg1S70wvPmw
WVO2ZNZ0csmDdQcX4HNMiokrI2gpR08Dk8n3nzdOhqyFyh79/eVJzQItyKMQmJZNCvFfww0mtX5K
FbNe2x6ria5jEBEBp3U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J8WwILioFJtk4e6vNsFHYZhWTjvAMbsqHcnvhYKYzsY6fpaoYuWnjTNNNxS6JYZj7bKOFgPjdnBA
rKaGPLghV6UU9fx6UcBVLjNOj95AU3CZPEjWGC/GqjGRPxOkhGtDka91PZuOBRTBqJT8F+5qIgQR
vO7WJHaKezpaUm2zbeC7+ShM5p4Wm9L4dzJ1OuUGZNm39p9FbORAZNzAWa35wpfJ6PPOgATFMi7Z
sN0Hg00oxMFCKSg1bxvN3p4iC3rVT+wV6yuzOecq97B7Fu+tfvP+shqnUhodTpF0WYfGWHeK9ocM
Mg7nt62XJybi4Tm5rgYGMIIM0i67934etK5Aig==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AF8EDKLpUnsf5U27caIfzjHsL1dKCT4FvrlOxjBwD3ZJ9vsXwbWO+EJTOJOFymKnoSSFnuslr7C8
ZCAbkJJLJrLXJwfvC9hiPRksxuYzuxWrtwsjJd+5KWtue3gL5kHClD8Tbo/V+Dnr3gvKzMRNdFRz
i+4p8dC6/32xR0/NITJMYT1uOYu0oBFDHGLR02Wn4PqghcTR3gQMVeL0RsDhJibeNnf4Q0NsKqCF
7OscDpis6r9ZAFao+mdpLGI93rreTlZvJBUPh2RcpqOjL/8IUv0iM922KOCZ6j1LtvD0igXehvHa
5hOx0DDcMjOoejqJiwIqLij0FB13lDBsu+fjWw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 139136)
`pragma protect data_block
BMP9G5RAk03qFRu5UmzfhEl7ZrPdoJV4zXjowSW95Dsglh6Eov1jbd3Ns5GU4UI4S6U9hKz6RpsS
CmOzramvUP7zVlmK8E622eFkoP6iziq1Nc8yKFjmkZOCwVc17IzqkfOmK/7uC4TWUeB0/0aA9MUC
m7cTHOe4yqM5jx16AuZfIzjQIMv7Y7GfMlmoYkhDj/H3Ox1qiYWXzJKmPpqPIYIFdobNa2FEYP5l
4S/p0AZgAVqh78WTyG3JYYDPaFeU9DRTDnxZyYuN/bpnId0OdmBJTkqz726GbHAR4aTZPG8e7kHx
S56rEN2+SSOexHzjlEAXOgj+aJ0QGn8D/nC+eZb2ls8x3i50f5lGCLz5E1cFNZaqVHgf4VDdEjw2
N7ubLRn/FvxGc+Lx8EQQQ4qWBlmHBLpML9qMsseC9s1zkz3Be/cmhkl0fz71kV32RVwSm9F0Bmsn
oV2D7G8Yf0U+govm1u+tWnUObu4iYN89PSAK+zgsrhRGooo/IQiSQ29q9FO8wI0uiB1rF0oWbjUf
Jr9j9MwrcPy1BTT5tOcbxqG9+VMMHT75E9AnMTbcHTFlBYtBi7T9Jy/uK9yRBZHNGkqMZX/AA7HL
vWy/t46TahY+vjyJWzn0JKC3wnrgRU8o/h5DalR9S8LzwL2lUid5r/sU7zKt6F2zbJTXcfeAFXy0
/WHw9kRbXbbvcxCTkSxBxhTJAOa8nVJUpC+saUaCDDA6OP14jGj6zIJOhFtPKO/RYODcYF6YKgN5
qBK8QmCQo+A1Kp10bPdEvgWhnWK9VjWvCYTFRksc2GqO2jtTVyui0gtCTzUEV8Xrge0Adwe5PJ7s
XoAqzIZsneXy9R0W60ZZX3AsUhTrhizIgN49fdCrH3f6X5L2t8SF35qm2GaXC+/JmR43nibiGksq
rldOCnkuGVvTXkHx3RCreiIODfH2ES4lFCtGQAgpPjvWZ3YpkqWJ5au337reigFgENFysfh30dRb
E64UGjJcFBeYRSVh98EQ6RGVqMcMft5WE+PU849Ajwu84DwZvZyOYxeagn6w04uY3NqDw4xDLooO
vUBpOmW6+JqqjCpds0tCQ5UrVfbzDj1GhIyEnOElD31ahiBfZsxXiKUd0WIN+5nVhmLIY8yOiisO
49P2oxuOYrV4oBXdO8sRZWHTHmWcgXkPZr1x0FeardDEW/ijV7K7Au8xQhScUcTBAxnZGIM5nL/v
+/TXK6NlKK4/+pys+RVYzouMczK0PqXsUrmJlQUAreDr1Msi4Ie1VRjQA5CAHbREMzaDy1AR9F4W
lQ2njpkHJStSFX0i2YIwWbtafAams01mL9Gzii7yjDSz4mHG9Uyq1A+AeyT2gmnrBnXSYGk5bckh
CEhQpP+PwSLluqoBlt7B0JwqK537Th4OtTSEu1XQjFUE13mLAYXHG6qGABFA4WnAeGNBD0UFeETp
H9Kt4X0kkIxgPuitCHz+23jh/PnAlotz8YGHGNkF/PtmXtaThDNMyAbfbAlaavlYUdBm2LMVGbB9
TCWKWEzqEl9MMoJs7qwRRl5PNbR6LpspdSDICTa1mPA0zen4y/YwwDuIyIY2wFgylNFgJaakmSU1
v84VDKvxZAXIvmcV78BXURc2izXYGtkyf2nsfOCPVkrUzXBxHMTd4RtKT5cOY3IuosYbAqXGACEX
8+lmZfoi89THKSF4ZmWTophR4xOqAVm26BOZ+Mu63Yt/YDrs6izE6M49DYInGOMmfD14SC7ILs4w
x/K4Ygjpa7D9/rfQaM/wr6VH6LMezkwQmVG+pckyHEA6ksEBF1N9SsX50qvckQb7E3aD0iV2THv+
MpRB3PRrx4XcBlB8XpGHeZBI2gJwNdabw3P/A2BcNxGbw5q3iRLqTI5XqBuYMkEIN3A4rUwsexC7
KFmfvyBmBZBYAWLYgqhLfs8uPqrHC0XBaNihA4fBsnOFW92rn6+GUNE4lmKNAwtA4ObqKh+FRVyw
2+vPv3cjX3YuiE0zPQ/p30V0tejxTZhqF3VZBb2Nxkk6iB2oC1q0FbZpZRPfXJXWcLVO58VpFsO4
VwSGTrvhYA2AvCeLpnID1UnV+yyQ28E8WC/KXbisT9s1RqUdwEeAgwDXhrflYd70hnjzeGbvRAJI
bLH07pXIHZB1kmc0qj/useYyqyG+Hywn6Olo5td2QkQOug8lnS/sTWWZn2tcwWLykIT9LR+v22lJ
0WaTnkCsHo0d6IXylV2dzisHJ0kO/LGoehssyAkFNgOFmSvCcfdflzi9lXBlIGVXuOXnczStJ3GB
TMxDN1WjTxmqJ4Y3ZEryarjxiOi4JxJ5wpOEt0tX4vjWTT9gB2imLEBGwuamFrasJXtv6rItD5JO
SWrBkDM0lgXDGTl1b9z+VQpM0bDCvSShw5P3tkqkR5Yv8SRPOeRheiO7OufVWA7vxDuWxZT9r4os
6DlqXu1oHh3GOC5bLe1kFoNojYLzZnf2UWEleXT18H6prYY+OD3c9tITBXYQPvV3kRFF1Ze+Oo5W
0ZsELDuSJPpmrJCD8E+d4duiX1tx/SBeV2PYmz6xxzT/gr4trz0huP0jpunMv2VziNKDr6oi+1uA
5JKwpM9gytQejvVTkq/VnHkod6CaClT/vTNbrrs3RMZEM7YZNOKjRQf1+D6lS/VNnTgfWzbp2J/z
djadwWWlY9VMEwflObI4W2u2geAglKZVXgUS1llGIqv82CJHP4CsPPU/z5g890NPJwyTfWS0qLf0
kudlfs8nVf1etko4eleSlHAwkf3XTTl8pzpqj8oGrsS2VECxbgQiJBVCI66BTBaBkGXtqihJKRul
N5bCTpfU7EHN/dbDSYoOSbNyl4AcaDWoqA8e0qxpb0UNoGcn5oREeXzNm7kmZcCNjqix0TVJuoQP
G8YcSdabAxBkX2RLxJ9vkgWAZlaGyVFmWhdhXlausk9u96jHr+q9r0xGSGeoy3eITQJOkmDt/Dpl
jZFBlDxNbwW6TM/iKvx0iwrEEIq8BWNVjRFphKLpIkVvQfWBtJrwi9dx+GxJwoHny362ZH1x+Lhs
8M92olueS9P6chEkfWWM/2t5GPh3D/U0d/JntzH5WYyPb8hF4raqQcaj4RVrJ/lPhwULH5nYrEgN
WsVJcbYHkY9jRl0rPj+pLuJ9HOVarlbUggxRFfmcLpTmJW+/4bpjGw5uI4BjuE/c1+Ly2rW8A2SN
v6UnoPYsH/mSM/LoHmk2N0x4KKeIx+ug7+CyZWrVWxi57U+b0gfRUg2nlLOKtHWMTMbdJzgLr5/h
fK7S12PJHnDAtHbnWepihfSV/ErmDae+td5yAf6jLMOGKaSsLUVFw3rwwfH1YhK/0S51mjH/6e7W
JjMNEJSCMvRmWulSOmh0foKSY/KPTHgswjwHI/YSpT/JSK9S6GxxEWZ3tp6pyAIpK81R+ytixhED
Wh7T7qPXszPTtjr+AnNX1sEnJh7F3GEQTlBMo3zSO9QLygcgWeEqZKjmmJIYJ1w98OT2snsya+nw
xGcP5LaffU+F6C5Jpe0+y0Q23veuVcEtLn8Q4fil7AlDLa5+JBtnp+eT/4RaJmBA8CnAk0HQH0jm
IVymYZWlo+gUTWFZYAlO7IGxrkO7KN4QV8HunvAtWlt8p0c8y1gvhSLWX1czijZAx9pYON3JIWUq
o/XPwfQGPK4FzDQ7vGEPHsc5CaYPhylvZtHPZrwwjFOQa5ycpxAIocVeVHi9PAkI2nmsl0keGd8g
QptKhAuOmtMgH5g2ASNjEIsu26ikqz/jeQZDbKCm8v0R4PCFVZAKQi5vnSL/KfRRAesZ4jUMg5Bo
9NwzOcOOntngpZIvAFq4nf3LiWHrfZ8JgNyqV85Pdlxzfg+2LmTZOSZuWqJpDdobrBQ0/nTzfMl8
07EG5c+TDZSp2ohR3L3p/rkq0fDzo0tHpXBSBpyUBTp8EZvpd6v2KD74rac6docQMPgHgpiGaOHy
3r/XhkMfb1QfCzLK94aK673da5vCLMHcLd+zVCLytYUVF1/emkFQ2VYWWc6u3hcOXG6IfqSiQ9s2
pR8c6LbhONG+332pXk9aCrpnREO+YzW3WT+5HXWIfGcea4n11W42d3sKleUw3aB9wQglhSKBDVMh
9dOwnjre13XxBHe5s3v9Yo0OVbXYyDsrTmsuziRW8gI/RJGtVixQWQqJyX155Gz7eicbZNgzKiJw
Rl/zKZEqN3FejJpMRuixePd1DEu4zQDccuj3GR353VmX74O/l6nQTq7WLlJtmoe+6hFywUh7nlTx
trx+/BSOF1R/wNfh/EpD8GSaUgU7E2OoIwy9eMFMabXHHvfKI2Mf5pXbP5HvXXAoAmzlUV48xKwy
NEADDOR2zUgZad4bf/4noLHgvZEAea+QTY/DOGqxn/M1bFkkj8ca3jIw6ZZ7htP4iWBRwp/Wjq0S
6FSfT6ZIC0Lf5fWQKKrFAX4Hj/iDpJ2Zxf3xmiUZBS77EfhxWhxvQa5INJU7NNIoUHJ0HrfjXuhp
0t4H+BQRMsno2EkEhk3Cav79fKNxVvHlGC34/14LF3FNZm+nq1h8R3olVC7FudgckRXqJ3uV1IGf
2GlPGkG8Aed1mByt2bCQdXHL8YRpyFEC4lvghDUHhQzF+TCCWRq8Eiyc2tylE2c+ucwjzok3b3bB
chNE08SrIU7n2Aj6s9w0i4SUM7ycY3EtGepSzvh3ic/smNvj6QZMXTYpPOgSufB5Njnu7ysdr2k0
IrKQpga5SaH+jSL/NLQquw6c0ptDBK1kr6Q1x1035fFV28JdrImq1p3jHuaKpOviqWglzaTQ9wTt
RrSv3pUhqh6VBDghPTuO7wO+4Ue+b4DKhZypWf1pISP0z6xHAoTp6g6ygdvod2cYwwHTpZs0k+AM
noOfNxjQytGLPugyS2epeYD3DsrCjxdG+5DrVuzmQGtKfKDlhG8Df4jW4YUca0wKt8EpjJQXwm/2
JIxeFH2J4BCQnsShTbq93zQrwmtTx5QHImK1uPlbvZ5uhXvf6/4SkkT1twzmGrUC8T1Vlq2kJTjY
FJKliyFnmCC71ApiwRD0sCgEg4Wyb5nMXsfwl6vEEddSjHJ57NFSETyuuAjegCcnCTPeZwwhtDg5
LsJ94huxes9GOnhET9qvsdBwXEZjPYvlpzMIhTMy3zS9Xn+AeK5qNJvekWRjMqFUs80L5I9WWOTa
+ilDDfJTold+Y7baNVgH2qgQueVoS0e6edcKosBLYBKiLRL9kjtkspubC1Bx5h/00+P5CjAKOMIe
PRQzoQc3ZeQiL8q6H9IFvW1L+kTznbyyKuby53nrRXFO3FP+SpM/6YmIyxuZq677lvnGUHIpO7cB
KIm0yI2Ca+FHB730rGZXoUHNWkkfMJ5PaalSd2ENYebsblhUWSRbjR2nJ4418pMUpoj9vYk69fH1
Ke1xwaiAdcvpw/r6p2G3ugBud6UeoVy7aniI0xVUw03Rv4E34TSFVxpsbw0Kz8QsZpkA2UjISNIE
gL12lzF3l2aFRcpDpUseneH4k3XkKqCuoB2EdTlzQOi0fWwjT/sn2yYupadR/+MiSJo+iDHbaqT0
rXhVXB7eizDF0eiWzdzhMKOqvDUSTRcJrRmMZHU0UJBWdCjjcJQbdN2Km74xTq7BG2D29MUDNbz2
5ObfvEmlG7+Fxm5YD7uweh6cSfPE0ou3LbPultnAx91n0S1cO7ck52YFpG/HQjNlZJBTsp0t9ihq
Z364WmDenWja9PzW5TBlSlxEZN26JAfT7KgbrlJOL/EDI8iFZS4ZijyAXgBEyShlgKOR+DCfhQ0x
EcsxhGIBc/YUXQ1GfpsV6aRmeCvgM2jh/5WJG26Ckt0/V3YhyhmjN6QThXHqTaHrzegS99fOqLZK
tA8drXl408bVdUSqGu0bAp1p2c0g/xvNtZrSU4OSbPE1oh2OQlUZeryDUGJbnZ6131GUHp3lGpdb
JVGnnmKB5lA1sOup1Hjbr5JGJTXurQKDXArIi5sRc2/dSkmvMEmWHv8Fms3V+R1OVtz4/vs2wa+K
n8CA+IjcdZTiuMWvQ2EzqA1g8NDFysraIP1opQtBNcq/mm2XxpWkV2tEwH2NF6cNEEeYpFjSEGbl
7kj8jsN5oXxuWsTB4mUo6fkh0hd8mlX81z6dgNStdyB7f6RcWK9UYDRvLvgMRWZbKfJjWWcEMAfS
ARsYaC5oR58lCZl3R9mVPbct5ACBqn5Obru8fzpItETm8lqkgIy9nVlC1XcOvvFFVYGpXO+3EaKG
v2EV2mPnE3PSy+I9s+x536QYoSW0dtYlAYPLK2RgwNz6c+z8j9vld5PhO6F7n9RJo2XkaLgNU7jr
S4THuI8H0YWfdRdgIkQbmavKi56It1q1eIi0V4V/l3ONLnj8tOU7S9tw6ZRoYomUxFa4e17LdJpq
rUMMj9EifEdmzrXvik0I0R94yilflY1oqbwkAoFVrfF5qYmaFD7vTE6j/H1obmY4lYgb9VwxDnuV
K3cAi34hYjS+/xtId3yyJ5nXv209xqO/GI6Z9u41xADjeNECTi1jFHA/C27/GAxBbBtNyW+ICCu6
aZ2I8l7CrwlrVgk5EjggvySTJcvDdm3yui6whkRQVsOCJpTfOm3pn6sM8Td6XzZBHyFmcX6dUDhM
qknJ+TCt5B2/aEEES+/JGWxMyl6P6/5kYVZE+Ho5xqu0zmAjohWUk19Rtx4+tKFO/Uxu2EMRYxpf
lqk4tcuUZz0+uycwjv4VG2qPiOdFSQ45RPdDD5z59zTIx3G2M+Ni4gjlCvWXGAxABbnKJUsFYhXt
FDBSMwRyk+Ywq0ZhKr+/U6sfwPVSlNtL5LbCyiDRPwP/2HymoMzSxikckYOJTQyw2e6DhkuKwo4M
FjGSSbosgdg+S4Vdwi6hcXitPkedZB9biaou4EYLYJuMX4ZV2GPcTymcqOteMtcxUGvmx2I1Dhoo
4GuNnzVKGsk8rJ61eQUNYIPOLymdSWaP1monNPrKAs4xN/OeWMjZ9PWjJwkaUxeSVgXGmfS65Kps
AQDVCTBTPVmDSJvnQho6E+r7DC0cmbhOpQB8niH4SsDrxXJlllXT8LXVLbkunQEQceMFo/JkuQdr
BtagJiJeSY9Kvs8ZSGDmHXTqbrrlFa+dpuHYwzL6X1z5iVp0i2GyLVE8259yI3YAVTD8qaxC4Fnj
4qpVwuyD8y+bkb9mgYmUtXlXSsb4LwUV2if9Y+ubTLkmQ1Zt99Dfq6dWssOcrU2HBYEVb5jmLTwU
Tw9AHjgqU+iTe0JKIDmSgDJ6rLrJjC2/1+8NCUEWGq637frCRspScdQ6JSx8GlcH6f7mw5WFJjpQ
dAEuzR6vd2yeyZUb2ZamkjyGYyXXWbkels3S9cGbVYQLAWnTBnJwzkHRJv97VWr9vJfVHeCERMmh
1RRUsM8ktS0CNul1ozWTL+Z0gu37b/yxR4Tjhig2oWo92bPdPjfUltSayXZbYwvIUdFzckD6TfNl
l1kMcVgiip5iFxhN9ukGj3xNxAFsyXUIQxTRcC8I0WETe3qxkttkm/tocNKTHEn7OYtps5uguSpz
H0HNSU5kLUcymy12pdVNcjZGKg+K8IrVM8R7RRIMU8++IQvq9JNWlrb4n4HJImgBg5CYnuQkCgtm
iUYZVtvFW5UZtURwmXH1AurycSM6ouQZBtjLw4YumQ29X3whazSU02PRXyt7vqdWNpBlFzcCcQgj
hxXWROnUrvi/at4EZOtYqvhs8SzlsoEYJuOb1Gnku8Aor8UqZjlI1vPe+I/ykRB0ZnQwbLyyPVPa
tZQwzZFaH9VoXmiiUrcZIUIRORYwLtNZjVJYmPsBasrHl4w8JuvV+c68xNEbFCpbqUlEWGve7Zj+
XRHMngrcD/LiqMf4+rnmfttrEJmube0tl57g6AAKayR5D+FuukwHyuAMbnr+cI6nPbDCXAdN1+vi
YdUpSmwxoFDwUDCiLcPsghgGE6mdPiVuSlDym7ZofquNNAD3oQlqjMT/hasb985s1XtBqsls240H
bVHSboNHQ5NRauk/x8B+gTlCDtsUTwFttf0hp6D9e/F77HP4KkwqxCn4WnNKJAjq00Dqs6egAixL
WjHtoehZuX5PkbMDMhK/FZdJnHqcs6v95AqDrnt+tWcS22MW4EmaJgPq5F75xNCiQ/47NQogl12Q
rgqaih0HZO7TPV/tsHPgbLLPcDnHFyfA6XxMjNSm5mD3aYMdaZfqFNUMhezqciwLURcJm5XHHH5h
sndCZX+SjdW7ZuEAoM2VtP6Z+TGIE2Uub1DVfQLhgfZz6VF+CGBjub/ucj9TGFSo/8BCRgVNeibd
ytGR+hKBgNjqcEZmCGVhDiMtp/P/dzc+Obbs15GK/LlJYj1odIw5GP+TG/esDQlJT8gPefUY6Jm4
ETmcndogaxz20tKmEQJFIc9vgCfSnb8EFQAnPf2VWjDHU/SXabcFVHlKhdK9WTLcvOMEGjIU9Npv
cYy19BR4Jc7WCdVbcaDRTZ5NFEmXAYbdD29Npvdr/RSHyLbmznHWztHtXdcnfqgNT1PoXZujSdrW
tcz1NETNDLX0D3goW0ljc1AouxC3Vz8sG4oz/TlVdqErtuy/6bW0MFrSD2dWJIhEf329vZDGgP84
qgJydPyg3fJEmMroOZGttZhqWm9C/SrE6rwPl8Zkqti8icz2g2Vk0RDDULrcXUwf68J/3dfnRzXV
Sg/+cie8uhCjlGS/x5xYKfvBGDOWgUJ/oHtMzWTDgWyC6yRZWmLIa0yUxsvB6ITODDtnak3Qw7Fl
L6vu1pwVTIca5dRXIQzPglDpU30mdxgLXWi2GklbkOU9fHNqec+L7F9wn2nOfI9aoU7I3/ZPEz90
q4IAUCikb7czztGq1Igyinz2kv8bZRhWH2AaOTIqwYPk0EGAho94tqNaj9xYRjxUlB0t/JTL/vl0
3yIpSx2lNbI+UPTsQr7qeHdqVgkNMRqb7l9rPQetVifGD40EKhBpgLDxWXxZ5IPt+pI2MwQTcnfC
LrEXbIa8nj9hbvMmf/17uClzZCWAoQu/yLYRa/CMQpCxg9F9n9CtEt0J4yARrr/tNru7bsTROQ3V
M/6zgCFD3rMeYHWbVEUmfZrcMv+ebVqU115Go/Xy3+wx6La1VTOdH8AZYpIqgARpJkglUHm8ZV4t
rXPTht5vJiOJs+Ffsi1lDwMaHXc1GF8kG97ltU5j1WoIe9Q/C1HiQ7ZWDInWU4r4f4Wd5wd0DKRy
/YZ0nTbAgVCgrBXpis6y9X51AtnJxffklTypuRjY/D5aepMacsBabmAZgREjagt8rgw/hztRBXHG
c3P8CKqmg53IMhMDWv0BL/mSUtdoHQQTb49pnmMYz1iBgd5xVEggX/9c9PyZUeVcTNehNUOWqliA
P5pEmA7klqw/yEbML8w5rPqeXxx91S7fbbzCaMULOwDbiCkh2DPPBksDJ9pTz9Xw6JZnpufyFSIS
rYVAk5vjKQyHzEn1iw6xPFVrIK9iWYmnmM2VWJClZi9a07Plfrg5nj+ny8SQmH4Y7gCUSN3G9W8i
RH1iPf37gKERvu+ELyCMfKRN+5Nt54G7tWFtgItrom7Rpn15fCUacd3SqLHW4q4Avauq+TL+FUUt
m014L5AmGGICYrpHJ/nB4HHM1V7LXPhj6a7Iny4l8eRgvmaFVNecUfA5yTTIKSa4piqaai5p6/9b
Yc/yYQHTm7QEIADpa5Pz6z2tZz100gc03w/kxFdoKRhKXJuAqy2IZ+2AFjw2k0/xuFqZcPmwt050
W2yNWOgcGwhPereu1WoYgkIthXmh3U2vG0zHNim5yr4f3YJhi/G0319Jw1leSz+8yn/GDas+0HlE
wp3nObEHpJf9z4hZGx4mvmMDGErLY4mWKVwxtY1Olp/Xir4WKKTC6hCFMRHH3TjXzmIGC0ETIR2Q
bjkMWnXPAH4uHLH3Di2PEx49ngNbvzd2vykUajVUwGhbhbA0oWNUBiX8k35AsEHP/d8w5UXg8V4Z
5kICYcGayFoWs7Zh8bya/FSKgL9Q9cEqfaAsd7Ic+mkGDgj5mJiJlgc6LDj6PFXiKPPLtx7pA/UX
2dy8nd3KSungrtmhvcZxsh5xZL6CC612LQDFcYD8/aUzGbjD7ImfZtI8Ng+xqZ8B95hTbk8GcJjl
cTX/WWTIgD1+jBxd9fi1GNqomUaek+BdeNORHD2uKkhhmXjH1PrENT2/XFH/PnFEEDkoWdfByOmc
nKCpetrIOFZJQIk+UkpyERnQBnmOhIgrtiOQxNHJZtS97bgcxrJdqo4FTFh06I6o68tGzkIfz4q+
1Fu6obbVznB/6ZszhtC1H2L/Xa/9YPWHfrnom9/fYS9D6Orjckqlg3U1///M5OoxQAtzgm0rz4mz
wIVagTG5t6ADmcMQucMQjtMS6EIJ83TDl/5eFxqQHObur8pjlzft6Q+Taa73Jlc0WeOG+Q6Ornfz
ZJvWk8b1kHH6nBmzWNwsNQzGa01KmuuPw+5wFTGXPn3lHZ/HEgLYtr+4k4ET47IgLKOLDJYF/N7X
sw4KcEvVG/J9mII2aMMnYUUIHNRrw2KlKWOQV7HXlg1E35KbJVPa1lS/epmofQVdxyqm34J1EQrt
iOz93tzh8m7LmCJPXUzxyzSci+4co0P4SNhec5lc7HmCBHIuik1gjzrvQ/xw9kkj1ljh7aR8pYTf
6nbLhO1P3pFkxr7rOW5r+/jp0Hen8nZ77sA7Ft8uCoFPeKVHahykdWrFkAG4aU3N5+TuGPq9CuRZ
gAx8ZAEztDm7e9QZQMYT/D770NfBNsbOQvGFRIalVQF0hGrSjR62l8Fes2HBVgfpgmRuDcWHVNb/
XtFWT7uo+ELeHVZ6s32A1lEbPQThsxqNsN7Fz5QuN0VSqhhC4IBgwbCcb5Lpd/1RWp9BwuW/2EJv
/N5uwvVj7FSoYVOKlVNar13iO+ssgTXJgHBGatAmNK4hL3/S1ICtPZNzSkEupaRPANzXGvOFX17A
UjU6G+AYto5DFZ9L98vaFLzITNEhVPElKGY7Ou5Qg1KGoH4dibaG5sH1JYP/yhdJejQ7KnVIrXEl
I4OQAtQ1wtk/3AIhlfFWInsIKCWkpr3Ufn5IKp56mxteHhffvMyZiUYp1Ru9XwH82WGi/BIZnwHj
n7vwmyNwUB+HfcB0SsjQn55cR0blHl52+oeAU6S4iuxFDQTseqaYpRwAm/TwhwicFAKPt9///ciI
+CE7u64bXflEUaxqSLw8JHqqmtbrQaQUW5mKC0X7m6jdPS+SUYlXJyqnRCgHQKhKOqO7L+/By3dy
y1MoIMSv9XdtmPiV14UCJuyhA0ebXS7TdHvAH/66bSFsLeZUSUfVEuBt2C358cQ2vSyMbOgMUPYK
E3n60E2OrREPy3ulmMVnYyaDhe1Mq8emhWj/VKqPY0foDxDR9DbW85f76f/i1zYm+Y5CqBHXjOfP
d7mQQnLeB7Canc4LDKYNbrL5lt0r8l2JqGJzgenzki0Yz+qcDMdERtOLgNDlS2LZ7+cCWb+Azwjc
7+tZEkKP7G14BCXvWYiJEx1pSriiGl8jqpVpL7pqpQarKsOyfYjoom62JPhHjG19DubdsVOALkg8
ep4aiFhR/xfkCS7i86sXbuyEJrbbWm9ZbQ1Khpe/wJXGFq/GrbCnGnAwT5nAKgu0oHEpYMTEeerP
11vFARTTlXWGPHGcd76jVAXzDb22ql3nfcNutWegqy1ljl6QmgCRfbxRCrm2KhsvVDe9DJadxree
rjA/D9+ns+G1UR+3rWpNl4ugpD0PySUlU9RPsVvvNm7MeKXmVzI4ofbiejENE5RuTGmL9FkA6pQB
iBCaZQidqMAOiAU6Qn04ORFRQTc+V/YbdQUsdwAmPHd0k83HCJV+LHyaQ0GtG4+lkc2FdeLorlfx
LV0p0eIPF5VSYFX2duE4778WL7y6yygxD1wmE77uIZLB6KNmvAkdh6BAFzT9UeLEKDZCKkHMhWB6
6Zd3VBT6tv3SFZ+5f3wuprnh/IHo02+yqP2Rjxt+nSoWpegcakHmkY0edP+1rhMAkNw3JdSNyn7h
WZT/qWeBnSB1VqLwx8vIGvhw8OjZv0VEJhsVhtMRZCmuT2ACr/cMu8pRoAwkRvs88lCgFEzGBrT4
wWnAL9XskOJElNiTOro6ucKWxxYAIqxeIFAJOckNtvvLUPgfo4GAWbUvENFfERn+R+MnaUWOBn7R
uYszwl9+ZZBZOnwykm3ZO6tLI4vqiAnxANKqGj56KCVTxoU+bNe5GObrj/brQDiviPOyIwNLUY8q
qgKxFLrcCnTUW1xy8tSeQjgR5jlOJykyZtKB33rs1Iz7G/XiMPb1bVwqYdpoMaOvWSozZUlwy+TA
cnJYSU3LL1ra64XfzRIN6dqYqqNL4gDXlhuA4Hsm9VCFhD5MvsYBsrpb0ddyP/xDrboxSsvD9Md9
H+5g1dNeKGZDIZxGeb3jL1m9btAkXleryDlOG/CHlcD4EEMVVQGxS5DgLseDEKF7gNV5uW0XIAi6
Ed/QiuSPWxelFnCBdIDaJYPoDj7WbatRzWr7id6LN+UgWtq0IdgJcJA1Ot/QdlmL89Rjr0/4T0VS
TrWjkVj/CHaKXFsHW/GQoMN9p5E+YZEV6Urh34ROfE8Ned7uGR2aqAeD3xkp7JEw64YDp8l7wzDe
9usgp3KF0k0apxzJq/ZSwdcVJxelAB6YbuhpDTAB6CJDHJgn8N1ovVSWd70jpi3gv5PZSCAuTm7j
Gl/GESCo4/ByE0BDRNH0gOr4h7HrPZyVd98nYeMQ4YRt2JutqjMk8fKjRvtOTuh4VTdfdhRiGl+J
xf4AEhpt3SsLWLGJFCAr5k7frKFWBXJIGbrPZ7+aAkixe7R23dW6ArqfBwrLxgo2UK9DeammtR6c
j4b13tgpqpWLT9VAGLpApt/oLSc/PtFd1H37Qmz9xY/LkEKJIChfCF9pKu9jQZgxGUL1MXiOGfBq
m1MCVczz/igtpLnohBSoW+F3YAZuqyjdmefg2CiZUWX938sRjwrk/WMJ9u2yjrj2PrLQ+VjpfHqq
WfLYkClzNzJYKZjHmGjjtvDRtEDfQhafecufod1iU6J+Vk7kI2sT5cyDxa0bZoDD1DvzTlFJZpgm
JGvLl3RpaX35em9sGBY5AN+xjN9xjMAfsgDm+tAEqUw87H23J7V6ZNmvU11O4PxfwcAG6l0eVAtP
beJbBoE8qzNqg/UpY/yukvaMpwv2g3DEDWo0d/th2w0299KKE5Su7RAyu6s3qanJJ+vgfS5ZBDni
lFB+tLzhEnUIm+YiiWpdeGtaZfJWqlc4t/jCleSRc8DKCVXUHsHdZipNsgbgAAc/8uFYCwO/doxO
DvEQ9vO6L3sACVy090zcYIcgyu23Yna48Iw9LLvAnatDb1heoodobuhvvhSP+5r/aLxQ14YPzIl2
6d3bJzoqk1BVEy7uUQxHVE4yrwXkiilWu+3+68kpE/8ygbMXMOYE3z39WUIfH0CVux2qIZJm4ly7
5I6kDiODUHE8NP4thsOS3kSCL65aaw2Hd94xRZMOxW8US7akSRXZXSRpsSGG/2SSFil58jJ8vWsz
j8i/ywxiIQsKYU//lZql6rjD/0A2Jgt/YRgVarDYsQ0C1fdQRwEBozyowf7HNLmHB2YfMzDx+GAT
MphkNSC/TWg73lDh85ZdQXfP2zF5Ow79Ck+fT/LnC5kPgPSU8B4kTr3sx0sTgmEnjZI21S8Fupy4
zLePZR2rvO6FRxtW7dijSeIYQHULXxU0/CjhFBRyF2824Pf8KseQNq2LMKGytvTprus82qtXDnQR
XP8sX9BgR4j/vR+mJubRWTsUwI/4cEx25jhaO2FcPu3D8e15WezkVkytOr252wsODxqaaQb+5Cvc
+oi0VtNXA60XdUtcnhRx7KARtBQkb7bjn5EA8jdF70U3fkSGRs+VWQFsMIk6Ie8xjNJq7m9Ac+PK
3osGMCo4I25xjjIyYcnxF3c6xdM3lCuyDNJTG+tjlsRbu7WRxIuN2IM32uW8ZY3vZ2TvsnzDzCph
AE87ZGbNdC1SeocrlpTEuupaN+gg3YFABkC6iK1qFaDWLMjipPgr/U99+gMFlGxYq5E6MiA4s4yJ
gyEcB54GoZEc8WqYH8EhsTpedym+opJ0uh3Q6VhbClja9I4j1sNahijIRKevSsPFDnuqpjPh+Wh9
Jh2VDV55ChYbJc245qXwO1ps6QyJ9lQbD5bNX63UZdRk1C/aFZafqIu3DPae+Qk83FJ0Ga7qj1mp
Ru70vuY0lKTLzzp2h0H4sSo4WnclaaM+BCKCqsmQybOluwrsMcgSbCwpxJLJEPNg7I2JJogpRhx8
vrEB5hZwDXEmA9Cph/0LyfQ+BRaR3VlxnK+09IREa9rvUVCbGmSr6vEwZWF3H3DNp+Z+zSZ93n9h
P07HLI9sEC9gQ1M9pk7NfHznvFeUcNX+uvbU8Gfl935bXaBOHo2unOQXsOS54kY+hF1arY0nMiaw
Zu9GCFcdnzPzWJ4JwuBCJUTW1TpbXVEeqx0umEbgGrzmOM3HZ2n/pyPba6rSMK8QFptekIaRNzgE
ThoIEZLIYiROl7vy+Ir4pCdhSBh1yvsZ7lRNQysxzzjnYbLf5NfgDVPev/+t+l2b9XQQXRMwXteG
N4vKAkpiukmXJwwqSh1xMMbCyCeQ8of1ynAd1gtx1IzKHuCNHSKcAy5e1nDX+0EqtvM7hVfIC0HM
6stXESKy3EQnTk/ami8KTYHeM2IL3l3BsxYystIb6qalaHRxnq/TXpezkkSJmlHrZe02mHVX+bu9
yUDZzDs5ypUF5O/Wp0Dhmryj+Ak50ZD1+H0eHgVupLobh7IvNMmKkd5I9jyBzeG7PZV/RSx0gGe6
DG5ihoX32tV1B9eGJipd/wcxjCy15M4xkolbp4lrszU7QqF1SbOl0H8HDP7/vRSZM9W9so8bdHjf
xBmJZ4HxKjSkfAgGl5XTszqq+po39foiVURt2cgVHi3Bvb4fGddT/l3ljyJj8kIp/nIp+840ZiKJ
gh/+2cryAVEm0O0pTXQ0c3sLDFoCStSBpidd+9Iwhqk2KFfy4LVwGUSjJSS9yVL5IQoSyVETkceF
NT2a8aunVGHV0xc9ECL08fkJGO+iu7PgA5Vt8sL+AKLBvDbTUg0oyN1RxLPUhAYtPTprHppaXizG
Jq6YIyPQCzw0uPFto65WEAoKgBDSlAcBkshqKQ4dNoGWmwWgqzJ+YS5qvIEWWCoWfT/EuJMnk6Hw
toVRu7HN8GDjNYWmV/4CFewMom4HPuRHgzsX5RKok1WpR1McEHdOS/MRXnNosZLdteUPzz6jm+M0
qwXEx4fUf14pc2pkQP03N36khEilbY7h6CHf5O+tkwXWV/Sawgc+SbCe21j1K+Pl33D6gKSP2gJW
yFLQuR2VVbe6ebaVw20S7+dq6HnQQjGvpOyy3W8Et09jWfjvbXux6C+Tc5Yeze8WjlXDKA8tSgMo
tAf0I2e7y8kkH2JDNQRbufpyuB9vsLQryyQz/p6zEklCrEGVlNmUILBI2SWbdvsOqyOxEKcLSfBP
bF9hN5qKxdZinPvb8iCwwJZ4sh3F7KoZvddGdQpCYwY9I4yvn4SVomnfbWV8e6XqH6PP68jH0DzB
3Y0stYIzVjHTw3xiHBBBOh34rkRUyBrLVYZa0X3yCeKf3tB3VFkKmQJMBSqbuO6x2P6qp2RqG8aP
p0hp6booMmBOAwtf2YgTJYKRByDl+ZFUytvsuk9/nor+5Z0I4Yw8aIlgWFNHSFRkmg9yU4LX5vK7
wc5ziZ6EjBwSNzPyflEJOXbEuHP0rwpGtzMrOhMntIey9jZJGl5dFl0jVl47gnPHdkYf1TDysO6J
b6nLK0ricOLoDr3dqBrZ0qVxegbjlRoDWQxqlcwW1BgXBaJHgLJsZDLgvo1IOZ9L0vQ/BAS02c0P
66EWqAIq/EieL0mqKJgH+it7qKATmMlAxRkbJEaOlHsHhG+aFxeFNBRojMe9QMyXsksaa6GNW6qH
4ewsVAt/s59wy8DX0iXJ6o2Gd4naa/wIbtn6t4FDKUCf7PwGryLoqsZ6UmG5truEXzCfGeY06kvp
wqIna5yTQAE/XbPnWji2PdMWiSGW6MOLVY/ELH4B/bzEV1t8iW0KduAJUyPmA6BirzhulEFjB3Be
U4UXlQW8vJduF/UaL3bk/nKRsQwJmQLFc990xQK62nnTEPgGb86m1lzfGrqEghtLJK79B1pZN6Ms
bc5EiLzfpfVRkHpJq/HjKQsBJdrpe4qon8832vcnyAp/dVdRcGdaztUiESNepM3qH/PlVjAHyI95
g0d5uCGrgv9/IvobvAwDXp3/EWvfnvmwlXcgEF/04NkCZnWN77QbWJq1yW2CrNVqTjkcU7BxPekp
GmWdj4c0VcxXBceVwY5RYtVvW3Dc9mg4Z2FBxF+PPj6YjHB42zIRi9BQVjQnjZ5tnxCPLZi9JdeQ
ndnRA04s4Y6elTjmEn3kyM5wnx6dYeRzrJZdrOxihfvbZJY2A8Xat7CQrlbQSLxpKVerhrPQ6Lgk
W3QoZs6cbKMhdS+EEjAJIyj2GDrnIXLp33b0o9f6OLFC+6xzvbMbLRnq/xcdJlOM4MFSnFRsPZq6
UjB33e+AiIhVi3dfkRSuY84ld1BCEZ7EawqxUI7536IZTm7DBsAvvkNZaZv5CtgxYn/ZZzLsxjRZ
FPtWiQg//oOjBWCtbmg1Mtn4i7GXdel8GAf1TF6QsHRBqQRrURRf8xeZd0vMmrCsmuJoH5jjCJQ4
eRyjUjT5mVZM/aX+2LBsSYLfbIyxBy0jDgFby9u4+/nZd7BqwAEuYfMzwP8fj40QuF7wLIdAWZpR
MqJhImrikVRw/wAFGX2B88yjPlGGaUi66/TfmRb8lPA+oT9yFGEV6RT2aDBtVLG5d37B1NmD14NT
Cmai6tTcIHqvMJmlBFYcV2cifIZeoZyPx/0fP5SAfS5W3+jBtmV3+5VbYlobiuu+WtqIz0/YatD8
8zOUoijrkKQwfZ78aSsZrgaqTY2ifPGp1JEXlMw7OR3Dy9bHVxqKiKRGcH32dyJiJBel1lxcN52h
G1mo4kmO/Ewiue8BaLz/a7GX5LdrIw4l1dJIaDN2NQLEAnCXc6MR+sBZqZvEnQp/LrXbqsAXwcCs
fSQ6S/81QU2GIrHZVtvYJFTmKN92+cv8OP4xB57cd4oygvGMGiOI240UnTkYgXs0757CEoe3ongu
xzTGnOp5y029M6nYD/I5aPWbjGpi5jv1KdvYHm7GcX5GSYB30DV5jcyQeVHV4oyv55L+27EEYl0S
bWBkNDKqkc2s1CAnJ3n9JSUppwryDz9LD5eM8RQUVJ/UTfSWmNLbPmRLf5U2gIgL+PqpaMkfBReH
ub6mbIZZ5xxUd8gTBVpE9grEy3tY05EXx+NkVl12jhVskj2brOjWcai0y+CmIQrCamPxXiRa5kc0
K7Tff85LSCgm/mSC1TcueSSsQMCRIaBLkf2NLjX81GgAIe8uZNAmtH4DrV8kdtP/80I25d2XRFUH
G9stRiodnz6f9H7VBF+1A2+ivrfomIyX+FgRCc9QHYWNQVOylW0vJ4wzvWg89eAPtheSJIHW7uef
MT5DOZn7Ik2r9xxzIn46LR0iIdPGvpR1e5XsElBnSRW8UojD11G1x2wSa+X0QKvGWByeEM3HMJ7L
epl0HvoTLvK6zlvMeHToj8zAmcyFla3rdWGIVhcSL8b5bEWXWdFbOSc8GItmZlbOUpTMjFo8lFAR
8VEBkRwxq/QdxsOEiEMwdjfQmKj7s/8xmCq7i6wV54Yvej+/qbEx6+UMIxATVAL/crg8p2Uc7das
oUxOvJ79gImVTerdZTunpNTpYlfAbN+esWcywirFwwURiqImblXy1r76xxTiZ5PjndqaV6ydFyGJ
6n92XIYsCfWu2dcFCRTb5/esqKwCpzgsjjQstpSNK2B7Bd/fN/XnyRE+JNhF4MIOgOD1ewHCqvTh
XVFj5j7CvsTAmBbb91x67DI6mhhUpm/ZzKQebHdxporUjJZPk6qIT3mR57e3eE2dFrOA/Hbn4mTV
CJxgRqNbj5JPG4t2Ytg2RqE84R2oDtYhBVB3ZToYFL4A19kH9hHQ9Y6lDtP6gnbbjnn0AMHSYW5M
7L+RvfKX9qVdOoTOcXdU98r4OhxbghVW4CDcluDNoELMX84ZTV0Q84Ua/4WCM/mPKypwP9WCzeUY
RWFuvPb9Iu2Dqe92epzdGp7ZcitKduOi5aqF90ybvoVwEEpRKBypGtMr/rteuof/aDjJkN81OjHY
mCmvWC+vOJko6wSiHp0ZFjDNZyqDvvycoskU05u17RQrMDl0S45qEiCkU6lgTPL9R/dfmcFQv1sD
814O5KyXzjJPYjHAw0j2XDxK7N80UsWzkizX+MMYMQD6ABFYA1ZEKLN/lFcL4UYwlpr+QGn5Nqh+
wGpwa/9+xYCvv2n0VJSjH7i22ae808Xr6CMtZeagwkVv8iU7KE8+lmtJ/BowBuG/pnLvr16qAhE8
917RItxDsqG2/eW0yYpCgxttu39QdM+nKo8u51qxaRufo1QA/0taYMr6eI9eS5P+TwElnwjThe5J
po0L4tt3tlguROnphH9zdxximaC1/r6zk7d6ulBTTp/I9e0SRxFyV3GoOYoYzYGEEKK9YMqSkTCq
K22XqBb9ifmCKIuzCYkMdsMa8W7WsjcxX/V0eeFtjnpenovIkmhxfWv2qKBinRaMFt5pV5NWtGXW
9pZ2sO0bPWCsmbebEPHcQZeFTBeDkrME3+NWYb/GgsBqkdUiPS8h30xnhT5T/NfWlY+A/5zPFVKY
IbPkcc5zYnoFOIVAb6+ipySlguTGXCl7Yb3EakZZ4jbRS6uARIi5HQPRwAEYwGy/DCmOZcSa87pt
ROHjbi5JUZ1DTsBaYrrE9FJT3NlgoO3KlhhprRrbdHvfU3zvXsp6Y4cISm8OQacIDVvo7nJizVPs
kdtcWwNzd1y5WUn1ckWMDkpuDRvzYsCAGn15dcT7Kk300yWWpztzjq5dTNKaQGftDftZwxN+S6kw
eHA9BmAW3NLbsJPW+ZNqtQxfyvxvjsJoQ4LOF6/eelVsxnEbaUM9zing0Hi48bxTQKbICT0SNo78
JINK8JGmGesLhAhLlUglJInb/im3gvzU53NRILVC63UI0WYbexDyXjkndDtmsh1nAdBr2CthuDsK
AI0WwWarF31zyL8qfSrDso/0RV1i37RWRcmSeOtqIR2rKOFdZVQYW9YZvOWVS73dfrhhZka9t/Yl
aEdBtSkEBa3hGhCE7O2Ue5eBeaswesMNfxQ6LN10vnncBRlaB8+2L1xut6zO1K9tgw9PrxIGeT4D
3XJ3v3a682udg6n3tHayShLFE5PCO/085dwEjrZ+4gSWd9Znj2AB3xkZc6QiE+xDsBiWFK/fDrSK
VXsDjPvGmiNgYRYldbks3IyJ0at/5cR2ssJDgCuIUfVPXj6GnjawO6Z1USHvu3+f8M7ILZVLoQzm
+fxtnooWkNaCIHn8eRs8P+zXLOfmw9c2KnVhcVYFNte74ccPMce69eiPwyGMTAGTs7uTMMQAsY5p
IDJ6rxHIfDlvP2UzfYQaWEFSHYmfhpzRUc3fU7rB4DxMHgsZdqGsiWfh8nZsk+e+3PIglgLfKcjU
5xMO97UDk/FpIF2240wuFaoJ+NBjSplaHZ2TlA82Pmlj8c5EnpcS4/W/BFBeceY1ueIDGfApxvWv
2tBVBSXBAhNO1LFg8MjY7S5l0AGrZoG//YtMwRin0x0jI9lBIgfGXhihMYKHSI7MZofTwFTsOZE/
iDkWZqlVq/yDWPCMBQraB+L5HFC7A/9veIfOqddVdxR5x6+hW30Zh05HcH7UJFb6hVe2/7sY274G
BtrpVUiNzz6r+6ehMbQ2qWb23W1AvmG57B3nDmTnGGgyAYaHm+9XB60XskMkjgYyVdB1pZVF1AgX
BZwKTrS1cxG1sa2P91jIHJJ05Ckd5vU58b1w16Urto9GPUN7Kzwn6yAPnfem9zKEQgG3ut9vFAWi
b5/+o7eg9Szx9aWYjQbNK8kh/3Qxm3I/P8hhEvCijMMiKPm+kvEjhY0lQPyndxQBRbj+vgobALS4
8DgVe7Oz2CzOddUuX6WE3USM515aL2giQPTdXi/xMbPNDLYOly4lkW+10/X/ovCSQAQrAygLPTF0
jGGklxG1F/6UUt5Sir2Wipw9bhtSxOwbPEzJwEAq0I/Ugc54eZR5c6j4kUf7+lg0sexGE1AkSq0h
gMbHIuVkWLYd0CUua85ANEIYkZnPumXVBMtr48We3vlU6Ft8b/GoBSupfI/FVU/7tpVXEE1Qw/jP
CVoqxpQp4+yvF61EUSbPnV9nG5YMcN63RiqTWSSiMrpzvQuCMwr0XzTBTHuP6ZDExD2g1wfzUfpW
EvEhTgCr+NzZHCi1qW7CGEmGZpG7TJyysUnrddOkdBA1uGPAfG7/eXBOcyFNnbJbiPWyBMQpPhAW
IGjpc9WmGJSow5oYyomIasZiKuHcvNf1AwhKrMNz/2ON2kLMxUM8gKzAY4dNp3E3vekUC7aJWY3x
oElL/OjDFnpU+6S3lFWybsbB64s5I4joVX3qeAXDS9hvDyEwjMqDVMs2xFKhiCFODR3QQiOPdMEM
FQL6jjgCShIx+uywpoHfcVcmuAzYqDlb3q+xPHaVuM8HOqSikRVxO4aSUWCpCel3zx6nlCGBvQ1f
uH4STTZeEYJ35dFbNk3Y0qzEwFg2DWfeDUBfSxxjjjZiGXP9x85NgYQndMvjd/4dHongbVXD8IM+
lr47S8hgzf9QGHb+4yrGlg2Z5mtRFi4yjtDavDObHTCuuQ0bNJK7k/wwMKW44b9rM1eCl71kZjuE
hAfzufSqVgVcxKvbxvX6gt41nqIL61y6qIotyfgqQxe7VSaVkJqf1DiWj38bIt85s/bEiosIHsnW
zy5qS7UZ0yBcj8iCDj6gkjTzFlqd4O6BgUv0cbumPCz3Cne8bbClDN6fQQdE01xXkRhrfKR4GZd3
X1nRtuCgK/mWX704HjHSK6pWoXMIkaZWeOGJevMhcBY3S9ON7Xjv/l6o8o902O5QAo87ltJy06Ek
iAQ1dWYMq4vTwhklgVpfwgNlhFi3hze2xikPmWgyMOw4HbHWQUbSyz0ZJ/C7DXyXCaU5FsY2gDvo
f0/56bxclXboDUaitNb2Syu+40/+x0Pp84eUOTtuMjIdt1axcXwLEporQrnIVyCdwmhDAiF2l9WA
sruwl0sKYkikKB3UMxOCb87RDTE6D2aNw8ITvnWgBQJ1oi+yAt5mdUz2EE9AWx/O5Bbs4zOTayfP
6TshianXSCl2GUVdEyz61qlA0w9o04GrKKaXlDeQTb1tWf7tHdXdbfeGiaWlD9zBl9QPEZjhVIh2
fdMB3gOnUaknVtxi41+QVlywbbUauYxqMZ1603jHFxjCVtY0Y7aViLEWhljNvojqe6yrqA1NqmB/
0xnSsPsgfzkYRPp1UVxhQtaehll7fCQMeS8RYnIHem7/obeVEl4CfqMN+ubTa8P7PwW+ZozmkL5W
YzgTYx/z3I2ge6jEvwwxo6PGbv/bUUhlgOdpB3eH/eKBYJUJEv/QOrz2JLcJ0qkJMttlErGW4ej9
Oc28Qalo4u6oncH+nbJLRqf9jNqQ9hS6gHywF2u/+OPXt6wLcyTAF5gB/gxoPTTFk2JaqYfSJbp9
G7t9nQ0pkip21Zbu++Ze6olRfNHUUeT/qa4eikGMnvQY1eX11Vb1tMd90zvfqNgt7I6DF7+vV3vx
MqiDkJ7HzPAIJ9srvBzAl6igHT3v+TN3VG7tSQqFlO90vlAYOEvQEMiE05Wxig66UnYqWRgilnA/
UWDI3v0qTGSCg28KG+gjrL7uuSGjOfzZZfx9V2gr95vlQ+yK/xeRVyiV55OFrs4M+sOaNNp+euna
TyegJhmfgJsH2nB3Ufooz1Vd6avv8hMPJTwTLCpdAFNE8L/kSY1jNWAX0CJYXkkjZ9KoFKZwIgv4
ueGiYrZl08+KuilbprHr8ys0G0OVuKub6JEl59ehzu65JJDyUQHzRVvU9km33qm27EBUgYTnO7q5
7rxGPtYqxfgcsVMMf4mfHk9CroGz9cnbttjwDLoFv/sjVl/LMbMVtqEfIUDpVns2TNebIYCjPjOU
q7kXpNBmN0zd6teIObpxuz4CHDLJcevXz3Aa4xHkTjXgu0spBhFNtvztapXRUqnR1zo8dMGJqVhT
znDkm84AWWRgraytMoLIEsC2zp6HYUgabD+s8cUERUKUqsSHSmQQUwuJOP9wCNVk29McWy/2tvN9
1ApylbnwX+yHVCvvRKteo8p+OAg/pCj95HH01o0aOndTVLB1gSsC7m9EnnW9ghxNI0mcPX69T7/F
SEmnkdibugncORPMPLaKAl46anrTtkRYkqP9HtvBqAEYoKZovUTOMRAPpc0JVN4Y+D+gOuoSnjLP
D4RL3m0yB+Ts1xDvlzVy10E55vHw/FZAdy1FbzoM1chiKXl+/1m/MkxgLu7fO0vZUb/h9OHSYYtG
/tKPzkeaWEAxX2O06K7Ywnwxn6IUU3i2r6ino5OzTGMti/jJ+YCpdiaLcJU+Hias9OxDD3fBVeOv
3KPY5bKp0KSGJDrLto1TEVmaPVYbFBhexqW/Z7MXWiebcvl+WWndIbjVFS8H0/1Ya75yLqFWf663
Ex8v9GaQ6hScb9YyBlXBNoSnqU0MrP4gUspdblt8CNdwV+6zxWsj77QqGYMmrOvIR/kHrEO1t8AU
lrsRKhJru+s1nziU9ur17saqi328YxS1FH2E/+PKKJhsYPXdC54Lhi+jQfp+xo72Ur7+3mkpPzG1
QZXB0s2433XRs5k9BpHPZO0SirTKwyetbS8hc+uvmRsisbdtTl9Q+nd7BL3Zk4e92OPovYr07cJO
OX3cLhKwWwdOlJ+B0I5jQEd0kLeILlUfqKcw+kSHc/yaWqgh3w2mnxXOvyz6aSGQR+4sjitVS3zf
fj2CgfFo5k9OcwAGlAqYTp95hGx7P+7hOz9SwI84J3aE23b9a4Xuq4cZKUVhHzgweb5S1yLh5VGV
1RQpfLjt10azX2WztthzS1bu9iFpv9t1cbxT6v/n8KanmQs2SoH/7o0dqkxmHpeYqZ6UrsscsevD
mhLIJZAftZtOkrr7cJx2FIs3AxPLQ8zREjPqvmZHX7Y0A9rG4usXtax67Dd9CS85MjWbIYjFurhZ
0e+Plk7uwMcAo81AEgEd35nPyxD4ceAJBqPgzmgNbS1i/u/m1gcJcCZ+cTgf/Km/QBFYfmYXgo9g
a7Sw/olF+nb8blXVOPw6VHgunTjjiAUE8XWwnAGBdKwukzTiLGst1tzg6lKo/Du3bRdZbct0cOOE
fNwwWe4RGkHfBoTCctA4Di7E+kPRgQSMtH6US+uQnkn7aXQzZ/YrBZ4w+03FZfL/S3wXKwEhfEYu
88qOgUKFxLj5Ut0yB9tYZ4RF75Xgj59x88YNe0hcjbH5tbQDLjP6hVxvkBYIoa8A0SMlmTYXfsPx
1BiGoZsGXJgGSfKeV/f7eOWltRTcYoW7PuTn+TLJFtMa39yF0QDLUdvKtpOLNKoEredsEL9kqFmC
2RUUkuuqyYuSAA+XPcs6PiasXa78fVmvjQI5BH+2azYdXLhu+BBNWWhjw4WHdwt0GTxZhUcae5bH
JgNS8hvSzikW7T9FuLVmwd26THCmldnJG3sL39KsgF2dklXGDbmLtMh0kPLdPh/TDY1KhFFiNdIx
Ogozs1UBNXc5hkhuzkb5WPNe41G2JqKZ/MyTT32M/eF/EyioA8/4SrDkinNv/+iY8TRpJCiVEhG7
K9Y1UaG41fqrhHOC++yfYyiKoYkxlbz18ZyNz3xKZGJ9jMfnk4f6kc1EWshmm+sq+jzKLTfTMoyD
/7U7xyKuuD7iBYMvwpe2+RtByIOSYWcg5WL5xkSsNMXQQH/l3LgmRr2pDWhCKFipEyNC1l7BMulp
y5HJlN/oV+VZ05ugnUGY4D44TJsQMIuyUNd6kmfElY5WRF9AtqNNpHjY0h2N3mPp9Tv4ng/rc4eB
YVuwlW5az8KWZaEzjCxXTmxBFwFzJjJCbzEqfDgOHvEnXjLhciPZOvibEqLG92k49Y1Rj80We5je
+hlHUK94EUIs6tIhKQL2yZViyX0y0VanYIvuPc7j4tGOvwWeMjB3syxwhCPTIApHHcIahW88yHz/
s4u8bbFSVUEOi4ISI5pKIozrMg0kdl0G1ERrqbJmNKDjo3oxkEoCLYE0G3BpqLVTWyiXA+Dy4IKn
4ks/rq2An1sCxMPz120TEhDE8lSAZlutT+UuL1NoiSWOuuEpKW2B9eheWHwkTDGcr5SQJ6Bx6OP/
1wRV9BpkE2tPjX63o3io2+qlFR00m6hBILjpee9wfZJf30QWFUxT+gCvRsfyHSLjn7wIioUbi65i
YUvtwW0s0Te6V7bxsazyVnf8Nqtses2RuVps2SpVLOMl8cB+wsf5RyrnMWsaoymVtdWLObItBUdZ
Kyk32M3bBxTiHdDwYUS+za3I+CsRDNWthEgMdXwS2unU9oHMUzMwGafcKSGCEtgNt3tOzV33vPgm
bjs+NC7UBNOexm6OqBquPW1MpD0ITkNb4la0xC9Uc62XWp1HrJnoHC7ZkF/lo6UTYhX3Ag0NBSlT
l/NewPaNSXUTAWxK5xxzBx68p4j01e8aiBFeURH0Ql7MePd5HwzJ5yJsy8L/QPqXFBUvb2cYwIOh
bpurm6HBydhYk1FtzYEu0+etdoydGvFdtruvH50//pXpogsfco5Lv9U6gmllrwt6qettM4vTNCcz
lXWzq1R2hT99/QiWRpmb+3DKgmNk5/ZCy1145ZLR/bFNs9uNMT0iZsKrdR/IqOt5REPNW+uPV9ut
Jl7epMCZQ62bBF0QNJVcaUV5tSde2pkwouRmhuIxTonkwZeT08ijgx92x7lCCHCQGEObBBAaAjFF
GwHDlHdFvecuJ18MAC8XgEw2qflyZbnuCmd1DgjYAQniBIOSYZIyNtziTCt2SKOh12SgR98TlnM4
l8CS76gNglhFYkBGlz/xGQbnC3+Bm1S5U6CbdtdXFxHNvF+841tKWBpBA2ky9fq7PP+KKxOduCCD
8AfPclRDSFtxMmPqJN6x8jzCHfCMbsxUagje0v2RXkmVPdIEKxPJdgjWpBzL24sOpExQUCAd9ndo
R43ldCZUMq0gmYVWlL+ckTOqnhbETWaLyeCBwDXEbIcFnUy0IkVGVy8Vp/4F3ceet6SMJlu4gJHk
W9LQeu3urV8ehtjKzaXlYInAnKgbrwtWfolTo1iHHhFwz/QvbqZxNvOwZnBn91niBvLohTwsCR+v
Ps3bYAOc6AA8xaWeG48zmE/CkVadF76XuztC1qYHl51INGbHaL3LtYNjG4ryYeWds1CybTP0NDJ2
xK+W20YJK2/BrT9Wo0VDih0k+0biyNAKHw8bgTdd2SG6o8aoSfYrd1jY34E9FtKBzirtNwL8jSEA
0/ZORWzbKQ2MTg/dyutDTBpCT0UFDfosvltwJhvcFfeid9OFS3UCEIyTSVb3mSYp467BgpDTvcXd
fPHGBt7yzOahV0tbXnaNArpYLlvUT4hCX0w9aI5IGdmc0PSySseWI+jaS3rmz+ZtdtBBMrTf+laV
RXrQHXCFPpwjzq1qCov0N9O0c6pUf883YPz6MgLqVAQ5zF+gw8muWmB4X1oX4IIoZM/3+SW6VzvO
jwZxZT+VcWC7a293gi0xCoNkG3WRFmHWypVV07IzCTgqqWI4sf0Ozc/gewfSo0qRPtVu8eGz5ZDW
r7Pvt0/1QKXqnihFlwH+3IkgChWZuoAiEO42wBgpanXvya9MQvGcXtpoyL8Sr9WY2rlCOijHogB1
3ACV0DyD9rMGigv6U5SVm+K1aiHT1fVETi3qC0TajpKdL3droTVAXO56AX9nKOC8/USMYtjlpg8E
5SexQgGtV2pfrl2v+sgnCOpuEZoEdhRI8s5oOneiKgETY51w+d1vR7FlY3vjzZEOlOwSU4bTC2pL
KbMaLk5yDnOcWy/OV2stQa9nlhcZF1A+8fX+ld0jA+cbAWX4Z4HnPOYGXAvzJXej1LmTsLZ76l90
EvwBo8JbMjXW4BQur/zI/s4NptejD9RaEK0jV4iPSBZ22SHcIbHnwnx94uhGb7wrYNpkQlCd9MVd
tZhtaRoufnByQDi+FDpAZdPfAnWp3Tlw8RLptBCEV3pHlpegqnY07yWV0RCGOZ4ccrhxLB8s2aCD
VxP7y7q9slEOn2Ne/ZKjg1gxtQ3a9rgLAAg2EDpPxSWDK/vQJbkUEJUosAQzie5Lc/J7XCtUNHX0
maB9yssxNqecVxDnJ/WaQN4sCBLU6VkXYxshQD5p7cM/ugvI1u9mdH/oNBu6cSLTRFgjHBCD0C2i
cO71UFBklPOsSDS07PcggkQ2vtsv6gqY0xZsW3rvWCRCh/TZ2TKUrmqYbbrIVfByhF9pzrsw8pp1
QUQkjvwDktXoT4Fiw01cJnTv1QQwe/Ol4wl71BI9zsIqYglqYDYfvW88RoSI9ItUqYMKzyyVGbsU
PQEfzkZ9fPf57iE/CLTBw0XIME7mbZar/JgjsBPoccxvawJZhoavkykVL6oIXL9moNG3nc1ikiLD
RfGfH7V0BxeKZ5VCws96XswdRcvPIX7NJ0vcwVEhjUSSvUIvZQUPb02PyTp0j4EPJQ4N6+ucnLmk
zsW6DoadeTKksinsqB5tKTjRl+L5yxFb5ROmKDc/YBYwnIyF1/V59t1kY6o3zGNWRQgCUns4WX2M
nTq2+m60zb09SWMlT2SPw3QG1nJBabHd+RALob8VxAao47ZGuUayJEDCN4oeqTMfGS8C9inxEAK/
bZZjeDa2XDHX3rVi+6+QmgUEDe/CgUy+GQhEFNDiDJSTh1CCPkhBhOtz+aGzj7gwI8QaTX3tHF8X
pcv0XWkW0ca8zATMpLYHVg8DZ6qLYX7PmOILza8xYWG8ZIu+EEhtJpcFdGkh5ZDPD++I55xsJ7Ny
fvdUxynL+e4cmEjmbHUwytGG2g+4IFR8u9bVfHyHn07TX7l0Dva55kwP6kO049T6Q41ZdUWTxYeF
hVAIeNZm82QbN7buqeOq7pBmzRiivSOswtzRJup/zQaFIikHNzu3ilXrgPBAIy9eX/hywrZQkfKg
R3uYCttfFNpcfHGBL9dGkh+WClTg1NG/N8h+lNeKwDOglB5oTQJocq58oNsGt+pFIkDH2NSTAOzy
AJybfLUOdqfrXrGuaGJyIzMqknEx7HVKvVqhnsvpBIl72F1wzlx11vPqSqAozpGoNggYXNPoxy0l
d+8S1dnwqzHkpc5DhmwXPE1iXUPvD8fs+/lyvkCxo79ZGZsscX5806bEC2hWayPukpLnTOa2vTV1
5rXBgrA/mZHiZKrLTXyBw69IAe+FK1TiD37W6Vj/HCWMCVt2AXe4qc0lYI4WtS0AWEmZ9qUuxmLb
pzEvXYj7C/7RGC0Kw02Wnqk4vcq226S7bFTpcDru0kNfi3+7dEmtRG6KEhKbdS4lHeB9UoXdZAVz
HfRHnFbOzLmjA9MpUUz0NajihBsC/yOZvRZAmZJ6QsGg118BiccLtjtvH5M8sHOiCCqAlUez6I7T
LK7MpxOvP6IbdDPu2Rk6O6nD8oVqnuNh/6ijBZijJi7AP5HXFMotiPK2a/AMby9XG32Rnb8qJKq4
1IwCVAfugvoBjVMuqwf75ky/BqUjatgkZsRoWGOLSyMI/bsgex7HMoyB2tovEORJMvODnejSi8Sh
2qRSSyr/uruJTu6LHdWjnW+LhrDBMOAkbseDw0UEr6fkwe2601V56eUEf39EcHDDuaq/LR5pGdan
ahe3Zl5Eri7IbzM+9Rf6PYFRQyOl1zkLOPY1XsEUYkuN7OwHo/2/lUBIaIKV9etvRwxWTcZTDkwa
XVqB84/G9WHhcNw7dBwuFESTHtdzz4NigzdX/+HWSoXsCECwBLq3flQVUw1LL8w+tpU3PsyKsMS0
FwdOFSVFf745yMdpP688obIoqQbaJ+6kOAP054jacslBxS08Ucn3hG4ye0V8AulxRsRez2Ne7Mhn
73JnEtCYShF38OJzny6rd9aSsRrf9eVN9BbFEHmT/cvoI3EQnlFLIL9j+QkKHCQPObXA5MJV/uD+
QsuVnFBqOGY9bYcOmkZg3qxYogv7AkRABe9MFZTYiZzxxreqOL4O8zqTT2Gt+2T5vFgT61Mv4J3L
S+tglLiYXWS8rH4XuD0DPa2M/C3QpE8UHkO4nsdDsytmr1/2A119RJiQTB8rI/TG04DsIcmKsGZm
dNNFGiU0xTNzWBfqOsWLogW3fukBomfHp7AF4IoUPgTKwGKDfIIuXrE0i+hdrzWAWZ8tybQL4GZK
PZpuGa8fg+jHOQdWITsiXif7hLcSrFc3ubLQe/P3lwvX9cnsZhCsnCjzJNOnKr8E6gbUOVK8KZ7R
s8+9Z2oOzwIDxB7W22uVSJqPNEKco/8ZrMNbJ5YdtNhW4YGKYK1pMPAiH6Puca2ewyAIrSDuGAgK
4+J3N8cIuu/EMah5vKNldsiXaEHDnXod0RsRftHJGIRW2q1/hWwcEldcL54eEaXX1Leise6rXYTq
hrOsaRh70rqrF+zMCNAyn7DmBWTqKrdA600JdAtohuZzds5eluKsaIWlkJke1TM+M0eMoetsGfGr
NCvnmBp6llvm7hMDnf/ENsXpq3LjNNipCNLDJf1XYvKRJ5w/WVxxRL/pujvhGiRFtHKIa4tpK1xz
+ppupe+bV1tv0VJCI4Kv5rqBGvdfec8WXj0WI8e9nuXc+A6x5wC8Y72AWkilpm6GPnUiF7n+6XYG
XpCTpx35LqvslgcmbDl59XuDC3LRmFw1QMMsXlQ/1iIzZnBKLVOwqez0s4sxzanxHmfA5F/alMMg
T1qhndGGMjxk3YVxMWxYYpTjh8Plncb6NYss/lJx8BsI87OJ/GnVEiHoGoSWS8fYHmWXZWXMvnYr
BOWI6hg+HxHhuIduUlt/J5vmdgJChdXOVBivd3n6d2vh6kyBnteWg5GriVi9iECQPBaRh0++qnbV
Ftbik24ibmYoUPiqfY/BwPoiHOYIMiW3rk8pFhi5w5ggpxe6C22uea8BgdbmCu0uuV1uRXbExNs6
FNMvZC3bYvDThDMHJGdJTACkaeBXbrD7DEEimDesrs1vloF3w+LXM5vB5EMXta8Vj/fpY3Pdyeuf
RWcdSZ0yCNVKMyfePi3w8Wv4KB6WDc60vpCC8nvDqDmObhouRvu9xBIVTy2E0eOEWMs7S5ZZtFHZ
zL0xsxLsW35HT4r8aqTXl84V5r/FVfxe5I2BRmpxovjUET3ijlcDcOdZgYb1ACmnjilOCa0AI+MM
kSjAtowEc5q2EV98dUkh00NF4FRD+EYzZ6AVrdUxhensPx2nzw7BRIILgoq9rrdK8aczrYAfUNTU
BF0b6W9cV8X2u/LC9jWkz+Vn4iSDdZ4Z1Vn0vt7AaG4oA7G01/XTUbwPPnzgFFP8jU60fKc6xoHr
mciiVxgYypjwPUyksFTZU+qp0hgVvcpb2fDw9FdPNIgIZBzgEfxrHTIP4CdE7BecQDW4izNzNOjl
Wplm5+FV4DyDGknevgTzj7elHKWaLU2YuBwYTlGJwO6wN/7eUP5ocYPwB4TxnEwTpX6ZFKDmLLET
G0yorUhZoEJKGaQL2QP4zj44KoMx9/MxKNqOVSxz73ignkjYovyO6DkGJOlWoSkk4CogA5BPM0mv
0dveAH+3+W905pmtuNrIChc9NSxUzETi0lsDP6YEe3mj0euAx5vh11aZZPzrEmy0ZLiI6mPYEB6p
c2KPLvCTOKSV7pDQymRRv3CbTjw1c6Z4WI38kabbyID3F7PgPDluFX/kf8KJqxdix8KBQWjHEqwK
F2eAvfV/yalvk9ZAz76vRof2XgFDBvJCQf2nXEoGijuAFb0zaLVi9FpVNP92AfpkWaFWbxfbEKLP
LsBudphH+nlFYGhhImsDxY70MRB0w274TCQjCZdZ9+tK5w2WKHV954tqweoatAFOMbFgWygbcw22
FKC27iWzdA5240YTtmFC5chhQTxSpuaCRPQsDifbzDzdgVAvSINTbLpUXdDIDZ51QWQ6sKr4H7W5
PFYr/7z4JAUugtajAdbipIOtVYZqUAaUJnH6pz76YRSmM+RpRZwR68sIAP1wNNldJ9yAY0qJwZPA
u7FaL6xrDxyF4meK20o10Q9jOEUfUl1AzmZ28qKpmblOIoJx8eUVijT1yK0KG0j5YdD/tc0azHeX
wlYJhDrx8rfcYaYu+1Af1MNX8byx2UNGYtTFtABGGX5TffFtzlFol+fRe2PQG1OdOUydaU2svp0X
ht2WCTHYI2i1uiBc9AqzPqSakSaZi0qcXad0EYkCskipfNk5am2hhj9dq8J3QZCEjBdhTnAJnvlM
bFfhSG/SLNhu5EQ7ZVJBiHcPZbMgkHJMJPHs2dVA98svXunJWCE2V8Kji2Tgi3WmYVpohJ2UyKX9
QLU1dUOoGP7UEOiECVZlvSYJVQxYt3yI5+zvqCFSPW/aJNGrq/81hhkJvhdPEepu2wnp1QpSnPAD
rNYehla5+XedhRKCb85Qsm9IpwyUtCyvfqpRF+4niVOZ2Ja+NXEId0GRzjZsTuyObjp7zo4IobVM
vYiygXHXoC6/zf8c1hdCXg6wXoZsD7OJELaNd1y4LKMs8BaS7Dmg8dTK+L9Dyf9d1ZADOWPLDp2i
eFInGg2DEArUExSSepHypf+dPbsWrxFuBbpYx8EaxkLUMk717t/1tR3qZDfeNpw80zCP8PWzZEzr
4ZGUCx/hmRK1F+Lu4twLbwa4hVOGO3No5xEuOBcR1q1Pl4bN8kficWXlEIrzrVN+/vTUdISX/MxO
/4GMT4PvArMqA+sH7bdPa5Gm+DH3qghbJ9oMwqlNJvnd93JDpSUFZMv5FWhFAgnKLEvzBl6+waKP
zhpD42jgiwz2NHMWgWBbUOscfwwBh+F6CSshGfZM03dJI6ZcVgABtvo+RYEjP89pzk+GuopNVEpN
x05zXFzUiX4f6j/FvTCT951waczXJCkehYYsGWe+7Hcwrwn+ZtSHlkieraaVMJzSekQ5WzJdZC2G
+BuHDA7cNr9X+wHgAcj8XAAcfRFfytwLILWmCyWA2OXIEuLmr5VxC1wD+u0X+Kw7yRYvj9jQ1mx2
UaTBUjEFfonaKuJlDTPvOBIbB4SF/6fBWmvz6bEQXwdIfnMZs9OJDmNrMracj99lXpr+ztudcGwV
M17afZlIuuopmtIVPloZt10HCVuMiIBk+VnqYst84Kr7Wd2PrhRFUWDqdkxBo+M3I4iahYgqTPoU
PopXn840gISA/iccHsuSS73nSrw8byVHK4VpHQZHX7KFhMvGmm3JbYzbxyMuNvr7SlReUnsfi7WR
ySq1mQbyAu+m3+rfCy8efjp2J2IdLENMlM2LcQdYW0c/JLd/dS/8XNEWDHFklNUovATBaseL+Q0C
jBnYWLcMvcq8msfY7y/p/zhDPo5CcNDC1uzCqqR4Bn7sJka0d7hsc2j9PJEv2ZCMYce1/kH6Yr76
Z3OgjW66nU0AE5d1ZAb5ulL/LmCI6BM9ejc78CRoFglvN5DwqTY3mFjhAUS622dvh7xPiTCzf4Ku
O351iXGZzlL0jg65wQm23zhnij3UQTnHbg+wZIHhyIxPjC9IfMO8IWblqXo57VBx3mRIaLYOLbJG
20tlNJdLXdRTp65R0by/3/4VqFcdyyzNaRW3c9saYc5dd/YWf24YcOqJ0DyKqlRq/47jrlHcK5/z
HqTQ8fmClf4QhYv9c8ujiNZBs3ZIxe3mqGMPTXsg74om92ctMkxj8VDxU8sw4FMDJNadorf9hInk
iAmFtTG5VlBCXXoY5SMwNW4RPFCb2iuRYJQwSCD4lkJCxiuUebZGn6toJ/BP1b1fE9Gx7O/AzIVc
0YBt62Hoc/cUYweaYmXtpT4UhmXr0leY8PYpqdBQ86BWz1Jc52gOUiAnhCX8mV11SwapX57UzxCr
al4v+JvDB1EljBecdBU1GtjFOEL0Q3vRFrVNtRh9x6ztcok3hpDHNcjhV7s3RHJ7mMRglRadXhPJ
Wx6kd7rDBzLptCG1apIp/Dj4stUbXouejnHG8AgyAmeXtFeXhwf7i0s9yCbs/SqZZrF1RRMReSBU
E0Wuj6NS9Y749rWT1q813JNiZahmIfrNjLYgkGGbl0e84eRZzjr4vHFzG4akSMhai3OyM3i5/rGh
F88muL/IT9cPZFdZJsTkeaAFHLjhP5a27jKhzE3BlsGbk7ZhStt8ouZG36f81HBjLNjbo1NTarCC
YxClo1cDV7vPSlAwoFEXg+Q3ohpFUnjVFnkXy6svrBMieT1atkmA2aRG/to3ZBarOaZMr7y6Fvl+
QmLZbjG7AOLs1lzfUFO/4Dhu3RSJ2IMozKg1hhTf9gD0mu3iRoNkMLR1xw/Dvo8pAKz3uToiQSPL
Iewma2GyPZh46of6zObHfSLnjnUQ8QJcnHAw1bF0ktQ96X0gtn9rAfKuX3Vb5o1kZ7+2x6zDDeGI
qgaq04kUgn+dgmd9ARd9ahza6wHPkDKywHU4OYNSImBOfpfmODTJ8771AClffMntXhMD5zGk8y3s
IEtz1Rtd32yTOQTN3g/6JDVt/qwO6J26oW9VdHRxwjancIY7fN88sH9UTwtGxG15fgfUBRqMLnPC
xxYI56PwFoT7kpa7CD4cJ8pzIH4c6fJTIlx6TjsUnY8QCViMUryaorDCEpIpqZxoHVOESEqwoAHo
uabjQosTxGWpoPx6BCp4/ICXcVPxAIoPFzWaZCyoqQQ+/yy5983otpI9HXbWq2sgg9EIV1EGCYZF
srZb5z5kN6rIqCCuNvtU8YHyIool2YMIBueaXTtDxGV4hilpIsIvEw84EhnBSnye1RKLXqHPlOdL
0l82b8v7aOiWmY5aiIsudBBkEQQaOBGUOmmsMfqB3iqO8roXVeuQR4VHgMVDpK3veEfn25dImOmV
GU41xDMZMQwNht0JP6SJBnfuoE9DQf9B9tjtNuVCfRuF/8dKQmA2/fviuI+IKgxp/lFVFhwcYeS+
L2bk8qmVBRZqzCBh7A+XRpqg6EFIJ13IQ9JQuVRYdgZNRSmkPkE9WVRbJZFpcUyIcSRR1kKI8QJJ
dinv3jGpMxX5x6c7kvHtalnlp8Bvrd0XGG1ioV6yP1P3nd70tmQlMX71o34T9waUMOVJWRvcqeTJ
WlFIJEBgLOQoqMrZwlKymL6vDkRbXI8GcQyJNhiPO8UhblQCy9VB1EOlW6GdOUp2ejUFf6OjDXIY
/NloA2JNywgXiazIF+rowYR0SBYxpx7sfusvo4R1L1uy73VLwFstwZT7bwpCsbnaJGHr84flFnog
sdAZAGXOfNtjvL4hF7ggLTIQJEkGA4Ka+TW3r8YCPsmWLlV9Qr1iBxA5R97Q9Ft/NDQDNN/+qZum
YXE+dX2SUl1SPq4tYR2uR1DxjZFgkKyV/biDEKBIegPfSdEWUIkxp8aE2YXm6r1vlBcfGjCSX9X5
+WMBrWlNMg6RGmIM/k6JMXOb7Z0T3yx1OSxvITEYAmFExf2Ot/WzBlbF1KQNi1ADAZB9EzjheCyc
39arqPzY/kFQtt20CoQscDijP2UjEqOdbLRFpDDM7DAsBqiMfoeKmYvsGkrb9XszoJ2aiDfzj3eG
Q9LA/qof2owo7PlM14v3GK91Xy7xvaEC+EHgzTZ3zC3jNDuvqhJX3UIs0MRAtBk5apfIBjj7IuXH
zizCxNveITEGUBdRMLAwL+I55l4b/V2Dn16bN32BMYLen5Xk9m1CoKgj1AiiE3qy2Hrwm4blNeis
RWMXlShc95IpM03IFVXgQzMK56c49QdjFibYKOmDDxqK0oJ4+z0MXbvmgrZjODEntjVHsI2vM3YC
cg9tYuJcXUxBeStdl6IgNNm2GBVNNi/Tv+U7PehuZ9CVd5Rcgn7wKK0meHkAqkUv07sxTqP/wx3k
Hiz+XCAC51Erj5jDW65zWlBymyj82gvIFHRsXV1QYB5oQSW/xdxfJKL+iVlJMX32oFoYPLFWfPmE
Hr4CWKVdz44kZYiRNElzQ9/Aesi6DDIySMMOoUrRDNJZTxqissIB/AG+n9hMcGynkNrDHD2ITzUX
Rn81lWVFNBMRb93C+Xi1l7HSSEOxX3JshQzw27SkBVcQTWrKJMLaO+TaEFddMM+EjkxQE9gbjWAs
rGje0w7z7KyOn0MEwt/AIu6PjkXZ0IFDTQCoNPpCXterUX1i+8cV2OhJJ7+FJIcNOwnhSBApUrtG
5DDagiidzQKbAloCZzCjfWwSpf7ItbdT16QdXYO5ZMFXFwriqfhouUSfHy99mVbGwd7fLkisXED8
YrRWqTgUJyUaQQA4nJv45EzN0gyfZo29QLGiGmkREHGx7XWgNy/PqksT+qYF5qzDvPcOOgYW829e
U+avyw2GQw+mzHVbIAV4wavbQKqgMihMxnu2AB7Cjm30QvGggu57Cup08t/2XV2SRo5ha/h++aQj
WpsvebGhFu7PKno65AHmvDZusSf22HUULNw7PNie9AQjGYkFw7E3GwPSHIV+oGsPFn0KRjryNVbN
jh0JDVHGaGIIolifDMhv+Td17rTQY+ont5RHYFbN0N7StafbicXYZxkqhPMYOcWzKpGVikhC8dGP
PLkGnqwhipJQvAo80124Lvhs8sdQbl0++jRF6fkb0CgZuXuQEgZX5otPPARJtZUg8DRI8p1MBLUR
yVF/tn41Izs5ytz8nbol2TudIAbNTXwJDAuKnhk5DUIRX/kjizLE9J77TX3TlvTEYxruHtpt8UoY
fj/oQavZogta4cTCiH3YHDrO00eaDNgJr88DvC1q3HlY3JNtEz7/Xey9taCibUk5rbiz4kRh05Tk
sNSj8rK505m6QsDtY7TELxuYvJrMFcOOxWdsjDiasfbz7UaaWZtbM/gJIcYR15Nz132uoDFAXXv9
2ct6ZnamaxebIVJJHoGnILe2EI3fL8F9giUdTsl24YoIvnr43zFR0pKLsq67L1wVHwE0a0yB7i8N
8amPm6BlSKctmMiJ9bIpDrGWycUqGzAV8K3IYfFFy2F0sGhRFgYy1pJE7poXa3afVN7AdIfqgs6h
3hvU3NU35mhptz5Cay9iyKHGaeWlFEXq/Wz5xSOPDgASMVIJ9Rr0GgK44mbyw6qnyhURAr9E5IF0
17qpLSwwlMNXfFfvbA2XscWA6JFnNsseiqYvMsWDBtO4hWqXPZfH4MnjS/uB969lNOHBilzKlPzF
j3RKSHv5LZeZpLHhq/I+YFD8hO+9KnGSVmiNVQttHvcv2R4fopk8SNLXKfYqkjwAn/j/OcM5y0yn
QAQx4r2DEaXfx2C8ohylmQLdoOe1KdYy+mOMOiQH3VQC9WTHAAUR/Xh5aUM2ZI4B02gLOFCCIL/J
uBES/LWqPpHaVj4yDlDqjGSlLwmyYQnADyWHkBVuy2vdK7tuvOlVwPVKvMBNfiyDHbTmKwib01Ws
b88BLETdpTB3eAHCjbkBEVFpLjUJi/LSd983KFYB4OMGWwio6n5W53dQPsA63kWC3eErfozo3IZ9
yd5MJJyBSVvJ+UtZiC8+uu65MXGN2VipRVohbRMzrIaO/+9qQ+PENa25x742STxJMtykjXQS0eQA
SZtVADPcT+GWYHUgdXg660ivLx84fOTS+qGCG0R9QTU+c5xCjvZabuThHjAKULUz2LaLGgph05Ge
g9RHPVJhtfgYchX8+2Fn7u6FI4U0idHtnYbXaWXTsFFb3sEbSy4o2DtQsvc7N6D/7bqh/m2hb+ka
jiPvIpvwQoJhQLs4ZSR1uN6eHT3XoO4TSmc96yuq4SdbPEI4LWgpetQk1/pOFpv0uSEF93c+zn5i
Awn588D/Y1qFC/CoIpLpIyqn00bultzTLkSTlRwaP8Au/AjrcVjE23/zcdiMrnwg8D+kuE0XvTaU
yoLiGVKbt10xfYCPb2Cl/D+TjFg2hxaiU561MPqhJor/k37CuywNGSycUpdKbQP90JJ4kKyQQRhH
qiTH06N62JIRHIW+KF6FtbBE7wJHHh00Orbn4x1wIyj9BDFYO7BKfthwsbooP5WoZMu9FEdVIKK+
U1QFN77LzNUdasOvPicAt+VPr2y6HTvrV/RaraSVR5jGp2VbyxNt3Xd+I2Ekrz7kGQfZzitMICzo
1g3zSjelYTH7+i33laslOIq0kyU5RLSQxBNDk96Lnq4PRzkHiXsabFXm8RvpPvmm+a+P/269o/I4
4KrhyQ+Jb7n5+dDJWbeibBrhSnBHr8tyzdTp9EYXgxUpL/NY6+b+Z5BjJidCjSuYsZHh+8/CZzoq
Acajs1n8Gk/WbhUR4u+uONr+Is+G0hvJTkuAUv3O1cg3DMFI5q4iQWXAaWFDfqOTntv0fCClJbkR
Jh6HgrzkaoZmrXStAmINRKenvV3byEkxsGh+ddOlJIG67KVxc2ZV10t7GZvdMtaRMYwWPH0KMmM+
htAE55kbhEhDlwTRs3/RNYdrqvYIe2pCM/eQ1W2w0wkyvwzMiFJNBWt1j4Qz2wvLP9Zgy6u/9LS5
PbxuD3qyOi/dYjH24XuDpCeQdvydLlBx0fEpHJF/iC+0SvGPTlmSKvbujb6+V78knV48QAKemymy
K6qPEkdxnLZ8JHNjCcVu+DsCEdA2buaTDUop6/4TRkbcCKMMKJ84ubVWhfr6LaHcVZ6qhVkwduTJ
+qjg8FhH9i5WEr83RfjQ78QzaLTZNxh0yQo2a4VDqk5ZimS9pOFvOY3nzn5UZ3RF47b5pVX+kamc
VKT9Z6bqC3NUyO/e8f9LXhzx0fmxwp4rN9IBUGSRyUixm2Tl2S/5o81NGiApGcZYeVVjviDDpe2+
h9B2+Vgny1wT/9Az7QhwakMwvR67HnJuK3H4Hh2ZDfO4DUq5BGBpahktN7oMefVzgI692FJMR4H6
2msEBt3O1A81fORHuMxcYvL1P/1itLr/e7OP8TiFqLSzbIzs1219C+U9UNx/tVNqlCenfwVUxtYA
rnNbegt+YNWKitVNHHzEqn/fJjyUFl5VjG8GbrhRKWKkFrY3+RZ9k0snbFfXfkDRj8AAXqV/X88+
Ssmkaa9BHoE8ggtmlh/X1IwxStWU6GvOtoKDTLCMT/NA5X4vRivdavApHt/ZQBp6A7XVH6GESw8F
dmX2ExstPmO3QHTqvrLTxnyu4q+hUffGWlhy84DO34zX+pnohJcbrhv5SuxImUDEpkY5NqZarmIP
i1QwVb5BZGpkWp7M7rkvYN2vikRFB5FiGkjT0n+iD/DUiGp0fBPq+BnqtBKg1e/HscN1FgFuTmoQ
s539mQ7B3KHRxTZSivjzjbzaTu1eMRww6bwGskOwcVzLymdlhLCVvq4Hsz0Y9p+r8qwTGirN6E+4
Zz+8U2DeVJAemmzXfvoWkPDnAXLuCRn3zlL9bXEFYs3lj5FbTsth/lkfUyNs4RUyaLuMja2JXf3j
L3+gn+tIiMPZpcKphqT50gHiF/mSc4HHyeafmSYh3R83A7aepn6ycNOe0fOemYXFeTE5tJNmzO5N
GL6MloDiPK1K/PeU/E7GY+U6Tc1UKbEa5YdebnaPHZeX9Jsqcju9m+uCLyUEuc+CiCSQQny7SDy2
7NdUec0QM/UzodFUltVv5hPq9z4g3xjH/8dxWKqdC0oKPk6NYzm3hnLpUOOlyk9Dxy1Ayi+EfPXQ
lAksapVXcygMevYUl7B9Vz61awCm0TZDLl/7u+rwTuAfwAzxT0VJyNgfepNCX5ukgL7ZyAtTPhk3
45Va5Aq7XYSdHG6h1SoJIfOk5nREUyDC4P2yI1ZEHLUL3vVca9MVOrAS/JH/aNAPiBXJgUk9a2bB
QKh5wkS+eZ4MrRlgAgJLfy6SeDhSHnuFUGPnrdtWkkLdCTKqfrJWoOmBcTRiAeISyIrym9aWKst8
7qNM+JcyDyuTh3yaxro5qD9GZtecMLNq4WO3+KuVBA7Op+2qEny/xb5uhk7OhDpsJG9aOtF6mX+i
wxAuSL6XsLLbZaIHgbPsGSy4TEgyxd6ldo/Uojp7S1StOiC52p9KM5QqRtXAGXlrMmdSvK6oA4cP
RVapTpYEAV0HmatAr3P/pru9NHNxhCvpwZ3RG2+zHYEQeYjiJkyWXzYVdFYVQfM2rHlyFD9nM+QV
sbcI4kuu4r18CpYy95jnxX5HbJIjTt3XfU6FmJGfoYPWtL3FjTCxqdHBRHQzAcB/3E5tmFMpetK7
lQOjTS5rNTvBJRA6zXupIwIgCRkUJgQvrHIaUTnXLdwz2TaLF1/r/pLg8hucJLzcu2FwDJhrAgoH
Gcw1rKfYnuiocbnT7/uhZuIRU0F63ImFfD08W75WDhZzbwndI+W9oi/NvzE6DGHYLazydMKJKGvB
vmKipjeG06ln7Zrafiv1eInNojWI5yISn3QRrTkWRgVxFD5hEFBLxInI8/lLxDRQy51tRqosOx+m
f9kTvLup88CBaT56nmbhGqtOZj3KS+T6l5+viKExcd63YcBodA+/BxwtamYEB3erJGlEUyVKW8bh
D7ev2rXh0bgqQnZhAnUvHq7/mcfZ9osbwTNjogMvsR0rmEdDYze1+KJcQU6qcd40HezIEVTHrBtg
fNDpTnf1ydcL6PxNX0ZupkE5W5FqovDL2/8bftuFXYv/s0s7D/cnmttZ8auWKYiHqOi5idsCzpvz
OSpwSobiYkOtVurQQATNtYkW1yOZZ/l6VSZyBWof/oWAqKeT8uXOcR+LiY6yeU/jsTr3i40FNtZb
GU2eUGeByjQmzvBUOtxH1HFQg2IwLh2KoUprfEJF7Cl8nHcDMzol1Fwrlqr05NPeMj3wSe3MKNwk
agiPMHdAKIpaJQPDL3F4Q22HN4NxHcADxv19kMayhjWV/QpGtOxH8hFrH1oGxfV0X8T0bUxviWU8
gPEU1LihzznkrvwhbzGlyI2cuXar7bFSuzK7xaeNDqA7kqIz32/u7t7XE8jBzBMHWC9X5XSgCEVu
a8WiJsFmWvQ3WZsyOon8MsQCNq/X3/jVifGf+M2uAB9+P++MjBSJpT+HkkpIzsRcKPScEr+9P7EJ
31Qwt/FXUH5nh+MNNzIvJ4TOscMpeyUTtWYxe3OhlABjxC0mUwa1GWcyfw44tNd/2ptzAltZzhYg
QMah0NgjhJ6IH34R7W5/5d9D7+wu1hv+7YuaEiYisCKMtKN53X4pK9qZT79epZUSe0ey3IzyvcMF
cqTF82hENkAZgb6WfUBPRviX1KKS7S7if7X4hrgAkxhKiaNK9Jv4VIdIXbJjuGyJwfJK9vUKeEoA
uk714lfMsbttj2fYIqk+/fGaVCqeNJt8TMnKbO9NDNE31WxG/6DqFa3C9EysOge/hJDq4pRm6WI3
HkHnIfW/d1I9F4zAVSLtP/vPmKfL6f2O15yG9XhG9+n/wZ2cJ+6JHXDm25uYMycd17ocCjeUfLIE
b56WuTEn01OTPLtLAEPTJLkXj5SA1LUJY0ZleJS0p6DmLSw1zOwG1A+jC0EiENlMzBkiHEBA6lq6
uGcIxRw2ltoRu76gyyAxhANA4/9WZIy12FNMhpyo4ifNsLOIL/Tub/r+1nnC8nuQJVUM9EHjmzDY
amvxsKUla56MfPl7q0BivxbKkasX0lVauL4UA4Tw4TtfJQ6zQVMM8IPlRpl+DpawfoSVP83A4Bt9
yS4y9NAB12hRNI/35HBm4Dax3BPE7/kxwYQJLMW2t/4eg/59FEgbhPwCK+bjliRuDbydb4tGpnR/
+FdqoZfB7uY9hRtzRGCI3XD2IhMeQf2cW5hNBsv59SWLiiPbYJMc/GFHQMLMH8wUzc5UGju/0y5v
UVVNP/AwV/xEbE08gqsufF3eUOWoIpBS9aOH954+KvxEhhbIR+rXZoXG8IZu2elsk7dF/OPVc/By
zmi0zkiuPJQavYJXogNgwluk57O6u0RBqzcCvZsTLjf8My/g/yQk7ChjYipdPDTsB5Og2c08iSCb
KtZDqWTUPByQUGY82wJxuFX/NbbrrE88lKuHFQJsfKlvm8O1miv5GtiCNS//Teuwq3Emzpfw2wEH
vLuKjKaVNPFf5AZN3Lm8NLxEtafN1vZKc9O8o8b816ULXbHAWrhJQfj+BYGcAe+n0BB/Gae6WD7j
WV2D6f/PYuaYKkvF4uaN1t5WRJIJwxzpLRajrPj21ymgr8bRtlD6anm3kAd/PdqXkK/aKtP3XfkV
5/3SxyIq5cglCs82/ZMlA+UA6aUDas/tjCHP+CWKnnecIC7gDm47BIXhdYK1zfO33aTk6KpeAolv
0ZpnUW18ZAM+q07+eTyKZxfbBC1ZfBVlWSUPX+5Q5m67eKE0FxdrWcy9/MtuItyUP+ZJKT2Be+V4
uIIfLotBuG+l+YKAB3roZfre1kmutHTfTlnGtzMNOyWPDrgs08YVrDPDZSM+V6c9/7WY8ENkyna1
Y/dElFzabLLe2p+4mbsDpUMLhauWQLTHaSngb272ZmFgClwiUW9SaHWB1AS/jxPW4AHBtCNSMVzH
QZuQJVeXVCRDc4dSjs7rgmpNx/jC3qqnBWuH84JrQe6M003V1vx1o+njtXuMNd7ADyrLy+A2w553
IEJKZNqt9BYi1cZqRAPTA5f0hi6Rv1YCtccSEryOY7ktOM6+3Udqu5wa6KbwwjCeSlOBcW4yONnv
sujSvQ4/QSs7k8A8Ei0JSCMYrDgmJZ8xCPLLwhoEaTIBOceepjkEQplMiABIN/LvSPqzb1La52Vh
AT2pNFb8aWJ6ZyvVTOjaesQ8xPnYdIqHWpYq5+bzY005+tAij8oki3omAgKv9mpkHFtT5dI8fl9G
A41EVu8dO8rlzbt/f9WdGxG+ncIJltGFcia1yR+meWKLCyr/57GEWnlnbCZzNlPunKREBn/sqPfW
KHk2RjFhXW9pb3FPWjb3tjx3pr+a94AthJc0Hs6EAI9NO+AGvx3J39nmOw/GMHdwONH8G6mIpNmJ
8AP4p5jQCK7Vyd1GBCuCKy4GSvrwwPTFD5UAEr5OaRADKmMq83tIJcqyxrucTuOb5oBhZ7A/c0xU
qnOvcxQEyiHWK/REj/MM90fF0TNf91/85bTEdV5e0ydiq4pHlUpQSY/p4w62IudUBT6SE9i199Kz
Z2qNC+Lfd9v2tlTHcXVX8bqOOITPOZ+CmqONZXZrM6FE1A36DkU6CbaibCvTDrFitT5gLoUiSLB9
ptW8bLMpWEsrjJK5E4ZuYqJzW7OzQtBcCZuhu0V//S2zvV6Em2wf9Wt+WkUjPkYq00+R9y/HOA5m
PNIX7V8HBJMFW6tnwt0qsTGgfn4rwWT8upiSOtqXuqhrRL3aMIFntidJA4nY2rU2uBXLuXvem5L8
Sk7QDTeNwN+5xFt4WPms0wXUQlsUFYe5lsqHAPEG9jGvrV6+cscoBYDsD6nHjg9F7n8c7/n8ZUFo
3ZeJjHII/M4gKYI9KxM2FBLkbKKO+CRMo4PK+hRr5pwzdBTF744QeMQCY9L6J+Xx84tL+sJpxRcV
s6zDKIs2E+VDhJoMOqZIIN3oi59XohKTFh1f0ABw0XsB6zGvIyyxjt5VAvsg9f5IdEVa7AQE/1Z1
Kg0hw/KE1w8DzPuxjY+ktcaDp+QRP4XBzuI1aZL3ICoja2wGqgz54BbFs/BjllLKB5+ld36+xgWL
aZ2J0dpldfhmtr5MqcRQILoXutuOqONL0e6MA3tf7y6f+EYqdQdf+iUZFjutcYYfKbT/nuYeQJ5T
LCimLfxfvPhRda5L9XvQwFqurSWo/eIE8aWq2eE4JF777+dffYNIu8/mCpF6NB56bUeEp75xdLdv
B5vKNgTwL4k90wr68SXPiHFGrIxbga52VKu8zxGG9I5QwcdQ5WLcCTzGB6U4Xoef6HByB+xQxnTp
ne2jljSbjVAqJPHazV4FiAYPIsqaeGRVp9Pb7kT6i0PsT9qaav+fKtb7avCCczm0XYz8fKgYCg1L
i6zfwgKPo5jZLb9e9UtiJPY+AUA9Gr7cDKhamufvQvKzT/eGwdnGyuAwynCx1oCihtDUIh2IaAzo
2/+3EbIeMHgISjbTgA5g2NuFBRrbCbD91ayrnbVKGQWXaDBb/XfzGXIO+aTR6bITS6iN/SZ2tuO6
RiY2crzaNt1zKUhSJkYfQuy6q75AkgddfalCvrmxkF1z295c8vYuOboq9XwQOdTejTFiNEbAHOqK
sre+RfP8FDXZ3Kbp/H7zOmV/msjA5NrQcOazJEhw/VVUyD38aIsgukIzWPoHIu0K+NR8iD0x5CTd
RvUnSfz6A+sJq+H9yaIUf7TkRn6J9go+Ojk54KeS4+8HSGi1xRCSc69mH1Ga0qtNMe5ULjncfc+Y
R6bS8LvOVgETKPu4QB2QuCOUXvwCdfUjhe17nxXmzmdw8Z3sqLdF7ODGCyvMW6GxgQMoYc1b0GBT
ngmVWmtcodixnctC5p9ZHhj2IQATus0gVBP4Ni43V1czu+6DUkK8HXF3b9cDmSMs09Kev/Bh7H3I
rprtV2q2TQjvIuEkXlZXu5YXxyGrn4qWW2y3eDOs6I6l0Y7/zkvEmWiR01l4/0dVq7lV8d63qwAW
pZtT+dkt4m1aDkTq8zH1e9XTKMP9hpk5lGyJ0CSAnZggffcs98zfiBrEyo5J3h4iJtZWWZaruzdo
caTqIA5yZlNG+Osj1Ci/Oi7ZaPGIoDIyD83b6njNWCM0SQ2tkjmcW7QBO51Boqgs/AOhJMJZV29s
lyAz2cX72e2s1D6botMAB/E3PMIHAgPBH0zjPqdjXzc9Ja3rC+kHQstEZodcTbh+5qEpCmOxb2lO
tPeqi47G7K8pB3gX2jI9+X0feJbXyuKseh3iaA6d8AmKGz6hyslX64a9/rxYYEx7A48OQDD45RiR
y1AHiqAm+Od7mFIYX8p/iQ0pwLtyWfpT22zlm3HgIBuybOW11x84iE2ZQ6U7i28oFX5ZqZ+RNMB1
OqBadHyw4+aKpyaGR3QcWhp8I6OToH3bfUtJRqA5U+h9I8v4B94BM+dZBlZ+pnmVQPMTDPQ0Rgvd
tT134LWlLbgk8R4hvU+DjTACx1hRPGuY2vJ/wiSTxkFg2vk95Cc0HuZQHgey8Jvan0u6snlBEVVt
AdEu58C7OQFcD+AUG67zaIV+ZDOCcsTaU9DeSu/2/tk2O8q3L59k0s302vYvHnbSebhwAf+hA87D
n4sf5K+TlSdrE08QhEd91xnqu2/2qncLQrB9ZuszWO3I2oAkzPSxQzTgVZLqFeKsiCOEy1HdjqKk
6/6TYhP7MZC1fixhHcMmFyP7e0WX8KYfHVaiYJDeWmpbgoVLuC3WMCGlX9CtuyQceTA+OzpFAw+h
LXmwFO39LhZxPXu99n5OzSFVFC6MsMnsQ2ycX8avozB6aW4KNJZRSuFVq+vSxdoaFuO9znvUeJ1e
K4m314oq0+dsLe7xv1l7d3O8PQTZ7m93AhS1kQiSYwqmMZaG0GjfTzhxgfWzqzMUvPH7isLnfjcp
VyIquzcKmXBof2GxFNQlGtAvu8mjyXXeS3naBDIRtH+ICTxFyyAOTouWmbZgmZ1onteUmZvSHlFG
dZUML3r0aAphV7UKLa0ZIRVI9CEO/CCldp3iH3H4ezU/BrwISxaWlmSLRpZCW4VnLRkarbKsjAJg
VHQWSJmQPgD9jrJdPzyocmDAeueuHXrhGzhOPRr57plO1fIbWdiQ61HoiKoWdaxHqUHyXV0QdZt8
lc2zmXe6ARBE1tyQ5TjFP5ixOQmu2TgfpHVKnM93K8w987oQONNRK3BS5wIj+JKGQEYbHyQjRict
lszXuqznY0pp7NmtoAsUqOA7D5eThFiYyCtK2ZvaBq7J406/g1OSwu+Xe2G9yzvWX92TwKH/cia1
QEzrckpzwcmjeCpkoBnFlp4zC25qgNU8vKUPCVxz/UPizemExnC97Z5Z/lkXTQwodTPyA5mS+acJ
eUO8KSEeLnfHtHWG2kTecwf2Aju+xVi55aJVIYZJVTNAD0Ek82Mo3hXeSy0llLYpodjY7/ZHXiUw
yrQqxn9l07koMXWN5An07qfwKo3HGLoDYCI4XxMLWEgvncz83kDFTJpDwOfAAEYjehx2axX7FwLl
AECbE9j7zXYj8U5KSd4lWsm6u/ZbSisJI0veob2HJi2DoIwEc6+Rn2an/BY0zoCuZ0+dxwOad1oT
xPtGqp1ZaGv0AA3MuDudtT6Aw10bGUwZa1y0cZqyFaTPVmywtEY7VhXuuZBwa5pqvuFxROAVuun3
Mt2mKL5AXzcDQdjtwPGm75fyE9IGOYUg5e/KfzF7jaTJGDBDBFQ/pvuM3gZRr7yjZfLVAw9O2f6H
j8e7/OdrNO8ZaWrP6JfMtkZDUtDcSD+19BJuVP4KRK+inG2N8qykpw/eHd+UVvONP0NCEFFz6r5a
iZ3Ag4hNnPBrKlwWUbHqKLRBzjaljeAOaSLlrCSwn+2iT/IppJYxlpxTGpaKSmVag8QPfmzHgClw
nJ6ZgL2Ve6vFei4+py1rZrUy68hbm9Z6853eqj3hYD9qF0y/u4THGNaEAxeKQtxOl9zvKFkiTyKK
p099bjLnE/SDJYi1WeZIQJc6HgqfoxULuD2QBQy0OXJL3HLJ7Xrr8P6jEfaCvpsz9Vtr+xQ9Ip8v
s3rHKAZZ/1EhbAvhL6cBLTU+/U+NTAyN4takYMiuuZhOkDCvpcZdQjD2G7ni/FY2HvTS7mPQAgiU
sgw1Mh7BGYPIiK1oHwmgx3B8I2sf0tShtva9Zc7l6PkoWJb599zGF4BExzgz00ZLT3yVeJIqRblE
ALHfAR0yDCm3VOVlztkB4VBGFtpiVl2ybgcB9nXyGrMSrmqkXmjKhG30r+TOlf1d2W4buNjIECzT
FTzLevyoHlZXsi+yOoZmMoMtb+7oN4bjvFdyS2TfKhsUw3NqjOgNC6l0M47b/StqtWVRKeDWxxuj
F2q8YuS45XX+2+tGXf+lpdx2AVXMJgVPd4R0J9qouHR088yProa5T8iRTn24qbTTwXE/5w/N98GK
51p7szTwECsrDYRFkjEHYJo/37kXmjHwdNyoZzZMzm0mzDVQyIl6GkYBiM4qGPcO73aVi523ggpN
JAosrjyx5je842ThU78rRlIx53lJGXQiXvQ7Qiw7Ft4CdPsOneyRRJdER6zjPejoxtLcNnBTPVJp
pEQ2ZO/wwLT9LH6RhHUSHI8dApeQfU1iOSeNDJWASYlCKRSlVla/Q2Sxk/i/bylzHEaRvyG6y+nM
kFAHMP7AYBC5MfGxgN3L7sLc6GRzm4DzXghIGZpxSY8S54XnUEBth1g0n1KpAUxGDN0TUOt/MOsB
TmjxGGPeyohYhLUnNgT3oH3o5vGllFgucMZRZQLOqiv3qzpTHEhi0e37L/fSxuvE40gbGbtJzIt5
AqfWW6qHZO4+RKY7l4DqavkwDS220VM18/HWfGX167LeW13YRxhQzzXSbG0l1QgAigoVj2Dfopzg
m42v/8ayauus6aAWT+oCRxu8Ji9tUcPUd+UXdr+5NY4VlW1H265qsCTHbaleHoSHhu6kft/odfc4
QDHm2Ler04u506x0+tvLdY31re8He49IPyJSerSaGntV2d8Q5ocvWJ+uWRoI0hPNhhX2xGBeambt
RVbr+QRQXhlY888ce/D3UHliRmJKdNEVkw8yfGIb+AjGfVZ1VRy9G2IB5OKBgUDwWmVcWqv2pfQV
0sx36v8740O96KIY/Y9x52nh9ltYIajeHh4DSzlJ4FHAnIUrO7ITigMMZHQgNOD82wHmEU8Gx3cV
11KC5yJauEsXQWPvISvlQdXK0A7Ze0nU+BE3z+TlZrgBTfT80bz1+LT1clZtfsDTYUnCvuxos8xS
jkK4wr2Ro5G1st9ABAulBbGDhvOJSakFsYrMsjyW7W6COWcgOxomc5oJHX6SABCoyOzAUb5JXMPm
SJB93fshsMQqeO7qAnypTFtpyGe18B4z9+7t36hCUdBEstNDhun88LW7fjVAon4b70AHrrcTeH+y
WJvUBreqah2JInkqhrQQxJrL37RD9uGlrvsw1nyMy9go2tdLQWvg403fcj9okyJ6GcPVm4CwPKgD
a5+bc+SLihftIe4IaIoOJ1hGR5BEVOum6nmtBlLmOcx5GbXT1/D+Foz8vmSl94+uM3qhEQ1PXf1n
1RLexO9HLWFfSVCgCnSCrxyxz+BzbH2dlXfy8VdOjruYOs5UXJumEinpFdSarrrK0h9A+AHWhRG5
Eyhcp7x2YfvOezYplJo5muLlCgAcA44ANNc9wKreKgCNSEsgdut9UilImpxw9ajn0x+5wzMjCyeF
ObkgpkRbgEAHUq03EOWFfEvPQo22M7Szi6rNQ4tH2jl9M4smeNRNDKIhGYX4o5PzgqjvhRRyosF6
RyBkMe08StvyZoZ5WfSQYgWp+PPbgH8bAktufnp7fEuT+loBq9sBsu4tOj2IA86ehujYYnXJMOAS
aRKYN5ZRs4fArmAnK8a8p27/2vcUu9zMSig2x7MUbi0ZVWrLqqF2TOPvlbWOJfqJytmnjFytoXQT
CPkyJ4up5sisEeqrAqlf9zl2W03BjFPSl/CDuGjGOI6uys3CDiLi0IbbY+8dgVGhXU2jOFMd08Th
DnsFvLuNuWjpdY9DOzDNypiQ8NjUchiHxRnF8o68jpCPXMnD73PD99kit9TuT0QijWcsPySVesP5
JF9f9tGZBefjOTbdEC3W2JHqhX4h3V2fzfPxH6E0tti0lOo4M5ADuVYIW665/RCq7UXQF0EDYGda
0MocZeZNbAlkLQ5ShozvFRVLu4Wr6b0p7IumCp56l40MxW5MdyOI1GZjxSjOjuJWHel5FpL1jDm0
R4+xYPMExMoi7L1Ki89tUTmMulrYgaiKOazC45uaqEpGRaiESSwrdR/oPtvxsmCt+gnug//52tZq
EEY8hZWAvJ52URAQSv7Y3EtZSXj1Tq3rhWLe/bVhDa5X1srw48g6pOMWbwIvYOS3eyQxs2adjztR
rTCeheWO7wbhTd5pEJ3WOdWLOIWjn7QeyWgOld0O9oKVboXqVrD0ADtL4IGAnYMX1XOU9p6lJNRH
UGKCl3URRR6WRtVe6sNOaNgXUmb8hnnqK8ppQa61oJNNQNKw0WvdslnrC5ZEZlUH/yxuh3cQ6XfP
W0r7X3PvYJ3k64XT0Ajo3maYAlQ2LO11hjidnd17bAchCFn+Oew6um0oaAS88pYTLcTxJ+xP7kEj
oai4ZXgp0TOOiKAi9MExsOwuwz2T+IBHCTm3z47HWeNZ/u4xgebWZkSaJiqSDy3gI9xWSKWBANuU
rEGHVkPCumZlRTU7D7+ef29Z7WqSt3qR8mk1asxlhIrM4VpgYK9RrPRYzQk3THgK7/1pCD4BB3TK
l0lvTHAgaN5exbLLucgL1sp45jh/A6TbW6sC2XfnLp1bUefSZu6v8ozReIgrSdXzxEot4E844FCg
ewIr0jQrBOcrh42ad+heBNvmlTBGo+X9xBIlGzgCZ4IB6GRowOMnD+yNd1WPRzukj/YwMei8yPHu
hVJQ//NuiX6bpm97ak/VT85MAcA1jO418y2tyykMq9OhkiOxU/27/y9gf+lQIAcf6Tb0Y9x1QxPv
16I0Ik6pm3ujESJ8Pzut2PiaANW+UTyR3mleidOA+p9PN4k6vbVv9y5m4yYtWGkyt4RTie8jM3l9
w0vl/E/TQRay91ijbKClcbn1/7e0m0zQYduAC5YpRgTIMbv3XdPWOuJeeBzms8N0SK5ZJwhUJy9t
5LUzCb5WDfdiLt171UwP5qYmenx+IeyfnszHzOEKJtfig1IUM56bRrdj5r7H0sFBT1SnK8hYkREw
wjh6DkFHgmp0vwxjYeZDxoUAvJckUdefsiAOdjcfYrQrgNjn2NCc+t0/7L158jdzNA356GszLVyX
qH/facJO9QTmWQDJAZgLsLD/rV4ToJyW8G/xThTR31bvZOPUcKC27VIyuZ/qYltQHE1mwzHdkYdr
/hI6s76MjORWDsKpKr7YEvKe2CJJSbGTWdwt9JYZayyF6iTMh41n7z8SIfkHzlSyr7HE1ALh2hky
Xdfi9HC38qzmK4+kkkNPIPJlK5R4HpLopWkLuZsru9gksU/6/s7alERQFxiapwA33AMHJEY4wCYn
doCt0dku5MJCZWbfsqIvtLDyFgZqPkOAZArr8qvq0NFDPC/D15nPb2DhsyHPzROLt0P2lm06KUml
CuSmpR1+QEXcAs2eHx4r4nytPu4iyVDVOVxWlYjbgiidqi/yR3hah+fqKikjS7Na85Rx5aECsdFA
iV15H9tN5bET/2DZuhGVClwQiDzbNMmB/an0G4L1C81FbmCJ9Y2eSKbp7n+m8eAPtvVSN7dS0sgG
c5ahVRYi3FnlGl8Sda3Nb/lWaFpdyzm6ZjigjllyvMZuD28byR5b7FD9mBA1AyLr5x43fQ1fLdkI
t6pEPkBgK35uM08qUqyW0RoCV5ik7wEC8dhc+pvoUyFC1zSpRqIcYTHjPGp/eydVFqwTnh6J3R5m
wVA9kiHgvXbWAA0T/kKm1UX49PIOLMz6wWP2GwzWYwNdvxWS0lvye4L4uYDDdlzKiEWVa2HBZe0u
xG0Ks+3HRV8w2wPlYZXrsPaOvqMcr6BfBJKN6RggH3FjHtFvhNh5OVAgFZi5Iju0ZtnYxBvCtA27
qnhSfGal5ObzCYASAVtsPwhUtuGzruaKGysqG5a5pL44sYyXXpk0UuOMp6nF5k+C0qyAh8T7UsU2
/U3e1+IbDHda5EKALAdJiXo3kqzeNQs9HUiqyD39ulbWR3gNxBsZt/kN4XH7PMiO+NL9/wmcTgyQ
kpkbJWIR/YM7OXgd+BajWDqRumfzKoXbU01D5aKC4T1/oN+fnI3BwrnMNawH0E1q4p9oUPXgbE5U
bhnY1Lpx2sj9SujDeRCOqxAdXpEwKj+C7XWqgjUsi/+cjhg5VwBwVIhRGBeZfFO+XXfPTJgNkk/h
S0y+fpL6tWsqLaxEpywTbTiulTnQppGJ0+g14MM6ctAxS8AKVxw2JbLeCVgtz259BOsamm5KJC5m
11HO1HEuO8WcEbg8Eb81IEb1XlUdgFOJ7Sv9EtjZczT0r29iAmVnKesgUGnh6uiSPyUJBrczJ0Mm
mQK/p5WiQ4VGEw/n16BDfful9i5TyAarXCV9Bfj5vP9nuvf5tCm25+lhgRNltsQ02yiQohxv/B66
Rd+1anPElQkJ0NhxGYvxeYLnEuTbdJ/p7YQ2hINWxk32mIGJFjzJ2EfFsIDIw/Wtj7Jsf/OxIvFG
8luWqysGutVN4LpdZohZ4HjYON+tj2dQDPbESgZAUko9vD6xMPVN4iCMe+AnfWgzzMUN+xTASVLN
v1Tk93FroI2p8ZT4fMReeKWAaGmHYhozUCFR7fz6jCxJlHDA+4WnxEuPH+Qdo43Iiu49Y+K9wAGa
gHLauBqxa4HrQZgVUxvQR4ivsQSV2XsSzto6S63+fFFGtA7Zj4JfLEaGSCq3GQvyepqmW90En0n6
q+Aa1KDITgzCEZeSoCl+M00ywRrUFxAUsS7Iv8ztrsHHgTIPwqMA1/9Xpexn/VJlGyTKBBLp76Zt
w3/eb8HvFf6hEQ6YA68V9pcbqh10xYpbHuctYRMppl6gwxOJqceiQtqFQqh/PBItwG799cXz0z06
sIySgc9OSUaprNT0f8qXlEJ3dvQaQ+jMPJBOwQaqPU99t8nA2ILFDf9GpliUbXlpGN1KCGC0kzZK
ni6sfVpwJ7stU7GG9fOeAFmBmkaiXLS6SQdS7S5oK1jN9HvIYFPzMZfXP5nIakl8Zug0y6tc2+fK
/wkzXqXUU429kkBU0eDUqkDYaVFRKVldjqty51UrpgK0xXMI/bnsJ1/IbBNfTnxQPfg19I+l6aq/
C9+cBfYuiAipcTJMatwN+q9IHdsYT6QayLucg0cn4uTJ+fhB/B3KSsJDkrfSBjl7zqjiFPdijrFl
mIHNCLRy0H2PgKAaHa01Z6yGoi7cO7irQVcgMI/SDySs5NvMzqSxUnYEa8zV8a5LdZ6jdXR7VpqH
8VSk0aqSJC7YFdf1G3LowbRSTD1V+57eGpYmYPZgYCRf4/9mCSBjBLMvA48fhcm9L8fALly3PNYQ
uWWpF2AlTuaSN6EJiiLIOLkMHs/f3Xr7J0rHdbFjBdFADN5WmpaGwMW1SHp6c/ZFjwvYgXFsSVfC
8s7Lf1uZalIyI92gC8VmixTOn8exqQfaBEJM0U4mmSAOzYNmhREt1DE33X2ATAMSEHGl1sMD9SvT
nTwG7w4XivvNnyYcvGrWFSZ19CB+fWpzX6hlOh/TtYKd7I5sp+pEW8mN26JNjof0Sah5XiDlYJS8
NmSXzIrUpaCk5LPjZooem7i7I0Ks5elIDqB3J54MD106vJiV+Zysh4T6HD9SE2R4SOTjU4yW85U2
IxMFGnEjKyV2zNchT5XYaGHN/3O1w1jgr1VwJblZ7CMset8sO/N0FOjhXkfQaI4j6cdJxKYPltrp
JiDzlnmZggYemsFCjKnCrNjI+WXddG1zvLzLtH2HtqAnqaWdCD4ee3zt/VMRat19QfFD6kXZOfRn
SQNaAnyKHSaqv3MqSaZ882vkDIeUXGK9vrRrwOYAWtoDHK4b5oWt/oirWVr6A9RmDNsLeS8Yl/q6
RGU/88wlMyHio9JNtLrr/j0PmC2W7SmqFoQqo6laN7E0ctkt25ijEzTpvYwFZPixEjY+tyQFZwUg
Y26wF+n4yFSBaWgazWR/H+5R9Wk+lz/p5Ul+s+ylLr4XeNf1GuAYsXrJeZ2uc27W+skHaZT40Yth
XNijQw8Jxz7/4jBjfT5cvMQEtu3fVkSGihQkPD3gxVUkDBQTnweAyZLQF8ea9hcMBcsdIj/Q1xgS
JfHRiXBc/pKY/gGjTRdmMaExSReG0e70i8++k3VuLcobvj53HmbIgadzm9HfDg1aF8o6jrUX7jJ2
hT8pH981tu4/MmwygoBbgIbcTtwYqawjBZalGmNsmFnhMk78wNHhX8x5RkYUnclhSv5tLpKTaisE
lnMxkRjHX/rKJ1TB4alU/Z9hJapEhwKuQpmHlgfnQKgt92OY2v7o2th8WvmNmfzhIknFyWfg39QI
O+vCPD7MVgwQptZi39ynnpdqK5nt4GtIGoJP+LJTv4xBlSw2EThD0ewjWXHcnQ172q6biH9amHu+
g90PSGPTxxKA3cj1wQCv1JsTGkNSe2bARy3hPxH4G5wNn091B6Aa+nPL457p1xv4ncW0RbgMM0+f
xaRhuXpkoIqMvhHwrgYOrDMLm6Pl45Ei4wLcBy58h2NUoch7L+JJVdEmAf4lDT2TKphwHQfQu04D
HkBZF6m/i6bwVunaLD/q+o0j/EITxNiRFJXFNt/x2b3+kNz0wCiZoi9KW1GKm1qigx/cbZHr2/Vi
2FEeALXjp+J9hClNEo4ivDh69p0J8qFQmImVWxZwT0N43CAn7TaX1iXpdntcoXdz06IuO3KOGU/B
ejdKzVxGLRV2VRCjNz1B2RDjVT04YIvrpUUFOcUlBjk3WLvV1xt9sPbRwr7z5Xdn2G+rnhfsCx5n
In9bCFmh4oSC++VPci0NWsNDmZVw7/IazY6b6QIlV2iefa9I47PSELPfypgZA6lZZtLXD2ND1Af9
sfFakqZM+vSr0eukp+hXj4tSi4wXu7+NvPh6rpCf/sQHr7ggRJ37p6Hs79FQg2Fbxclrc7QBUgzE
fE9UC0Ij16tLpJefBrSiAoG7WqkYedYpW1O7pwCH2CRaO5Iu9K8le99a7dldVjF3wwzOuh4AHP18
mO9Aha9arB3sa2yc1ZeE3zVrBojAZa455vgy3uq8KhgVvaTiPj56cMm6xZWElO487lDquswth6dz
Bf8oBtdgNpgCQz0ae8nf+UQ4EnPAHOpEIoKHZxCz9bN1Td/vd1gUt6usue0PigEsEtqHfGvyVhyc
ZOXir6erbwCjjZAIzyIfDh9lqKTG1S9MqrDLBi1AOAIaGVUnHbYcWNqSsyRrAZGjOX6ENJN3vtWu
P5KnmDogkvmB3+XgeSZuqPka70d0igK8uNiQjatbBDLoIyHaPWAu1euWzuR6yf6gAIhNNrgC/1am
7D/CA1S1wikaElNDZPa8Bq9GDNrD1DJ0dk7zUPzL6A7Cw65qRBATyZtQQ0MCudTi8heAn3GIyuqU
VyXfShsCLEhjWxois56DZTFvx+c1Hx09Tc7dObpN6uba1KKhWr3VI30PyRuWhAAe2G+CMZ3wYDiK
SwY7YTcIN/bFM2VB5qalPetA9gfAw7lPXWkaMuNN9vUimsJrzqgsJJ4fx+SSAE6tu/GdNWoEMOzv
0p+wCO732uUruw/wC/PkW9TjwmUcd2YDqnIZhGycFV+0WpwVMPvitcCQlrevNHWssD4fvCwJsb/Q
PnfzJI3AkBGOHfIet41QRjZl2qq2jqb/PP49Kh6Lo2iwuK1K+swTRV9mlVU5UOzVwcyAWEHWVnqj
HlwWdsD6PH4lJpM+NGYxgQ4fWv7Qe2YxdPi/6IZH9ijobXgUmWTtYTaDbUf5Jv8xr+/OHY2tY05+
/UQTUPrKYSzXDTk4WHZLJvnvVftBLiCBAV99JunOfznWZHA19RFPIcoGDOJkPqWE/xNcZ/pZ7ZMw
S9+FMsa01dcv3t1XB5oiD3nP5k1qjRo+NlMXmkIFPrlSWTY5jd66Amqsj6CKFmLIt5Ntx1Ut3fPc
OYXOirJ7ELhOiTIU65FeFV1euoJo9EVmlbbLcclzEOpkMbLG+BLAsWQ7i3RNPL7n4bQsxLSnWK6q
CdeabTGUtiDi6iq5Clbj3OwbmltBKgP5vsp1E3BqReOlj8ehLECz/JCIqYhncYahhzKFJpEj5ojF
kvdu6BtQ0bUlQiVOaqC2plXqfPtrsUSQyT3ViMEnPoE+m9T9brHyVUA/0ufvPNBXBvHAIoNbpgRf
pkFqB57vJcLVd4bGOu9/CxNdTGTG1D+oeU/cQHmK+W0q21WYAAojilYW3sU+n3agBQA5nMst6y7k
Su3DAYS7xa7YHxRNaGmS01R4z04xgXGEzKli5qGsEhoO+qxWLfL0jKPtR4rfxsqIdWW/VfwlXgbw
wfJaG0X61n9L47CohMWbDf/4IM/k7l7tYmzpEjlRf3f1mH39qu6Wmdw4q2Eq7bXxTbJ8e7Oxutg1
9WE26VZbAG+UMqpHbN5yn88xxWD6UdPaphJDbKisd00a2WNFVLlEBuJMB9hHbL+h5EIs8owaOPbS
NEDYNmAHKZW+PPIM1da3L3tUlIcGRT80ngv/m1Tz1vbLw8fTliZQIAhnAxkl3T4W9sBRni7dgMMU
dD/bvciAG5J3/vk4N8EgGFla7EIvXOuEkDU+xOxDaPTZyJzwp3Ry6JqfThsRPtgeVMu8zyWWPTmq
V4VYFVBEZUeVsI9GZlAw2sjqwfeE08WBaWw9p0bsE0ceJ9/BSQIH9U+OpVpN07YD8hMXcJu7oMto
aTIAmnCNl4XnxIpTDVyNSw7Tqhvcnds3o8Ches6oXWk8mPdrchxgNEwcih9uh2glKiHWTiwZulTq
S2W2irKxCmqAM2xJ/GTCyTnpNe4Ztg2IUxiEHHWdsxofYnsbitqdmaZTeyFzMzJUEMY2OQ+6nUAL
H5fLGAUKfe6wPxfOuTmplR871qgk3clWZq6QM4mBgFCid0dNAEa+dWDNsDH//z4hywN5PFCeOjmL
i4Z4VJvFx47yVhbURM4h1Q9K9m256Px5cBVkl+9adj9z4/BGWIKhNQqHIDZeyJ2C3sWG6lvBqIuC
nnvA7CfhwaKZDiQBEVDHSGeSq7ihhBuiR0natpelfL2QdH3QXykxJnPekEfoPTNWbIN2TdXmWfuJ
z7X4iJE9Rjlcyjm2nbNhO8zpHKvOgtoIgj/qg2f6g/539ZMH/nNrUiP2HEl+/0Ue5sahujFgfTps
hzWHFmfhMlWTgrzpsSJd3eebjM8ZlVH1ts+MV4ifCNrsj7/nbrOypX4UQhXkfkZAejExn9+BeQM7
jRhPbydm81WdVUM4DjKIWH339IrHs7oLairWpJ1UuA7JTgycd4CBzb2C4OwOBdi3zaHoZiqfAF5t
glu0Ara89ecqoMArlgBS9UWNFPwvi2DOppu4p38TUK89qqCbbFQPCY062OJ2lvh0PcqZedmlK8FC
YTo2Ubwg28gAAWvopGFjKLpniCnfRg/94ik9B5L6F18/yMQdjnB7Xl9xJPGSFX271HI6zjNrKKFS
1HU0WgMnj5cmv0W1R2D5Ike+2KHE8AQQdiOpmeDgHTxP6e0x0w6FrzJIRo/R7wdwcmKDGLMOIwfU
hJLunGIfMlVD9m61cvjs5WNz+FIsaNduXXVbnu467gKF++yiaTpap++jaR5t1Jx3QmGC3ipSQmKT
m/fV/oRYHR/2O2zN/IGeFL1HhRRLUgf7lmTZpGx2vst86HJY8L+z6891ykLDd5EH1qLHfxEAEOa0
+oETuQPGDQXszmg6BnLl86z5ySoKvMuVeXN2dtlv79nUack6KdcDBhx8Gnce+bxqWenoNcshxdkx
fVdEBTAwWuzFxCQtFVFnK+/aQvTAZYYACzbvgva1nQUjl1GaJEqMb/dAyD2yrXHH/nPPwDGByc+q
mnaNAdKMeNt4dnslNb0DmwhppYe84kIvTOJ3p7ZKnQg07ReSpLUeb64+i3//6v/nm3FtVAWDCsG8
dMXj/cXHKpaxMhTWFvhI5xx7HHbdy16w3tWHUu8W7Koa+aci9Uu+WXpBJm9/nMhquMz7/q26dqRb
IRcw/NdLILErrhhAZEd9DgHAXOnSK3Hkp1PPypIBeJSfj55wKlOA0/mB2UP75k8pqKaioqy3m5vE
MztLY4isMvoluhJjhAyrGg2hGLN9DFvTOK3eCEnf1NvNh/CPgRJYUzT44AfNxSWeXIMjv9MlLD/1
+wZ4LknsLtT6FC9l1mz5cfWcJvqQSdn7XomIteJUPAwg21r8IU4k1eR/kAft5HF6DWYHygeER2OG
56APeJ5CxtGPojBkM2k5AuuCMlESxP7TwHiqummnIUsET2tB7Tyd62Lu/ht9kzO6rcFnRY/sp68q
ReRqsK5zoqyOyIW1MSfaA9fmDRVJip9/IYGzvonXvOLUqpvLmAvHdGXgi7ySfx0tB7fxKpyheOlr
JgzOlwb9ClyXjCrJJuCAAm+M5HjAbKZFjz7tM4nu4bL48dr1svh3CE3x6E/vzc9YSoOauuQf6rgU
RP4qeBHs3y8VkAXLdTb/coEjpWLyyVcy8D4c8TeRZjcotI7fqZTPQlq5ETMzhyc8TR6LdXrMSZAe
5GmLUh/Td8jZoZjoqN6wQRUymVvM8VgQ5MUfvpC9rKPT3qKODzMlDT62aoIOvAnj9ghhcN74yhsR
FxdIhFi1jKnkBDa+rw3qP7eyAWKTChKFQxdW6GP11eT6GRZaqwmpSZ6iHz6rZ6krr2ydgnh5zCMU
on9+fHAyDZJTcS2c1Obv3KYjL3Q5sziMDtnJQnmJsbc+T3+yB/HqA6J5b0OS6LziL8MK0f2LwuBl
FrBAUVaB4rXEmCMgkfSv+x2gc8q47/w9nTGZk9IOA9Mob1G7X4HR2+nSWYbNBV4Xc597G7695Etv
mO061qyGBnnpVULLkIzEMogAj9fIq99b4WqzXbEj68AJP6/JOhpq0CVBmwTpAFIFaiw3VUh8eBnG
xz/5inCAcIKQvl7lnKiR2jvoMuQ0JSA5CEy4q87t+l4PAjFjwGjTHJQ70mHclcTvT8G+BIDq4QzQ
48aZVSiko3DWoWFKxEKQ0pBd00MclyCmS8UyBr9xUBNQDKtYXhn0+m5my9a6LtVNEfFMUdLg4oRw
Eeyf67+fdV1i9qUSMXuyUuo2Df2yrxLa1PfvMbKcy4GEaVfq0KQITpNxCC/wmRsKHorFoEkIIyye
hrJ+DOXQ8bxfGCcPDaR4OdDv4WS+m+GfuGHm0xnICLLPG8XVOguMCa0AK/2ErEPcZrJxmg9R8q10
2LVVNJUCV9An7DakrQAH1O1gEhT8szgI0eFK+2Z6Ilk2fPKmMN9x/D4YuBFhUyHS38EGZD/yufjp
uxRQt/vmhKhRGqgBxphdCU+gsIWFP/RqfpA8vUNAaIk2F3fEjOoaYoB6w8OKK3eN9C55KeSDHiAA
WXqNac2nXzoDJONGV2UI1yMk4ufj6LVgCqKCM++BSKkhYoRopv5jGDfxHwKF53Mwv93+0j/arGcE
2/ix75guul7bN3R10j3wQb4F2jHjLBX8wR1nNVJ/vUb+sGXeZDwvOhlgKWVm1FA3oqE8k31GrAgj
xedN/I4+4gZAEUHt+8qtKTI7lNqwxYy6fdBw+i+U8aXKIHdEZpvMM8z46OPOrGwHuCkx4FSL/we5
pBk+VSfBB+Cj2QtVUx1EkgsHvuErd2cqTlK5WUHfWMpLyeRVBp5hZqr1OxfSi08kZkFe1aV/RA+g
y5VBVyeF2WHAGlJU4dQlUH4mVlijLjNB+GtXUnk24K1A+yChIrLkWvsGtSFe7zTe2dh5gvRtrlAa
gH8y6T61hJW2pv6irCzyuezcekyDYTHCdmUqEgt44b/ueENb4jwASoJvsvV2B4XuYZbh+Lopnuip
nu4BvcQYMr3b+uCygVNnw4UHQorX+jmdJlkX35RgY3pYe5yrLbOE/iVx37ynxHEkp6S7sMqn0lUC
r6iPGPOso+MAH7e+Al/Fgg7YsSI7onoHguTXglg97bc3TP5ZOz5GRZFKKA67xkr278CX5vxTo4Hd
vCBhVkqliA9F2eRDjdZhccxuN9ZARSNMSrlykPcr0v1J4AeogefAUxLHDbVU+Pc368KKhJMdOEs4
76QvVVKWZ5U1JGsKPQOB1p8Gkb/m+1ZL/50ZDBHhBRg21+TBLvgwn5X+pFERsg0zzmfcKe+QfV19
VlznXCA3fsPY5CThdjkWCvuSQFKLLky/EYmh3CppmPMqYK6kWFHgGd5ck93XAHCKAkZHzQiEYRgW
PDkiTPPiLh0IFScf20tu4PFOxr5n4H6pCRyYFBaaDxU6Zz+Fq7FfgWGkN/UW9FKKJJhOKpYq4vbr
K8cCZAVA9bTSLLP6HWOKAwHwhV4dx8J9bQiPSBJsXh2QKoNCm501XFNiXBC1ThI/LoPElFItey7r
2bMnFNKrvKsltmLyq7UeAE8WkPsRy0b3M/UHVUQ+obxwu/enRHm5y3beDOTd2bWtqqcxXsMIgcl1
ZFMWGW5/rzceTkGSJpdClhbk6TmtxudKj/c/77HJnNqqNyl70NfTSoCP0yejfo3k1cxhNzmrsWkN
IoQEp6hyruVkuguIfyYkgUpYuplxDtJsqU5tmN9YURkiRLJFDOduvkM2UgexF1n6XSj7PLGWvIIx
KTeR4/fQjeSaqomAIaT0DqcTT9drEEoZRRZZq9TW3ukrzriEbzfhtT4/pJBVUwUjmaddoaq1a6Gm
qZBTvAZZF9GNt93jTezUI9PxzTcFAZqeGiM/tx3e8tsYu113i2Y89gilJI90HnxS/q6M26HCYHkc
343yXxV+8Gvvb4w4+hg0Ig/1xDoVhHE1nteYejAiH5/nNKLrqCNdfi1T3gnEEGvBy3rY7yEUvUCG
ZRWbHODWn+S9v53RbSNGrBIx4k5JFXHvGUXvzKTg0bDMBkBeAK5oIuOfZ0HwNC8k/lORs9jStrod
mupOJoU9DwPKe3OJzx1eES4grcUKvv8eAZwSUQkmO4lB0eUJ9jTEj+C4O2y77wpyo1+TiyclqdjF
yehUb/3K5fBmRyTMbtg9QXGV7m/i6TfCWzraYHzqvjnpqV6Tp1gVvxxuMXVYnCyIiSM9iieMLRI4
yrngg8/Wq3S/mtuICjo8gLAjdFUOf8ps4kghNcdPUn+9RVrLOndCzYarJ/Stm1v9r/r9WX1wI7kU
Qwsm7BtTP0yHC8lWKzf57vZGerJXbD3ujJfIOvFhMX5M73kl908An6vEeXq/UnDqlhAvBb1e065Z
70CIw07iY0tzOyyGFbxtbm172ADvJPaQPpaLZ7f1GRYV9Lsur8CqIjXkPoRGW1cFO+MA0QgA2Ymd
Y0U1xYAklG4teiPFDpR28vi0m/IS3bFX7Gg3j+FC0JeFuIp8WygEbdfNBrUkmNxKAQAlNX1wRppB
PjgJ0uUcZkn9NCK9XYKQc6+GgQ4jW2b9agrhME0B1+//3Fs8WKyhBgJHyFjshXm1XEF080UgKzwf
FBVDIUO0M5SdtoZWXSHArzsZCXPB0scp0PS9phYlnv8DrBTahs185h7jO+kjXh7ogYBXOIafPpgp
QOK95dDhNb5fxxNTOCj9PPK9vO5tmYDEG5Q7tWZMhoFGU9WHGXx8IFgt34MZtJ6XPQ/40s+Cbg5B
3PzUZUqLsT9pM3e7kWna4jz74MYnCYPtAyDKStInGSzaePy2eFyOg8CU56k1u/YRD8TE4JTIxYzo
IhG0EQPD4TglTAfEcYYrU9Iub17kIY8VwpvsHj3aEf8ybK3nZZD4FzqqSSuV0WyNDZs3P6zrL+IY
uAoId8kbEGx468zWaBh6SvTcSVlINCreb//MMPRrRgFzrNzi9bSkVjSYXxWO+e1/6S7Kb9E7YVQ1
T32c0CMeVFgx9NqnzDk+SzFK4eQs7z2rWgHYu/XTB57zTO5qw2sNEqTbajsvH7al7ukjX3l/7VW0
Dpt6Yh5gw9Rgo8UPpLOQateNVmBGNgfk5xNKC4xO49ra3ILB3brlK5jAVpqZ/XL4ddqrsSIpjKD9
YjQ1BY38OvCoSvk32NC/6qiEDW0B/pWX1vcPsUu14Nwm+PBQemHvzOmnKetmiFfmR8It9TboA7CA
mDvPhjRfethuL2mUHxu3b3H/6ZTJeScTC8/WZN8enYM/nm1lQ3SHyU3zS9z2eagQ9O+8I/vR89bN
XyMocnVcGsGh/UzKLUATzG6TqyT0H9719ym3khcA2B2Q6gLuiVHaG+zyqe/kQr6Y8EnicKdc4cXo
QFkHnnuoA/ZtY1RTc5Ldyjz0j5mwq9xL5jluxCXaTQTTztI9teN/EhbtmLiXRhpbiCN6s5Rbm/uh
58+9Qx+6IB8/G4W2dLp89J/q6YmUfL9Pd5SsAfawnHUrn72iq4Az18LZyQ3sG7k544RUrn0CtNdr
hJ5YFM+q9+s66hz0DcrEhLHmz6B7njeY7BIMxWNc+9ZiRjqi2f89ysLjqo8P6qkZyP2JqCQ3NkJ6
p05AvSAdiyyfI10IzfuChycy6qgKLsM0Y515vm/hOj7DqMCw1BiixlJZVLmYhA5w/qtUOal8uwcA
rhKoLHtXl08JCuNxzeHeQntUUvZPJoSgK23gYCFNZySBr/kLwO3+yRu1g9F89hj7qC/r12Dgb7Mb
zpnJ9GNrm7SzzsGe3S0+MOMPIjT3nCh0hqabPHFv5Nn+kIikF8MQI4QHgYST3OB/QmW9A5C1CtWu
TLtd7QM2TPeXlIPzR01GTcqT7yE9pCKn1ENig+S7yDM12iXAk/fj1NWr+1ZEJ+nrLCYNz/tGAN3y
mROvj/WD8JZjDMsKaOWgg+USFPbJzlF6dFRozMAy407MfnzqiOjQGNnYGXM581yEj7wpMERaWD6X
YYqaIGE2hb34fgeXKkYJfF3sX44XtolwDVXo/vXbdgZF1HM3+fSPGm2LXIU1JumPGgW78aLvLC98
BHl1VytjLQb961jet43BNtljLbnKM40zpVWPHdG/c8CcAys/Ve7/DDOM6eH74ja7HddiNA0MQYXS
uST8dns5tYWNs2F7T9f4At0BsRhTrhf0yfbZLEMB+T/ejILvcAVxyhmHBHyLaYPN/HmfA6QQiHGM
sn2KO+fCORfRLvD3EPk6qI9i0uv59awPObPveqyOgui66TW3uxr6ukGgi6/LpyHcZLsWQzcWug4k
C86DgTgoyMtFun0WzWGUXlM7PHZqNgOmgkdnttqM3gGQt27nqi1nZnp4fmNPbm3AP+hhoofFkuVp
/RnDWqnZIOae6mJDhIdxMZ15MGSPvZrIpsrFSrltbXcKioM2Z9CTJFkBDLnpYT5EbXU1YvLW8q/4
ois/UHucIW/CeVuZ428cXs9T00rDePKW0Me/Zo5RxY3Z1w8B6d+48XqKd5Un9v1q9CpytLQE7y84
jq++pgvwVb34yCFdOjf020EsR89Nl5UcFLOVfG7fJde5eretw28SY8oaUsG+zOzTA/BKtlc3h4Cg
/VEgaZbLYOsJKEUPGHIVIkHa5HmxQO4AI2YKDn4EOWv3/Ldoq5R5YmNEv6Z7tzkJMndAISE4AcHb
Hdv2tNQeqP1U7ctKpkaAl6ohVUvEj496tpjHBDeek4m/RTC81f6IXdnCGcGovmob8kbIgoXzHCTs
RGVgJ0M6j0kI8fQm1VoCqGGag08ycdoMc4CkLmwDcedyS34VUATqG/+HsDOPyU9oYkBQETnCIbz4
TGAqZ6/qXP82HchP4LQOxBqpqpdf49/dTeOqaUELCSDJGfCbYev8ppX8kwh55ABDlq0H7Wiaqpyi
c/pnzgEerZE+hKZDPN7OHEvYEHFIQ7Hva9AfIamaZ0td9X8ys8HjPStiuQ8abBtQarm0M8qpwVu4
CMd+1B95DstIhmULPtaHsAGrcIwA2KqOuzu5f9uWVkqha6Pin1y7GWyohmk2yWRYY58eXUIpro/V
Db94jT1eZIkm+z3SettFVSvhU5HXLU7GMvfKzXX45V3mKDb3aFJBvgC1Bn9zrYr7UEYOkTBlhl0w
ECTN2FtCxLLTkSZ9nHyc9RgxP11ZgeQz0GcJYdHNaxfDmu2xuGcf5pcb16Toxxqm+ow4yaq5wi/6
5pIsO3j8VvK0zY+oTKSsLssXIatEFjsd6qNKKGY/T+dfiqOFrgU2pmLKiIA2na8iW6aEM6cKn7pG
Huos/Qsg2QZ2VG6kGZRSKRaYjDq1tqBKoVxZMuY6sZesdvFJDXfd0dLY82BI1BAs7lffHJJAUSAE
GEZB3+Vwi0yk7RNnkx22m4L8Y1INAJq14AdbicQy5B4DpIhpzzmFQSE8g5QcXO00sWhT3P8frEzk
7h3DEtGnwRMMH1XOgdmJ0Rp4TfbYBoSc8pwuotAIdU+/WBBFfBd0KaRBlLn5i7Xi20l8ZyHij0fH
gOi1ckmy3kFEBOeeCQP8ANxuketYZWq8PvufPNUD7xvdDb8x/S1vBSD4S1sjuUNJKJPgOTT+hC7O
uCnEEee8QguHyDs9lmyafpuRj5bDTtXtODHZGQs2QhIouQfBsSWgJKta6mP3gHxKUFcusn8kmwOM
/3ET0YuGY/9EdmrrKX8LE/DkxSp1UI3K3DF5MAe3vqMHgPhQFxmZ+gk6b2aFN6evaFg93xrnjJcx
u0QWR0nFClEH7TDDDMfXJO92lCPAoUHiPWdR/MOUy+5pkZm8hlrzs8KTzl7MFwWp99LIWQwXUKM8
Pa6iwv/FzLWSQe7a6cgQWlv3QlyjpDvU0ghOmrs3txaC8tXOHeFjokUcbd3nsJILhREUOYAx3xCF
RxRS1LaxGJMIw2njpxS7I5VdD+xO2d/S4GcWjyyJRmrNF4TKYcTv6UK/tM0uQClHFQxQ8Lx5j0DK
GbHVEOmp7GlMk778+rgpCLurrZgC594LWEjp+Wo0qnAmQ8YyRyev8eTCJCGFyJ0zUwJ/wHFWxwDp
L5gFWLRedAHnm/xSJIjRgNc3ly5zpIK57oXatW+uuAgCo3XCtOqvQUe7lmSuzpRuJRvIHN6r1JvY
TrhxqX5bTwBOULBBfoju9taBpg2jRwijS+od4m4Qo8Hpnn5xuCH5L3Zu3YYSThti+v25fwlL3+eZ
tbWXDRWzCIEXD+2gT5ozeh7xJvqfmepD6gRiaNendodAlkSzV7W17pABhGfGYKoKO2RKirhF3QHz
Hm2VCYR21+oxg4sJwPjTb1356qIJAkaIQn2yhu+/YiyWa2b8rkhM1YZYQ+7izM8nlOh50UYmUzQE
JbdkT5PBQl/mv4QbAusmMszuhI2cxdyE3IFtyTIeNWJ48faOVOo+nSsUHvDtnSEG/bxvlOmoJspJ
urQo7JUgVGCl9rpNS473p0pX5jl+jnHNxleYTfXtugMWxqi/LQeCDaVZJDvYPKT4QYZyLdHrsdgU
uiP81Dly0otvHMDH2n9LdrZwPIukCx1GqiN8QlYw/JdNaDoMZV356SaKmL42tYCEKUDp9obtfNKV
bELkby5zI8nD3WWsI/Tzr7S8K3czqHLxHWtrJFrMX/9CJg1CY15uzPwLI8TrpgBSRft0Cy4lRDpc
KIPNXA5HoVsE4ymRuW7rnrD+Bac4yKlK/qgvw0NP/sd5DVcpIOKYW+lfl9HdEtWe7468gNbQN4F6
kqulS73JYDPMQcpngY9R72aEN45X+NpvEQiGhzZQoIXcjttoeDYyyWgD5bc9M2glkc7/XdI/6oOT
iJvi3dTT6+u/XKGjXg/XS4sw/N+IWKAaZ5Fx5JDmN09iDv1hiyyWBmBk8+N6v/HBOsBo8ZFF48fn
Cuz/880vx0cHIP1qIPVwVk6FpNCxb2GPH57UTP1YgAWCxfTdgRIFa1XbcOv/Rxq9JiajpUXkuGzs
R7WJK35qlxe2Xh0QIwAxvAU/Dpi91lvBONVt4A8xjFvIQ2u4M4y7WCKiN/SewWYR+AzXwBEU//4D
LsQ8VZHlFSEyqQexQ7O4t3BCoqLPY8n3A1uvPI0nBhhi9AnQT6gF+22TQK1l7qlvd2tXNcBxPQ9i
oX/f6uA+LtclMEARp6wlqFddFtzYu4Z+33zHN4Tkkyo3buUm9Img4pDR2Jbgt0JiA0qab5xEKuiS
OJjILbLbHgUv70BYd35mm19cCwDrj7APupxpNa5roYZEtwGEOv9OduE2ApoJWhMRNhumFrmgoWun
+B8l4J40dQ9a924beBdtcx+uep4PrhGF33GhhcbJOX+OdWq8931D5u4QmoYHfVsR0SgVYJyembQL
4kBW6ZdhadyvDWQJNcW+9sG8vV+8MOwPBc01qud4WWORVwGOwbXoPQapmmG1yPsL83Nx/JKsqZ5V
wMPSzIlMWquUUYX816300cjj6ijv8bxR7xjLSOiLljgBHifhLQJNmwpijGZ87pExUF2wry9+z29e
oNA7TWdl3Np2i7oR4FltQSIhh8Z5SjSfCWRMlK4OVAdBwNO9hnkLHZ6S1mr1x5E5UYeOJsKYgjP/
3a0qIXZHUMXkYgrFNcJGSCex5X7Z9haChSDgpyCGo4gQllwQfoGGidh1dxF3IJuEteSS/nH9CBRX
5ZqEM7AHVm3Fo+9PijsHN1k3dwlfjsYyem9AhR91DZtkQrpZsjR8Bxn2gxfeuWNG+oB4ev+MZVeD
7bemuciAgCiX3a9WLflNou9aNvXJCMiV20tUho6vi1AHon0cSq1/2UieCyRFxzfdeLA1ZGbtBLnI
06MTG4osjv2EbI66J+WuTs0IE3DxdOuJPNGQRqrkAZH6Yc1XeDeBBNUaXyFM7SiR4HcRQsNsh9DT
mQDrh/RlzK/f6Tb6zZkUG3YOsUHIm5F2RcXJl/xOKOl9k4qEXtvi823v7YVEhA8uEZdy33NZ+kTX
7DALU+43sq8w2bvpwS7E0MkM046GYHsEsiUS8lZv+d6WlTgUa0wiW5jzQ/eWJs9N7TyIgjc+IAA3
ac+7m1MZopDvuaHHo3ImDrqw8ZsMvI3V0dwZTXq58tpseN9/necrFg7I3w/IIth3Mj0BWKRT4IBs
gwSgAdNY0KuFchrOGFHn0piaZfzSnHPgiDt4B4FMLFY6YP09L5AeFlz907qsuKYeNg8nj1A+wjoc
dSPm73w4R1sBM8qQYz9I6tONwghsX9aHH++Bz8DE0rC6u8Re/jtlY5YPa3r8+x9On3gWS/OQ1ui7
ZjVb8S+pFyj01YDFrjaMLG3OQWguRARfSRoTto+ummN0dMoswrHyLJr1E7k5E3cc+9rbnGBv4L2J
VsA5EI1LSiKd155orYrBSQLLBxljUXYNuyjTxdlfhn4cz+bHEQ0FLnZJtwWZcXH/r/Qd7sm5s9Qv
P2Mvx/27ysAx17bH0cY8z8xWB+COn1jQPggQHGm1mS/+NibQz+AtN2U+pWU8cSdcFvZD1zHJ95RK
obkC/xvSECNnslvPjasM2Rr9dkxKpsaRwDLHVsxCBR3F0K+iEbmnaX1hDoM7Fx5uM8Ob2MlCQS0R
xuzHSALs5VqHO8GYA5ZNtsbhytUmWsrqljehKcykBrbXpNWwf1Cxne/VLPbdZPf+NylGX17hkMoq
l/yLhDM//oWxplkbQCPhJWxwIvxaDVregOYvWzMEemL1ZS5pQ8vR/f+mNvCaGcuUpaR41CZU8nkx
3WFdup1ZP6Sx5IGtZ8/QfGtfU8xAFm+x0B246lJIhpaf9kBepTSh/rYw4fZbbE3jDZl2vjwcaQ7b
pR8eUQAo9+ouypVZh4nG1vzopiLrjwNJRGXRiBeTU68mSgUQ+NMWROD0D2bCwZGszQpcBDPq7hBM
+nxAjhU/RU3XSWQq3A8gCs/YLfdzJrWKiDPApe5R9bXB+Ajo9SdgYIBKt0hEHiyVn1Y67YZtHQRE
XxTcbdokx+NJImv50Yd7p20ftMhe/LGhdPmhquyCiVveRyWbWn7XW7bUEkhwnBOiAg9FbAqLAJDD
FW6juqmDx4DfnAfB0V0ja6aHAS0EGwLAfcErm7rUjufGxAIWBcLfUjCE/sSF2QmUKzHR5tAO9qbb
TEGXnnsC5APJwpskc8VHaPP4/TPzHcU5lKEVV5Ws/DXGVVkmVrHHvlCXNRMIfhJ0+S5CIUc3GBgq
gNj9Ob7HXZhKj1URRhS+w6nspsQ53588ds1gH09grmSL+mdzMuOabV7R+XDQdcGz6sZSLpIkB9Uh
jtO4XZqoNEvhL/mM4JMsurIzUWCaM9zdHQPOzTwWWjO7jSLAcT19sIE1WiceWmJT7dtytK11at1i
DXuMK8atyGI/IMxlvz3ftFNd7k0SqC3Q0job3jC/OIAqiNsMxyatDxW2U1ltsNYSIUNMXPRhlHpg
nThU2iOoqQxrKUucERjO/DqhyyQFJRSFz06SAKBJEuTVNbJofPRNOGwWBfj+ES0FibxcfyYszr+j
0xpV6jy/1ira3Kr1NS9RxSwEuvm/N8vEFjQ64ZMhrIJY0TsMrC8aDJ/UhsIOKGbdaMVrFqfVk9kT
zeNnBsVqIcSJGhj4jeSij0aQbER05+riOsMJ+xvdjFaZS5ISryYlbXTeeeiht5zqILvGZdPX+4AO
qaH3EjpgxiCcriUUtkgRaZKOKDpU1plrLBAg5ezbYaft4jdjs3TUcrXpr3vnu7dERSaP+nfeQtLw
a8YSbE1Lfy6q/zT6qYMvmqT9l6JmsDWJSbSl2jQNf/BeX5plGuCfAWk+Aep4WZI7tUrYDZ96UxMP
caN8Edo+SgW5BnRC4QetLRQgWgVGT4G5QNKGRuChU9JZ7J2VvXAQ41ym+dYJl8WcWZWorN2Vr+UG
5Zu2+KHmUP3PPJDkeFPN2Zlmia7Ppo2W3Mn3NqOroX4T6TqPHoSaImq+eAlatVBXVmTx7SuYQvwI
x52u5Gf7QPH1FncE7LiJdBznMhCsLj/K1iz+mf/84rBb5CU42IroHn8QVBUQF5h63VzQ3uXi8xLa
0Y1dOhAs5Jpo749U/iyqUyjHz7WnQupRUfyVSdN8jiAaoiwDtgHfawKQbHVnW8wzRO0eaJEPyRD8
w2zD2CEwZx2D35sJZb85Hr/bHxWyvGgdVREHei0oHAKgCavIvmEEvgOJKmJlSILYKufugWLwAiD8
GGV6mvfFk2+lhkPnbEEobmPlvG4xpnaoQrEi6wTUdsHESEGqwn1zNAZtsp3x8YQecIdcARZ/T6NZ
T+RviWSiV8e6j6e97BnfCbPUic3/SeodY1kJCQdTeQHl2uZRIMrdJEhubxLjsUGvaLX7byN1HbhU
ERQ0hNo/qyK4YQiyIdIFTmwhH9vufuiSLgkIqJz9dte6kRxGfBujHerI0oz1CvUcRdOctcdj/Zk/
uVmsDU6YDXh90Ok14oK6YNeE9Y293gIL1qYlARKhExD0fsOGrgF1WGDOfPGvuow7BGPv37hP92np
m9JuXA+TTwEgj2Z3LQ1Zpge7HOJh/g9r31ofP6DaFbQqCVuzqk4cE3rLqBqaGz5SwCfXFq5aGT3i
HQc0/ZNTvUsKLrCR3UhsZTcJvMDQJ7wahgSnikc3D4H9tpAR7iT/s536vbfMiIjtFNIjTXnni44v
xGBcWEDWPvaU5W3s8WZQ0yPzOqRHEay+gxVYV1A2w45uCiLuNX3QbfwcTezQe4Ee+E3DPXnuLoc2
wqFbIYwydA8Zz2dq/T5OsfEWIvqjYatDI+JcnPoWk+24zdxPKfbMsxv38d0U/C1T8BH4AzZvm3f6
ADM84CyATXzHGpcU33UgngS5Kzbtwf9XkQMNDOlSZyNdWxTVux24MOAU1FZrE440Qc8wKc9r6wb/
HTm3uDN6Mn1v+KuQ1cdRhQpqwf3YT4r3VS+d30a2Fmjdjkes/vUwWUn0xXGk56rDqMEamZr8XgWc
paqaM8yhjdbv/NDta4+cmZ9l/xcB/+shHX03SRRSbEs61YHfYHZR4QmLJF8iCZZnyrDCNzmUi6TM
7GAe0BDC52SVR5jbUocrpig02tlAYUqPungg0RangR2BVw0Zn3JbqEDQ6i5j/RhlQXzPUl0ktXxD
dbOKHRn42gkZHhYga6ulUnQzSECTpvzkJOkpvkkYtlx4I5/KewdM3qaAR59W8ZcawhESwtGPI/GG
YEQT5/OoNuLcugVegFgZGIU6iVN2+5QsnUAYB9BMPifMlo9S7MQcX/cvzvuCOdqV7uQdzAS8tp4w
lVyGKDjFOurulp83jPOG5BWFdrqgo5jw7N15TzOrhD3Xr7apRcW60yRyWTEPe2cK4yTxcsnD4NiU
QFFwQmixLB8E996Lc24vc2v67Q/d1flnnlV+Ij2j+rxlVOeRYnJYeX2m3TK1eUEbaWKNC3AmEfZX
IFeTjqjYki6iUIwBY1rreR0IE7HJGwrdse/4oCn/J2rZ6YE7lYStTeqIQlVLmAa1cpBsQlG+p4W0
Rj4p0QLoe6nBz0pmG0wQV5smo3NFYe0VrCcwbt2zQf/rv97fNt2pqcWSlmbDl1vdff5buFooUDZu
ARGfcFYrYvPcPJaSGlGQXluQqpKGVahnKMj5s+FK5IrcuOs38+lM7LWWHWXv3kfCdSrn/+mnjVTC
ROBoxU1dG4EwPeOHZfCi428NzpNhixVqETkUzOWZ+cOtI9YfNnvE2uon1ZxHqANaZ2AcaTPRol/v
7+qNV7sWeHqlC28ulYp++UzX9FelDVFWZbFMGSfuMGYAUvkQH490beuYZvR+xc/NiyMzYXBKFyOJ
wlXKywINimtT8IuG6pgrohlo/89LPRWwSHEgyxYibuj5q1Bzmb0dWJA0WvJDwyjWPpfBF8RaAWlo
EzLNZpZoLCXFryq4MwG06YlWMLOw2AYoqm3qbtTYAhOMGz8lcyFeHUt/YYGcctLqMOqOXnXe3261
z8T7+zSNyNlubDcrSYYEkQ3S5ELW0zC1zmduc4OidshE8q2wdrYKNV6jId2Zt5Og3qXTczAh9VkG
zodrOSkUz1KFXAjcin7flC7mhO94oZtxZd2u/MncCudyiZG3uA/7iR1rOVbfTCfud3I1F8cStKwR
jm/cD/Jd5gVxPUxDnnL9jJP+ss4SSqTwa5IPx6jWblSGR3Qz3/ri7hIkEys4ZWSvdWyecpGtoLmA
Y3aaEmoG3E+auDchXEGcG3oQNo3NODXU6QCjUR/BQQnxxRgEBY6XPp1Hvz2QpNNCxf0vr19Q01X3
B2fi3rFsEC3sJ/HCIr1aJ8FMkO4IINkrRW+r0tLa6pF+YSkFOiloCpuMOfYzi+2c3tPt6IlIc25L
aYBhiU4KMHz9GNOp/AUSDseBa8GnUHvEm/se6GokqjyQv7+3cY9BTcQaLcIAAZfp9O0lNATgebUI
uNBgN6HjiQgiwERcODksp4sLd92WX2AxuZ90rLCFfV5JkWRY0YcCzVoA1QsxPQhckV41yPbcbQsa
CVI+U67mkNjWKjnzuDJ0cMabfLzF8RGV3Vgas1g3N+aXOOrOQX8c2wpZtFUcnUeTFMpqrWAz7mG3
2K3oQgwtgThdzcQXq0oMEMu8lttitbuGEpIFmpRi9jQWO4ODk0DMGma+XWMP/CLujdbsfJDjwN1L
XOMh6MajdHCh27RKP6kwWL/k43X4BwaTeQjb9AJNz+Ia3nGc6AVYHKJGf0mwLtAmnhUJeZPnFZHg
9lFM3bvzEJyJdc1J/yPxumgt8BDh5rLgG1dD7YUtBjsVfXhlUYX9UWLc/7ab+xQgHJblwtH+AOSf
XfffO0Zjv8Us0ResTmejf+X5ZtaCcB6Br739ZmFreLvAX1sJEdTCguTs5DBVnDv0CeiHNMiMR4Xt
FUo1NL2e9V2Hs87cAGma0VvHJqoSXmXPf19FBrcOFCAaxsBh77FKAFS1x1+ODQ4vGkGe0+DM90jy
lCESKelu19R95uVdKtPByuFH1448jXXFxNZoUCKQPqGaWSbcHNkbIWkpfGEWA18/SGOr3p82N9U9
Xw6vyShLXGmBVLueNwTmn4jvioMGQgJeUwQOX3+IJQgsBP/PmREC2OjBuUvQRG/aoehvTp9yikcg
l6fHdZXex3HFvgXqUWlpRijjvmzCZv1FR+o4LAxStVAPHqsM0uVzMoLZHekymFtU89oDjrwX0Q3W
SorRhubUIPKyFYtOFzwDvaMIaULlcln53N50eIfVfnXrYVfl7Abrj5qY+1OuO0zSxvv5qgPWwvGV
OhN03lpUo01SKyzD/pG8FmvYeLTLZL4pPCHNcMaU7u4i6xHkPyYkORbJbSL895/SyaULlkrCgCtZ
r8QjeUw8XHPFYhBZMJu4Q9AD81hJMDu5QlVyPsiNX9jIteLyVN7Qfdl7P/VWxAHMBEV8jkTGUx0O
4BjsDdGAHjcKSaYFMypR6K1EgLxZFqo1H+ieWWP6rYs81eMn3xIC2DycxHOt+Z1hP/wQdJ0z1gPL
G7DwnatwR2MYBTjRsF9rbId5OBWjsAk6hzTUcdsAgQcwQmF+IVmF5qSuto/jbPpRveRc486lsLay
hQmTerDfGXYSoiFKPzhPhBdYLEuHz951EYVwWYaZc5F/VbOXcPjZ1NFGpdvSvHo5moCDIzjSDb4l
Dl6Yc2RZ8FICOe+Yaw0sEyhzdF/j6tmxcRclYKw6IGbcb4wOWgu4LxthJZ44+kpdszw6aYW5Tg22
SNUuDUA3yNyD9Fd4jU7n+IDYdcq0A/WMG3G9XmV9cNQaUALcm4QeMj6llnyFPVCgnfvksCV+3ZV7
H4rCdYnH6hbTOf+gPkYZFQO1m19AM9u8ovwdnSNj58js3pg5O5oA+oXXzONorPvB8r5ziD1qD3DT
LEg78rI0b15Fpu9QXOj+Bgq/eUpIrH+ZTGIWJ3bzfNBE6Ga2ZuBe+uy4uoG9KB0o8I5oGDGhtEsq
uc3Nn0adLVgKObBJjweyAP10HRQpEZdivY8WdtGXQ1k7oUQgLLr01MnNGf9am6fl5MR1sNaa+VOZ
2gPSmhW2szuI/V8vWFzCOdmpKGO94tVex66syyfmwZh24gzFXU59UIlOaqcQp1tSZn5vKA9LLkqH
V5NGtjsNQmqbE2iDCKS+X2vhkgGCUzKFnbvEOhW3ShTl3ziD9OpqRWUEMb6HC+c+klrNeICcjz1g
k9AivaieQcVo9mepvk/yBNGAgXTmPkXPvbMr8234ahvYW9tjN2Ub3FKUW5d7650L0bkOV3E0tTU6
4PCHlKxOH1Ej5bp8GB9SP9F8J+cV78loKxyiJEXwKPCDAgR56w3ZHe5s6xhDY8UzbdmcKXrl+Jfy
3eBaRvQ6jRnxPqPEhMoyIoGVC6XyW1bt4qyBo59Fmv/2cu/wDS+TjUlZxnizx+B4ILfF86ZxFE3n
eB3QO31/bRe88hwShWXJsRYbpurFhSbmABOCpSGJctzk4KGB4wmTy0ohAeXpLJPjVz3QyY6eoHYw
NfPnv1TJ/9CnU4x2Vd8lm7HD3Badd7c/QbYZeTa8lPhbMdTo6r3QRUihngWUWdpOkJ0Tm2llJJM5
Hn3rp7o2Vn4Jjo7dyGtnCKmn0FOUiR0a7S4Wp/PNMuwBr8uNkdwDAjg3VKQulaf3pWexMHGgcswW
ZIraWv9sYKzWs52clzMmkmq+PYzyRnjamPLJw5DaFccgPE+K0lAN+5q7jqN/U4r3VKLnAsswoiqR
O8IslxK/m18Ro3AS7gjwBU82pvsN3XAE58C1SGzLhxiKFcC+lSsoD/DQ8x8Q6vn0OzpdQUgCQeFj
5vZbG9x2exNtdyJ/LFgP7ATvbEJu77GO5jc8SAPPvluxeltd/tONr92t69U70ooIux3mpJMimseE
uIj0APzBCfSneEUfdoLj88GBnOk3lhQ1BXKaPc+H0q9IlnoRk4Wy/B7fXtZbgSgKNSn7c2KgZH8X
XnVUQlaMVkZ6gfnfUD9AQNLn75bN00efVkjbHuo+9+9Iuwy/Y5zumN07bEwGykcTWKyWzPgvJMN0
KM1+5msu2932N23kgvS1Ita02SC6hsBs6sqYMS4DrZe8Ol7tX2MOjJTxcWv/yGHqD/9GZLqVzXb+
XR3C4NgTAcZe/QweEucHINzFyWTnX0J8x4PqZZrUof04wX0TLsm13rIP16jThH7figY6UugC/YHh
LXWlbnM0QNRAdfAlR5h/bg8e9sRUiPL/ds/cSPkdYaq8th4nIVnRzxjD/UJxdaimDFfjnPP9KtaD
yFgwNIXQc71f2M67gtdgtn3vhjrUMo/s738UMxMbvL+ZmdNBP7GJeglVJ/fcA1bY9l7aF+j6wSAF
VR5ngaSgzS3XUZn6FFUvkykIwUh2PYzfV+K66J2mC9sTyMslFMidyyI3BEeRKWwc/Lb+GwYrTR2e
JxCgD/PNovSCApTXLa479+wAkbktFLP2aYeC0ZncixMp0jfzCajHbrm/fMVGmDOnJvtgJAL73Ptq
RZj2FE2P++k3zSWKcN9R5yNfeEMfS9TOXe9bjF5e8pApxZAKhpETO947onz8Mbien0teWotNoXzf
gGB0jNKTE9DwN2n21YgtaxBCxkytShyeJ8ZIqUL/U3ePh8bxjNo5pebxd6+OUJu89IY8nNha3/tc
hA8p9aPs3CUvSgWWjaElMnY4jxUeWaOL3nj/m8kD1LMNsKlAiSt6E5AiSE21KMr7NNaLmFlItkw8
lsyNTkXeUiXLWzGnBjbNZ5F1IhHO7sBbcWXo5sAWzh89yQkB+0N7s20gv/N0vx0AsJz7VtqJa5OC
yNt7EsSwmOu1GOI7TKqRZg97YmQK/W33ZR7ExUFefBepNE79Ux8qdGiQ7Hj1M1RsAUqXNwqLBTYC
PNjVp8quf2XYt4L226C4XqFhryrPoxFsS++9wzigBjlh0VYhY5gygYyc27Sc5JP0q9o/MPM4GY1c
L++FmV7wXA7HK8oc7q9dpexIk7f6OMWFLnSzGbtd7NucVK2c+OiPGhC87KxHSSY6SUl20CdVxib4
XPkUuxKhjtbaP8mL0x9Jbb29rao4NJLOe3xVrT1t5wnxGlp+7r8Ccf4yuqkeCODyhYMf9bohAwAe
mHZB/KL8qZayZ9W76/tjUWMQZ5Cj+n2hgbnqUjTrvf2eACqv6OzO11UAdIVNWpaSMlaabuHEiGu/
Pc++B9UfvSpNXFM3USR5dXeSKzzoFdpSjVqizbibAp4DWqy34fhW7+/NcJVjYudVGCRzEU6rMqLY
+fOSFTCuCLqfkmAptIRVJrFhCn6us9EVsiT4rt/WVTAUhYQa8GCGcJnxdp7/8i+BgV4Drp6SZtzs
7Gm1tB2BOlzR9ttPFgnLqkIxAUQDo9ROry1UOkHBkV08rioGG0g0bgOxaDpSWTl618xplniQu8VD
0a1OieORgrFEfFkv1TjmXOImZixkic9TyijPmhC810ETY3BVQKXd9EsfC18xunuRt1WF4fwyBelj
chjEc66lVif4tNPIYMw7/kfwrNTFf3jlyTzGHEWFDqU5cSsLOtj6O7w/76cCImkxOQrXSp7tf8F7
RbsPgoDFEIsUoh3n5xc+gHF2MO6T7JxwxAtqscZ1V21ouDBNJc7xojIhdsYExy3zhr0XuhWWGFLf
ZebcwA1U7zDJUYuJGIjT9I34Ai/vFV0ioLrogE5ZJzcg6axsDrvcG4MRuc31CQ/03zxkqYvLpN8r
pmFO5TMMKAgUAbgbT2OFAHld17ocqGg3boNpWhJPIRDEIgjyBj9vKL4Ah9L4nwhb+3/+T5OtTxxO
tuKx5lfnqBYU2VH40GKOAgNDcXMGo2gcmnnLJkYL/qzi8kuwIkhb84rV5RV1I3swMs9e0dslHBbS
/1y6uNRtCGamQkQM3motcW44VhV1hU9bwxR1ux83xu4uRc+O75FQvLbeL/3Fg6aMwO1ukt4B9fZL
HMlEKhj3YSOUNkitU9Q3JBX2RTWKHAXE1QyrrRCvas9x8q4RVjxNBnMgOY+4tmAjRV/MOK7R28dn
I6hSZTDkcmFIq4eOdEpmBzO5ZPpdP/F7XLoAODEUBorZ4qdAquVDVj2fIMpk3309b6FpGatyjd1a
mqICMpR5OyypobrPwOHCuhzy5DGXHrUjetfyyvIg6ORzTxHxiigbnaf6urJpZXraWT1R7zJSu646
SUDkiopCDuogm5yNuZl/PHFnJ9wcUtgmtaERkG9UirMEEpPGIXONIt3UTXO4qXIGz8UF+zOe40Me
6rQ0jytwF34Ev06HY4TVbYOuyEqf81eE0TSdq2k/UXbzarkeYvC67+lA2w4JfPV80yISnGADFlJJ
5fUpa3ZkYV5dwn6z/jur/lSHXfYT9wuNLoofe8P+cjM6GRjN9veXwPrc8EOi5Y9LL1aFB3y5GDbB
26+G4GV+xvAYCLBoTieQvabGpHOyYWbFEyqs8ZN59I3/S1JmVtVWs8JPynf96UOHmp6erX6qOWdj
Wz0fWHc3WKXejEg5nBGwRNBMaKFTiapPnrsH6wn5YjXEIIOWp1lb08MR1PGQf9SXmTFRRfaaG6mo
wJ1REQvj53NHGwCEgJFNPaim74YqyXv5PrAk4pCZ5V47/oDMv6qz8AcH38mlsM9v/euQdxKRxDCO
SPjWOnhb1SP1wWqtKNMxKS0j7v6Uct2u8+9J9kGge+P71ropjaDbhioaeg98niRw8LE0YbFLl63I
GW7RjINWYAdgNA22KJDMHR8EiIUgD//pcknPuo75ueaMZeoon1ysobB/NcDIjFQjcHlYEyEFTN7J
EI1e2br6/4C+2A0Ch/Do0LHSh+qG+zCaLt95o9UUb3cojwh2ACH5b8ZodQg6t3yF8tiUkia7b+Xa
lFSdmTThdWy7tCQ4VJy9EL9OAe/Y/XPMt0MYxNpG3QkbuE/4kUNngIob9azM7hEO658ct1BB44NA
ysdVc93XZhbsUUeYAoBaV5Z+5VXgiuxeB5ro3XH8BIwErYDUz/pE9wJW03eo43FF7jvphPhIVHiU
HMztQ+pf2GBupbMvF3ASePK64s+eZ4EyAHEB2BXwxSY3w39vAOgQVxWLY2fb0r/gRE5kuionlXPY
gt8IryxEN5aeDx9fFEYtszBnkJmehmq7r4jy7dr4jn7Udhd5ruDl5yydj9qvq07rzKfLP2M7KIqF
R8k9/ze+M2dOQO5wgunUc8xkkLUIecv1snJjuy1rYDw5IXvsQd8Im1GMhyEeKZBuGM6GggzZq1QP
fg9SeeHJXq/o0EEMdioMYcumFJB6DwL0N4vfxQXx9dfiWFJHd6P1AQyXZMMKSJureXt+O802CMfh
5/BnWFxT5TZd8b15HllnxSo9rllzB3DIBZT+M4lJo09tWT/0OREhNBvTQq7F54KQJm9B7aKZEUa+
d0d167uPiOlDKiI2CnbigYIHYhpKeXje06/tCPjrzB3sVJxzuyCfZFDip6xP/XQyAKMCIfo5XXKG
zpiCw4qcctgZhrRrfcHxHwB3klMZVBIRHcZjPqEplkt+nPcb/9ya5yYAskGJxzqILg/Dr9fuhdaz
Hkn2JkJOzQBveEnvA0LwTkOOQt+IMSterxMMiz5p5Ay05iaDTklia6QEYN9gLB6y5rZOBOqnedYb
hhPEj2gBow0UHF1sdoDHVpk33kYPUuQ5GJ0YPrBNEWuWAURAv79v4fBts4PP7OdObkmxtyB0rIGl
GT1aacSvySSwx+YgreE0EUPBx54KJM82nLHT+jYVFJbwVJpV5/q5KumG2CNtQDwj5vDXACN6fikc
NeAX2i0i6jF2O8enTNVf0TRdFjaOABX2kwQ2btf62TxzkNnGXutIj5XJ+4W0HfJqu0d+iiYV+Xyi
OBLwcm4dEL0xXE3SOWpu03M3fbbvtm0NkQSAzCLJCPWLz/G0eStFiGlB20iTilPdHqJeQ46o+3Th
XqDHp6uMtkg3QonpzpT5dhlfhwDgG+dKc/TEDCCbpiSlbVG755CMI+wf5HZoG1+6HAbMyARmNXtz
AcUrHjk8Wej6kw8Vn2L6A819K2kpHhyhJItwuTX/sBIMG6asGBtQY7lU0Rwse9qqQfu03K4SUGEB
TYTii5FblVrXnrti+UUkogtV39k7pbG/+qTijsb1jSeC70pjecKgroVpPOYRxTBTixRa+7LHlqRo
rx0UE+2Vu3LdNKDztr8iCbTRWcAaHR1k/sB2jxxzK0Y92niWMdCr8bw4N/GE6C8VEcZbkbLBS3lO
nVQvFGSsIR28eNLmoFjiBH7bxR4xLoiyRofDKqZ+w1PgxyNLt8aSSBd1gsbo8uWIMxBkLUKSzujJ
FiZuzepDVFgw0U93+tdosv24eWQ3iOdaRuYotgWWvuU/bRFkF5LhvBTPYZK3XZKeTYrJi3BBlzVi
OmexUBIiKC41jYJwsX0wEZpfZElADvSvyFqogSjpVUYo0Hz9N9ek9TSb1gO4jsK0FyfeWKcz/lB6
ZwyqW8voGNT5ut1qP693SvmBeqe/RBX2jwYVYiQlnvgjXTzSzoEnjPevGTB0GQi1N7x81jKLYrB0
3k61dMyfPJZWuZdSUhVNVTvVSt7PgWl8bxSjRm2PMHxymwMXHI/AIShkPoqKTHsIMcZPKmPFhqqj
tOe9fTOCIL020Ms4SZhYOGhWwPOPL2PwY2qVDvb4i2jFUXbOO52MAuHs/qV2+yD+uvwzkyh8wGnm
ceKcjP/Vaz20f6OlLHxYTnVEU10n74Oo4hLDun+hYnbMkYMtdYv2d7b9RKEGyaHjjsVAn2mhOb2i
s9QZa+KkL5xTnpzz94TCx99LLeX+Mn+vHL2mE+ku2dGVNUti1AILaBdcujg1S59eWXEb3AhlMuBI
tha5OmPS2WKZa8Y1lNAQd5K2BFmJoPuu+NkGOrZ40emZMaDgmRCUkm4WEMPEiqz3GaAmXrEwQRnh
+TBTuhIguAuCCakIWyEptgAu4PskJcQe8YBZ6ZoqIvtSv/tk6WCOOVLqROO8P3YiWzfJJpj80Yj6
3ZAY4nXIntmgpa81wAqc47VjMWUhERZuOSjh5gp0MsT2bJALUAtqaf48YP+KlIKQk388RmzTcmcr
K76mZ9nLImMkdNlxmhZjvOirwuh7wHnmAtYmmm0M5VFnzpgU5RA2GYXdeOarklif3mL1Si4zGjOI
TRLI1eal+NJ2LFeALYjZ/6y3EdZGMdDGPYSpFUxUco+oKTpLdF12G4rn9TLYOOwXZ9GWe4uUS3LN
D9PRjgCdLwmJUela353R5hWh6g/8R1uqf7ylAZ6/A9o0ad1Ty9qtjg45WiCAe3WG+18Lp9lNhw6C
LDuWluqp2G8w2Nf7gPMGUEKVTiBtCS4T3IDQCIJ+gv7f2O+RGw5a5WD+XXZloO9x03KeBai/dq//
Gi/eUGcZBLs1yCxddxxZ72M6zZy/a/0bHiTcLL1yqHw8CmxY88e59c0fY5S7STaAwgAzNt6gY9zU
BIU0+HhEYMiGrO/EKjQNYO3IPV6yHp1Xv48QnHj5amwBVM/VUO83T62nf+VRO5vxfPC5G3Hn0I2n
xGEwQ/2z6OzrIQP3g2ZBICdRn2l3XkxS+xwBVEryo87pB7kikdbULrb0YLN9Qpwnj4cJ0LwkBlVm
HyCNHYVLewILNWfFZgqVWtfxFT6OhGUrKn+E8CcjJjkT6FyOsv8RF2IJodrJCLUFM6/tBUjrFa0S
FxHpf9/uBWGOQSUY2sME0ZbueytCyB0qn+2nCCLeNH8JuL4lh61vbMxJLBX2fyxvzh2c9EghFs+n
9RQKGCAI9mxJn8SHj5x3t+gglPQDTyumOK1em/1p1ggPZfhPOMltKZzMOyAehF73DdL2XLpzKZpX
9NiAtbArIchAFLaZBJZdJNpdLQ4pv9sbOXQkV6tZ+W0K3nlXNrBe/mFMzJvpmaomCOd0qM03K57F
MY/Ca4GUT4p15LL26fUkKsc/TB1tbPr/LRxwd3ASWgHxrLlsNBdAE1Fh6gKMA0dwpj1clxA8HJEE
gAbovSTHRDe70u3FINcZg4frw3qhNcEw6b/pbhA6wrvvvxOMhRAhvqiba9Ys//6ykd4e9niiMPkY
dBt1nk9rV8FSsjH4t+e4zOMjPqlTEqO4yROv3udHxNdeXWtl5sGTyos+KNyEzg1A3GMfAJ2Kio+s
VtexxK8wiYpOJxd+bcTWnG+klFnezMvRi4hdLcIFyDg7TlM24mYmlllpR6qdhchpxNmefEOF8u7V
+tJ6BCnBADBfi4gQRicdRWv6e8QLhOlySdAs1m58n1H+rIJ38T7jsvC/i4V/7ubBkf1oxrbBosBp
ZMVkuW2q2Vcke+f3PRR6cR8vzA7IZKBJEzU/97eBRAUe+SC01t49TjW0d1t/eqxhIBL+xOTIs1m3
COHy7uTITmhSaQw+3PCjUGoqC3Eb7JaaA0OjFTcljPXLFh3hKDtdEBSjYL1h4s0zbVWjB4Nhh6Fh
eQpPkXIn0BKHN6QQDSniq9TSE55CaenQAT048xMm03ZNysMVt5phMcdEeBLbRaENDWXRoSt4dSGF
VikVIQEcVxkEaENQsvo9rNGyl+biKTQPsfiu1OpcFn0SNaBd6tBBOlQ+l0BzxMnr+9teoQ+un67C
gof4d4UcmhUSXr5f2GOAw42lLHByVBgJINxSGG2vhUBu4P998GwRNF/IL9ElC57IR6eMirCU46tT
Zpn4aDQNXlLzt2zTq/PAdiJ+KghqqTCKKDxyBAT2gkDEq+PRyjJvSY5DyEotV1FAQt8pHumOgV9o
ZIus8OZTiYs7AjiSH16L1JvGJ0AFYIGQU+CsTrLb287Ye9fwh0TTSr6gn86B1aBqlhjwaEAeVBGp
pxlS0H6ugBjQjXBnof21b8I6JwNY4zDF/4TAv0gEKe6fN0lmriMTLiCN09GnornGUamDJYgEknqT
3UYNe6XYXBlrK2dyP/mz5qjcmxvJdodY5/cR7FclSGmTSCLunCXmBPBlHjK2Z3KOGnhkRWhSSWhz
VVNzftToriW7nXfVStJiz7vClFkWmFuWUkJZovJ61g8bm4l0Rx30YDjwKT9DQ4DaRSkGb1KWSy7H
anbVcJM/ocgrBqS/jxRiv3mudZvle+IleIqGxFs7NX9fXMEfWocku9cbVn5KZP7r4e9hvl2SWu7r
msRkJJsIiyAXFBqkA0CMv0VmKdQDujS3yo8t725D+fUiC1iXr9DQTOyCIciyjC1QBO1QCtB0pCKs
zmx0v4evxQJ6DRpsLoe4WhuhXuYq0Dw7YfphjbRD8vxPU1KlMgdzofvIrIx02VxOi3pquZKVTRF/
T1ENSWqmrrE9SwfiEy0LWLbR/vgnkbzBSnG2hvuA9KvHhO9gjTdGbDfOb5wPegXI2lckGnO5N6dW
FYoOW4uIyJ1ncZOnPJebd28W03fF7Wt1QzrtSgTNEr25CVLfQlUT38pxOt14wWfLAuYZLM69VlUQ
mVpGGyGWI9SebazH2DyMX1gFWKd8S/nacSd1gCUIBeY1M7aB+33AajhFmjOa0iHEDjO9rxXsMxj3
wSE+KizCNVKV4WL7s4t41JVoNwGZ6esecsuSJVk7aK4z4ZeZ+pdrMjBhkTUX/MDkVpuG+MPv5w4z
cBOmHSpML3iIhHy2zn8RCa08fEtAeFCuNcF66dB0vdRnlyYQ4/DQfg5ampw6T8IZ7rFenWuhPJ2z
m5aBZoNL35l1Nddp98c5oLuohlUYkXzYWCFERAEKio2ZUmCAqwAEVLFLcJRX8fPveQ/xZGDGL2Nt
OwKtZyLb9/K+dbZl2pa9AmJawEgklMzPwmTO6+YMn9ZsPNeoPazz7jTiAY4CoqJAI8uBT+KQr5mg
lymbVMDifuo6bkC+eLhqTZYuRAPtXOxPxKQpDvI9F7URKXZwzFOhhhz6hzKnQaTSSBmdYcmxtNAd
9dyDI2pQgNF0LUoM9LYFxO7qeLju0IJXg7MtvSMJDDHqaLNnz2r7rZFd2CBfF+WwfynyBQG5n7/L
rxj/275O0u0Sg56aC5he7e5iaAD1i3vFYE9phd57HL10mxESY3Ha4SYzyQj0Aj05jcYUVrsJXwbV
q0fCnbIls5kYFHLmoYFwIoOT51acLeHQ43DTA5LmPy/cYHp0ZoZNo2rRYfrviQWAZLgM/1+TnytQ
dup9dRefCoKE6RhVqQIkxDuwkjvrenYawu9ynJ3ChjN3sVV4FVPMWpeBfrfgXWdYpZ2aXSlYPKwp
8d+cfG6gT4jtJh2qbzM3+n4o1Snew1T/X0yJsvxLo0O7RxDnFGeoWKMr/e13TIhmL2rb45XDMqzI
RJ5ITr9XxflDWaN83DXHG3hJXnZsrGxnKyET5UNKtQS/CnzWCXUhnJYnpa5tGoh0AfEJO9CjzCsN
+Bgy/8/RnY/s0aTx10T0KZFdxfB+z2uJdLd9NBfU6c3ENZ2ahUfdtSIXsvwyp4+c/3fJbVh63r1c
vw1i48GjyQ4IYstvlby5/v3j+Ejq5SX8LA4gz+J4YwCeG8C5wZdjp8XFDYgLFCMdJBh3gMHWfsop
OmNbYShZ1ldyzMipWxr93TeVCPu6ygIsiUdEP0SLNH+vCX/s0/70rQSZq2VMwwOsRrkSK3oOave9
S3G9T6fqxIdtLCUeDTfA0MCU7F982P8oc4wWK5ktR8yYHtcsO9ozqsXJA3Gij2P3g8bwkFWue1sZ
gmPR6cT7p3M7DazERsN1klw6WGLOrX0KDxlEnCwxGi/YUK5rZ9iELr4Y/ryRqKScV+RLcaIMrfK7
9EklfyTNO1fkDrfpaBeKbP7noAt1N/t1A51YsJs5QKv0ZqvkbQa0pAJeqsRvMkVRmUb4dBwZ/eC4
cELUEZNRt/DL65vJ4wKzHdGIBZuSvuqa1QAkJmU4lYGf6Zn7PhiRn6gd9iz74ghXTJ2ujhHA4cDu
oCXPMbDh00uaccChZuoAI07aXv+1r8IoOQQOSJpXvChbY5Go3uL8D7WdsQH/nUEVSY10UMhq80SU
AVsm5Z3d7ZSbEIoC8u6rzdQCV/bXL0NZkbwka4i11QrIRo7Zn21aQZO/Iy0S4+QhlXoQwlFOBW1g
oZZiKV3J//tdlewfk1VKwU+tFuSSAuJPMBHUIxTVwNfRGyRKKY1FeFewxoYANdgtNBYPaYAr1aZ9
vPh6o65gt02Ak0gJ339c+NGjzI2pk/PZTGNiW35nHZTgMAbVxRTfzpRxvAN5NriO/l7l5fMgjj70
1OaxRdTC5VAxRXMsE7QUm8+OzpKI8wsZdk0KRHYwJC/dE1Y/zvLVzysmaq+bS32VL8LgdVFe12kG
2rMTRi8aoFu6cd+BQ0Bj9KCG6fw8np7bkfeboTlHaS0SlYc1ae/RXZq16SAZZglIvEm3duYvvh2D
/qqbuYHMbgjntOg3U40IzZxiQtKrGrAYkEf5euFN0y7dMFwQmocgfqeJIAKAnKWdygiG/FYFQGA/
HEJNTsfwTCaGWSbFnd6rN5nLhQRWQTgo6tbHr0tNJg1KoYfrXKs3OB2FmLqwdyG4mV6opCPhwDVw
fkj5SeBf11k0np8/LMlPdRwB1um/IGyUIMdYAjfhffw570Ra/WZzznANbL+ilao50C+UGVTPR2cH
r7wFMeUxOfuu00UrDGPTkzWcriOsOVpI9iPJ/SvSYWd3ZpJ9NHoG8ZyybuYsx+KxLGXyIl32iuDZ
FME5k6aKebuKgfwNR9dfQEwxXPAIY/KxuaG7/Pb3iRiasEX2+YhqegnIUx8EBGLse3WNpJ8DxQv0
qc6IOzuNXTReXBmIV1J48qlp9XGbqMjj8uaZHxWE9CE6jCGSNaJt+bF5oMmhvVPTHCaeHGvblFAx
L1WjwxCinuVE4UQzlR/ZDBvLRolRdyGD1fx0t7/h7oWR9Ia7v2OthsYtcRMiFbuHz5hLUpg5RG7Z
UCMZ4MYWycPX8iTBEbnhpf5MajWaOsCAu4vCs+AT3HN9puTXKBsDZgfP9KQbAEwvWDKqyHB19WQz
ZZQ0tvSn4oCF0Gx6sahasY9hUwJdLDK/qTsvbUEUB5KG2FA1QBpPOERDSM4ks7MWhWzqiyBclrt7
GAhZVRhJ43PA3P81gwQM/zz+ic1+K+zpqZiGBvT5x0xz0kmxJqw+Lfy1hOuyPK32KXGrTIHl45el
goMjOry+3R9DjfFI/ILRTHsRo0rO99Q7LvElOmv9bfF5h70UOv50TNx0Ktg5CCCDvA2x4FRMjTHf
dkxm6bxneh+JNlEfFQKRcdxRZT8DWuGRtevf4YpXUhqazBY5Xe2oSIjafS18yo5VraWf/IqCXerr
6LZ3S2DLGYjxLLA4TM6duPJdP+d9WcMR3YVqjzQ4zAp3cgFPqRMBBHH2Rb0m7yq3FkXwME+++Kyx
bZJsNyWY6O9jI1tDpR8KkOQ5lUXE8kNJ+bI0n9GMyn0MDoFEBglH1yxb5qdccd6AwmFKuHhFkIgb
6RItBddxcgNyr9a0qyb6FHT9ogwCLlWSPy2z/VGOZd3L4wO34z1Cl6LEYOD714/hdH4qCk9RCRMH
hY022wb6uMRoUQ1bBoM8fw4RxLU/4PCCc9PgaZ/MchBCN1gjgcm+TeX/mSYz/dMKBA3QDKNU9bkG
5moLapqq1Xm2yjNqoC72z0zuTZfgP1qUteBhmI2yQmcwaVnq3ISDvu47ABT0H+EFfrCZUhrxB3br
I0+aLM6GEFFk8VxHLi25pn3ze5sMis6GiVqyTavjeNWEKo9s6vP+4NY+NaZ6/6FkBILEPpjCREjk
opchlmkMZl1aNfxjbHwQFhXt1wQmXSSMWKMfoRSDxTJjiXVewm3prwRwY/xJBKcZPdIwugtM+Fru
/oL0WYZFNpwJwbeeWgTkHSJg/3XoYjhUXrsb+1MuKuTiSzIfxxS32hPbizyqkiUbfbXOWhoZRKPU
vHH5n5/2fUVMRtabwN0Cg9CRp+OagHnaT2tcdTL7oDhhqlWKnzFBJgnY6ErDfnP3PRD4AC3Xr+Vo
n6izXmGOumPjiS0UtntbOhuAaBby1Z2EN+orgA+eaROsEt3YTfl/xBBbRS+eeoBLq0E0iM9U1VPI
XfgQbM8CoGWYS9I0Rb1TGZTSJXdOizQPg941J2ZUEiHBKVqDskvLLVLd/Ta4/ocHbKog0JcJyze6
4eaB8SbzJN6r90aIZgNZr9S4Uv9GGa9Bo2JMDtZmdV7iEjOO9gg55aht0yZaPWOAqj8BJoaNS2ac
VxwHOzpjiMk/3ZCThQdPSpoCctEw0M0LKis9lP48Ikl0ZwwtVLXJqc/hzu1iibtYEGAztS/NBFKm
YiCER0YCLb8HXVG3XGkgDlbPRZlqv9il/7GnYmh/R6ydz6fHM06HgrfpkRLKqtG1cPJJ8FmDsUAh
qROS6UckN93qhBcHUgMF4MG2F/9eOKmMU/dq1Q0XZVf/8LHX6+hpwZ652peHX5kf5dMrikQJjaSR
dDXOcw1e/pbElnU+zvqyBO0CaKgjHds3OXDnw6mXR/RilqNGUKYFYfCpr5gaNFqFE8GfccmTnUdU
DQxHPBio+ZNzXoek3MAkiv/jSDbe0D0YWVGQDLF80fSovz+/7du1hd8Mnhes4G0qrkHlHGIEwWjt
eP8NmQdO/VSwBnQy4Lf9rOwSyRnvddc/yRuFl1cRNA031DHK4J/WQVb6Jnn21VSMDpqCsSNb6KSz
uJX//uG8FV6H76cgbEPRqKJE+qcAAWyoDjo5b4w+xBrd/slt6aWX04objp+tRdOAPakARXkwD3vH
09lWppTX9qn1mxxL5iNMPm/bKLEHyqKqqXj6GZJ1oQfHJidlPBJZHu27SYdk39s0GNi5b88/3Jpn
UerwiGA7eIEftAno+KiL8aWjWs3n2E2o/zEt6ToTypYRMVnchzRde8i2fKUZrgCgcrFzFljR32Ys
ZL9oHAh98nTohQAHQBTQAvbE+R8HSDQ2r0V88OosAjvH2sjjz9/H8mV3MLyUHRgmlXjlkjTaSQfV
t7VQqJNPBPtLXNqGoWjdj2+O2WO0hiCQAYjJFgRunLXapf00OEQ4fNvyPtItj5dSUZjK85iLxJzX
QeR+ymF0C6UmFc/mw4x64IiLqPpzZmpAAQK2MkqPf8yMEoma9f31AHqsiqTMIDZq+CsbmJ0YI3GU
L8YWDEn2DD7JYPwMe52xMdQeLjGQcSmFEFnqpphyMyvUE1yYWW2oG6fItivo0PNT24fGSpx3mwJ4
q9QLQg2OP/wVVXK+L6biKMR6/BScsOwAvG3TlnG1mRPrJVUmAi547jeOQswMkKnJoWPHyWV6eRwz
xyT9bqBm4W2f/GEuSCmp37cVHDNTILm4iesNPoRlV1hpVlUJVJeJf3VN2379EmbRtjGqc+Eo2CyK
1N9b5BZTbyqU6Huxd/c2647mtKcUm+hM4zAC8ZZPIOqcOGYUEoADQ3cuatkh4uGyxyKWwCq5jUn+
YGAGqWtTBmcYBVfv5QNI9F7TkdHgi8xWPLTRJNmiIs5TYiNtjzmHZ/S/xtmZFTv1IFeUjikdUBYC
VerC6IZ15S7pxrtl063eRDqO72+bR103itPnlsIJSQO8SolVahWgoYFG4XzCgaVid2GI+WPR9UR8
Zb9OeqkBc+yIhdjWXy2B/cD2vbsHdxn87I+O0BsK3L6Z03mvM305oSiDq1IdzqUTDLsjrQrNb8xd
oln6n2sA2fbb+Pv1dt53D6SN/G7zAgUMZv29NI+CHTAVCa14l23jSSWi80VqXzCuyce42ddicOPL
INlzM5AT1On+e3+tK7aWSnVFauNfULjm4YnXGepqq1jx+PHiHhyJBPNFPtpzowFJMm9kH7vhqmqd
Cej8Hkf6IYLEogrtBs2iw7M7PEpFRYmPFEmxCNmgqnIgk5WXggJdpYJOF0tV1g2zgVUQEfuBCUik
fWsj0sP+aHH1WTjZ4NuW+mXuc2f0pc6WvrvdqLmN5z9JKtCBOEUApuJCdphI6rskcmLl5iT4TTCT
Pgr/YYdPMFwwL7Z2oTvaKEbTfPJV9CDM7xotIDtze++ed5pK5L6FBElwA6PD1HgSUL7ti9dX90Ea
9LDVU28X9rhEEFhUbb2mXcS+44LCFBcUeUsW2D3/LbwnXrSW80WZLYqv5RUdm36G51Vsc6cOS/fZ
1zXRs6648SJ+MYnBhKtkKj27Yjp4spfcbod2aTtxLqt53sjM5EYLv0wU7C2dVx+cwxP42zkP/49I
dvyC0JzJZqrXpJX7UqecuuEzvdxYf1N/WEaGUUrccUZdAgvARujozXZSZNOTcT1h/ZfAlFmG/qjX
Bok6/AeKt89bKWEJFBNU/8jnssRNlUxG7ZttgQewZl8XfCaKynhzEhvJ2yj1nAcDksV7ifNQLajx
9DRNrGjlhJPtL14Q6edPrRKvTdRJSDivEeMHf5aW0Kmdv8fUJqLZDGlN20403gx2nInjhKBQJ61E
p1I/Cl+Zn4qpDQPDiWWKh+6EkuQioroMvXwrixAUPd2ShAcFz+y1SCOVquZXZ8OsSAZhk0j9h5OP
iFiWL+1+5WBsZ/kkDyqrG0W/c5+s0Zpsx7Mbi4wcQXjfVdMfvKk4IGWxgLm1Ofv7vPHSmGd5l+cJ
CqukrgangEYgqcYUuWg8Ni2OqVg7A9z/1JCzKpGfLKx9Hma2XxFuPiHKiYjBgHFpaP+pNln8JYK4
A5m6xaGng71NXX633VfVsRhZXyw326s1mAaaIPYUQdtKgncfS9Kb54ft7yyLjMCKAXSoGRqwN9f9
70LGuGdEU4zOhoH+ETutXqzXhsrclId5zV5QKxoFp9trTIsGhUDn4UI/+dIpPWr35OtI783/6Njh
4ZBpcRzDBNe8DwGMHct+0YMEFN20ZM7I6GsYVC0s9RSeUdCQpLyaqIX+qSJ/AUBy/lOXBb5RGYkB
qJyTKfGdYHwZhUZyUl3Frwy6cMLMFqVU85AOgcxAmXXWN+AFQ2ilqgpPYidz8+ROiLv0rMUiWUOK
JuiXsmToeX+t7U+3HwnIfjylrxDBQ3H7oke6gVn8yDuAyk8ii/8Ch7/PlJ64Jzfr9Ccpta57LkVV
S5LPsyGjMHdhS2CKqRG+osKt87ji+Jj9B/CFz/nbDeO0vx+HZmIvWbYaY9rMIEOdx4qW7X6E2LZ+
6SsMRzMOFde2rP09Ax9kZX++lrZx3hP0wNu1L/2+48r+7qGBdjOiQys97gvqhcKkwM2sovYeWXhF
CsFNwqw61lke3BieAzd7rmyo5a6hHHOydQQ8GcPCrQEWEKjg0dyKGRQUAVvk2acpkw0wDksOKxm6
R8oC6wk7flHQ5yMeaAZLi0ir3xHgC5sWafj4wzaBHAAC9SrhOjlcAHBGElLg5QaJXs4wIl4gmY45
k0krlUVxV4FuH49Mqpx/LYLwijIEpqCMNeObwC2sbINmTljddv82uknXVTj2jzcYZFZKEMh76qQw
7peA7jm8XCbiZNs7pInjkENK6APxY+TMHFZ4JFIHbuzEU5a4I38i+JTXTDVLg79edxiti+ASeO7v
ZKze0OeIEnirlJnEVJ4lIso/wRKEVSuWOsxVebl91p5mthvgdH6kHd4f1LaOayBE7tHcaWDFjlrz
dqkNBy3YCLsjn4BrSWUQmZsWPzpwN9KfEXAfRfxNh2Lx7sk/q6j1kYKa9l8+3iZJinpiTYEpUExt
0NBO020qkbr9OS6m2LKvxPY9YYbSCYftTr0384QeVp6FSJcdKpMbSdIw/DxUbm1bZ/rXUbHOY9pf
0LoKxmzUS/Cj7nQHsrMpDa/CCZoUEvlU1ZinLO9PE66H2xBbbdJz9PiCFkBv0Cn6sd587e/kog9X
3cH2paZWn9S2lAOEfimQPU0vE0cjADXheaPOg6nG9y6UCxA8coUKFXyP+2eXm1Wk7mgQ6m144aan
2exBPsV9Spekale2+qome71rfR5l+k83HJPa8NkNhsNhh7oQCkTidCeBbe7gTCdHL7CWu0Gz2sZO
QDNlX4tLHhl5w3IAXNJtqRU2Nq9wOTHHtNmDjkeBk+ThNYECcPns09ECKxvNK/Kjm3y447kj2gwm
TaUur8A2PuW7vlQrEH+nqRAmQd5JgdkmYnOb56mfcJ3zGSYPy9NzLMCy4280j4H/3bi4fNDS5nyq
XHrb7jZ/BWpbd7B3nfW53NXqlgo3uh6psqmso4PqfBZ+M6AH1knO33shgtpNkcDGWgEPRp1FmGYj
40aIDi1/2wDxMyBixs2ZO1120yer5CDvN2Zr8nsa7gTDTvATB5vsONlT592YxPa1Qzvf11wzjrHM
oIUolrPdSyS/8AB7wkIGmCW3Ys5EWkapOy62+GwsnWC4UH0pxy4577etrxPOx4QkobGThyTPhReo
ilcoc8l2oY/Y6wN+VKOW7lAKS1kcEXGSruA7hQpDwluCEzGlHxKY3fYHLzUddEcdAJE03W48gVrq
u/pYWXD2J1lKd+dS6eUR3CoQ2+Go0GzmTqSBOZMYfavlGcPUIwjoX7QIQtFDi3UkwR6p27BflSFr
W6JAkZA/SxKZTbXkzSi/wAysNMNDncKkasjYJgVRkCNgkawR/+eli+0zH26jjvjdqGBqJlJVlfnE
jJy3hB4Yw9Xq2qM/YcFkQ52uDlC60Yuga8q+9EAuYBB/n6KDBw9KGos+RkCVoHcsK6oCIiyHkOP4
MT5u4hIs1yaQIig47HhOaeH5O1i3o4jrsKYYUT05eIGN8lriMLaZJ7UcMitRe6Z6nHDwEbEmTJyJ
Kev9mkkKqciJimpEtC7hZSmPZLf61KR6+0DCzBW1IAwj1syJTVHPzUcc27qtT0uxtHh4IGVUNXin
fVRyZSvXTSM/uwdvjjD/iN3mG556iDcagZI7oqre5O+feZsl9p8qsIKuaiMF9WH9XNTvcummUcPv
eYOhnzRQsRMUZzYfb3120MNbiAJe5Ucb2wM8ru2cbJRTZZsCxR8HtWsQd+g14OVpjE4oQ48CgPNH
7taXZF+JrYJWveF9n2Hs9pScjT5ag43/2U5oujilv2AtK4GYrtkf2WqTTxLro9dhB8/zrUgXuxH4
TLpG6BpN8tcDxRVcNl2LOVLNsq5BVBGogqWQu8ytW6RyHAqmm4Ne0yH4BGhJiUJPBvB8baLEA67p
7skGgIxxDk0nMLczYkSGHc27FMkz/pmRO4va1LBXAcsOtQayeaSdE2Z7G4h4rdoqTujLw6KRe7Gl
l6vUDu41U13qDkd9IXgKRsBlyJOd+cgd9Hqtip27hiBadGD6qwIzCH3xO8KNvMsiw1QWuMqn7Lu1
53UCFvjRFlDyefeI0v+5mexX6KZSZ5ZEo647NuYk4/ByY7JDFpQYBi3f3dI2OLH8Kg/4Dn7+7hng
jj8t4LaY2//XQhKtuygjFE97aYdJQ5cpQX74rDGYD42sdwaCgaFw9vNIY7ynoCjmRRH4earO4X3t
Kcr/lNFHHL386ACk+uScPI5JIRcjDqoZ8DpdnxnVV08mpZ//Rx2/Er8B1FPy7JikaXERNGDPMVzg
nHk74/v5VQPZfX4KCzPth+7JKEyXa/cYUhHEpxIOVZRk7wJX5GO9RBK8h9lMwM/1GEP19fW1oXOb
PHrwpnrAJ0YaLbCr7MHmEGme++cJpFWGSqlLxqtZ8arJGmEOqsAtGSjiLqeMzrQ9evfzyd9DKRQS
z0dK0P7KLTUcT7kM3wILrfziqp1k6n08NmmGeTEHuJKAp8MruEfgw6rqRJRCeoconNC07MxVMpEY
62/c3f+i9ERt5ja9Prfbf+AFNT2UKmeddI1HeHgn34bONsDWbZjBnmJJ5Vkm22gwM9kz2VYj1aWp
WxRfeLamYoAN7woYj4X8m8VNY8Ep2N4QSvNn/5bPux7iAROGO2fGW+2w79/yq3+w7lXrnrfkan1+
Y9QKYJY9VjqJNT+p6w5cPBU8WkKdOX7CEGyP6aEXYkzrRvS8az/mZFd72RPP4J0FMVnxMbKZaAXW
IaiT5EQBtY1eOzIUrqwuDoPhab4zMRxsGu4ST95mnDy4bf7Hc1ATdeGuk+WOEMnKriikUBhbZaXE
t04J9svQC6vEmO8+ENPfCPXR/UHvieiU77+V9ehgAvp9FYB8BiRZyGD2qXwastDpU6PgUBh8LbER
lWw+IpTXe4A8Dwgda3TrVct2H1pLjgvbzItFtKH1xk/A4L+z3inrlIgh5NkI+wnO1L1s0+7nptpO
G/Z7FZ6ExUgo/BoGlpD5d35nbkp3GjI1bOxkaGzeq8sySL2GuiBJ3IXY2zuoJCRoHIPKzZ5GE7Jx
jjTzA5HvAXJb2gh3wwt1tkECqXNPUzfFQxqrVVq3hLQzzbUG24jUSNIXd0VmJ90e5h4q1xTQhXKY
nOt1OvhLWf0DPjmxMQkSr1v9q7hYXiijNpppQtIwWOqV9wwqC5m+N/EBcb1clKZnl60FsVN4K8uw
XWfNRAY0cpk2kM/+pXkwyjlR9SzllcCO70wEpI8aiaJJkt3JlX+MxLj5X3Z9pDTpepL7ciXsEpNZ
jKP7D/+sw5e7qUyMr2JL7q620+Zb5SZHX4RrAkqez3m+Ad9S4/7+8W8a/yOmsMInoZiqPA9DqAuC
L0+wCtkxDBRVVH9WmjPTcntYM9UZZYvGyYeZgdTh4r9WaCpgPnHMP7xrY5mXoRrpV2cGFOgESvlp
m71NPHZ+xjuaWTqh4JALpErgBpyztRUbyIyYq7NjhAWUz6idIysUgW5rU7PD3XGT0VbkhE53ZXmv
nHhPQ3m3nYvDdLG9XT/Wo71R2tn32iydUIIl+zUlw+X+ukOveD2Z3UR9M932ml87ZSiCg1LDqVh0
DP0Y/AlElurYBSJK5NrZXXCFXoYoL4w/dg+x8ecUNWwraJfvM7qFVpASQTvU5/2YyvOQtpMeyL/x
IVqLczhnxs6E8GqV71FPL1m+u/6+C6ClfGExYbGagPO3bf6BqMTASf9c0uSB8VwvGbAwYXAQXTJh
Oe0fAY4FwmzY1OB1bpXrZ7DL6t8Mz8slLiMCnFIOEqvcBdtf7OaZgU3jJ038mSUvSz4fh9rTJDh1
SskbuGiEKAUW5NFZUZK98EIrO3xDo4WpUbeUl9p2dH4Um4Z81a0qDoT3RgG/P1JGvoqzTizk7Z/I
mgfO/ptQaa7fFDNhha6KCfehwPDpq1kS7rpxPpk+JrxMnhFtJAKI0ctcbiRUwUiSLM6kmZPdM5sQ
Hf5u4OKYb1nl/4uKV4/XlgAmhD5ZRPzVIK/ioTj3wHzcxQRmqnxA4iHDDeQnEIFm0QVjVqCcX97P
i5Eu6HQO3a3ZBrxcfEH7HYqSBFO5BFkX6WcYVsNqSVxAu/zTZ5n5fLWXZWDPkP0ShZRsvnFuTUzE
1vfN5iI6bvnz22CGf6fiN1RczvojkebgKtJhkSwQ5qFfa5IYN+PhWL57AOcr7/ccucQzhqhEFXs6
cTHdjBraiERGAZy7s0PzOE80361woFNCErG0CHyL6zZQJcU4UwGacizZSjFThyzijf8A+2SMwYDd
f6+2rZNfBvMnZnbRlo2uu7grV9FBhXQAdFgToYA/6RosGyyQ8mdOqVSAVyCBUep+lej93ljvw6GT
t1Y1/XL/FxxPwiAXjvZ1vR+PysoxQZQr9Isv2bQ0pcqTxHXMG8mGgyBnkaOrGjR1s8OSgTD3GZaU
EqjoWbu+YmzcgEsfg52j71V22s7iHxq6VmgSxGkud1WbGRIvi6u6HSVokPuCTh36+79uKJ/VdXpC
B/thQkpjKLFQ3FaNWLyb99Ohy2C8ykrY4XF3FL87zZzutmNKkXInbNqhfBiDCeKGYcQNjnPkse4f
78396Hwi3XrB3gZCLogds0lEI/kEPEzfkJllZw7AZK/G383mP6AdBTLjlStcBOCWmdw1/nZf8GyC
EzezfiAdt4WIAD06rfZoEOfGznvLjraRgZHDHuRktBuVitg6OQ9fpXY4zGHUHUbWZM9oI+JqRtkq
OtovbxHGB1C0Y2BbP2OwYunmdyn1KGcRiGykQPo4hzS2zxCddYbSqKTQIZwTO+wztjNDm7co8i++
4gSYpcIdHW3epX6qJyXTTP0YqXYv9/r0W/R72fL9kNN2njiCKLpqklAiLpLv3PH2UC+rqhszL8RZ
zN9QvPDNUdOFhCSiNnG+sWVHmriHLLwM9YGJHw+Wj1gMsOtWn0GgP7RrwCQCdcTuA8mZaorS5ut/
qPyOKOGYq9Ai4KkrFXj7GIs7Oo9uc7jkLhXCKoDtkEOwNeWKhVQ7r9pGgiFIvlx0SVz33WKn9mzn
GGn8RELiRhyGfoTalXRtZvxnzemrwKSF5Bi9BODgYSe+hpHvfxx8omlf4lc3QMl8ouMqmrXjBhsr
DyWlnVfaSXlLX14K6ayiNoplemWGKYUyeVMvaHhG7tptgzEmgm5rT2J541KRyFf0XHT0WCEsT43W
kdgDq+d6xP8nIlOWXnlppFI5GNMHHqW4+/9uPMV+igeNn+BeclfEjSw0PwsO+PAyVrfkPCt+ps6E
ZhhchzKScPK2qgG5cido20iO4yrvlc9bC3Ra+g1nBRhfYdtdoM3tHCSgDinaQZ1sCaZJMEXNe9Ev
LcYdzZ47hUTS8yqcZaq9v+bvYnTcEc+tdBJBrDZbh4P1U1xJTjyCgJdW6IJQcZJvp4u7SdPuCqPC
0diUwUf1VQ3q/my8MyqwW+lvWP7SwwGiHIXx7+dk5XZYe9HXB7x5wWcODNgjfbILTNHGaafT7e6r
Ap8ula+wEOSEgRBZIRGGKKsgOWTKWFy+xzJqhauBpqShCpXLpj/HKv6IXqKYZNm9cbuWbMA1IU3Q
5hvXYeixCpjvEAKrHg70lo/bfwVpY0xoiWji0j9lvpiWYisSpdRvI+OzbAOYZbr5e64iXi3syawp
ilnBXHJlOpZMD6mkSNkR8Res3Zo4DMruQv0PafjVAZyHcf8brLY50YgFamGR+uXdwpt/0vq1wHQr
xggPqD1nG5Hy16OLK1uRaG9cuOULWaWPpllm7DlU9TsRw9TbtuI2O1RgIGSwPmwKADRG13iyD6co
0KKDE98VtggZg++gIqcZ2UK9Sa/EmT101WQZcFjB6p5LN6x/lrdU2VXoePrT7xuv2kS7SOqpFeCs
q47H4rbv9FuZ0JjM8oFCPbWZkETHHv7lps6lk0GsJXqO48aBX8p6EY1S2ND4JBA/OP8ZN+O91RJ9
Jxa3/93FpeaCLkvYOpqCMEoSYE2AWR4HvWFKRECmqLA6jx+etkeF7Zc/9LEa3iepxG7egwgF4tBZ
QeY4ibPSGyQ3mKGn9OvdLQW2qAJMhjhLwrYJfxuC8IQ95AOX82s6x/uIxz1fNr10Bs9wAAHQBzG8
lilQwGQcu1bNlMElRHC9rJzypOxc59Qozoa029C1yujpFirdqDUSE+ssHqmTan551Bvlxh7p4xxt
84VFS2WKhv+aiB+0naRUNS4I0pJPVJEZOMYpgHLtdvbdeVMy56SH+8uK87MGFDup8LPU/KAnKPoB
8CPfAemvZXxoxlvyWWwX8qOySmzYiuig638AietQHmo8ahp+aDXf45+k/Xc507I9sx0h2G8CjqTf
zjFL0tfu17AG5TzJaWcADtSkANrsLG9ASIr9jxYzknSDmTyV8BF3+bkF58yxF3pRTXxpE6uYZhS1
q0XcYtDEI62LALBO2rukuvR0mafll1SP6/SJBpNCXGLZ7yMaqSWrhnCzaS1MWTkHUgYMLNImi+bz
9N+71EYa3VosNc/RkyV+aYIYWjta5NkBY+PVwbS69O1Ov6ZKeQcK4cHAQA88L/PRLkWi9ABG8KdH
7C2N3trxEl44hL/Hcsk2SwCpHi3ND87aNvj23LTUiE+r+p7KgCpqz5ldql9kWQqsfjqIYo8919ft
fAH2XY//3JzdhuHuu7C9QwGZf/r3us01yd3w5SX8KkHw4mlhSdsBvnk0roIgRYNNuKZO706ipkF6
tRgtyRGGSNgcDdo8PgJgJAvLDJkYK9seMDDID55qPB4qxFzykllMROI2CcrWoUJKa1wWpsPXiZXP
r9rYoGYkBlwxJawDxjBVbdanXVtWaJ3/AH9S2hOCdhDy/VEdwi97bAz+b6sdcUUYnJlaVoI1SC7a
AWeokdTvuIc0B65cAfr3j8tj5NrvT0BLsDBJmHKqAqmbrGR4nXt0iWIIzSofdwF7caNWuBRJA4k5
vvS24BUYTRNbPXloAYp22i3VvfajMNPvUKhBFBatqW6+Z0jL40ejDJGABuF1RJi3EXzgJtm0koO3
pKsZxEEty1knXamMqwkbRV7eZOPeQ+/Y7vtvMEA7SsihCya1Nr10x3Sq3hRPY8cG60pw51Uef92i
4XPkRSbgWQcJ3UiGQtm4wtF7Q3rrsUB6UeClrFWX3hOjeTQe8oPxABZu66lq+WTH8WrUpbCo1qT/
mmH3ch9tj9oTj/5L6gZwk2op/mw+XV1bTS0SNvYG0s2dinbba4U5wu/rJs1adG8vKYUvtUN5qs88
qyAZk5l4iBhMyVejeaKUbiclf8OZbEzTpB/h/QdtihCs4L+mWhfHm/uz56zgAu0hkV3J+GChfkpn
gl6oHlOAvvUcoLjIiZFVNUbmocdBecN6L8FNGyW1bDFAtLsmXTZtDc5pJrwl6HeLA2dIrz5Mszx6
E0iEKWveujA2BMbzrMLNs63SgdnC7U2uouiyOiVtezL2d+dlor1P4x/ooXPu7s+FcBU05e4PN6xb
5aCGPDkxF0WRNEqzQT8OdZj1seOUmQcvImHqBI///23ObFt78X+4no3nYllxwAAl+S0YYd2Xh3zi
cVY7ctjZZnXND6x+DWXQqrIBCid3yXYcKXkEg0Am5JjXWO3y064etvZjemZB/baLGDUabFnmlceC
2KAk9TVyRvOnP/0CKZZNUdxmP9/oGxE4++jvrAUdOtezNmH6PT5fatANXkfvVUcoycEue8WflJHU
8a8xWhYWIzE9xxis0Y/XVFNpaj+GVbEPdzPAVFXc322VNISeoQ9BzFYxF6NYBj3HzwQ+WgA8sp0N
sOm1v3rffeH3P/yAguBErjjl0T6kJYhEA0lVZZZJD+MeJAy1+TtGlXO5kH8GSAtLlBeO8tSBVzS+
dqqZo4iHlEdl4xwUtdHIOFLr9r7BtNKrQUWObHnPyDsCGtdsk7SECcs4VDiJEOu5AfItf5ZswVai
yDveWOfCfIXXGKG7GmzJCrV7SoZ/PpYHyvXSWV+9LFnfn0cdHYaQYLTYRxazazp3hFm2EMwVc58b
+UD3/ZHxL3quc5kWMhwrBWdYNt4NBNvjNF8q0ZZ3HRstxI2ZciyaQ/dSobHYRzXxivBLSUhWjKbu
yVBRZhEdmsnkEUZI7d3WeUcjawC9ZKVL8boR8DzFhKUqfHFvybqRflTyJtEMGOk+OYgzvfMVm16V
RGya7sdIlea9uTfE7rXjDhCSQz5lVKxV/P29jJTm8oDrMPt6gy1oVrLyq/cmLI9/8pCwX401cKZX
mVU8MxeTPJCNbbCDntQTUHwcZeCC1Nd2x+XO1ntvJt8cEuOooe4Ey7AgaK0psr2xE4OGyoHMC4G0
xHsANVW2xlk+DfA++qFWRKs/UB8qJp1I5X1Lp2n17fl6BCEvlfuMHVsWtGcytzdZ2JTVAclgIJGw
2zM26fjF7BhMjwEDlpPzWHdkU9ei2Ytvtdg09+EthENq0LPB1j23Pq+RmF+zPvOd+qBhwSnXHi9R
S0etzT0a8Fo+GVO+mYOXBvk0SL/uHl1cxXZRLSdvR2TSBdijXNqOQia/am8rH5afkeCGt6xFY287
f/ykoSOiE3XfJvVYBJ/Gm5hrmF9J3RY0L0kxtYzWXuohQ03AS+nitJ/7lhFcluu+8AgFSw1ZMMv7
S2qZ6JPW9DnG68+uKcHeucQAv3BijgGwY5om19VybVQkOI26kcMewv/qKthRcLDa3LJgf3XhNHtn
P0X2kPoQV0Y3AojnVkBixFCxwJxPOqKkcYi7efDNlMSz2/qwn7XX2EkYG36rBHnrsyC0Gb5S7u5W
ogI8YSKSunR0JmYWZfr/t9oqGLh4E1cSlTHV6/tfPnGg2jaVfXsEnqmzjuB9lWE6p4NukR5uZ0kR
J/NtgpXEb4Of97BgSIXKALceyfwlsEeX/C//B/PeGNdXVfVAlg45Jj9Ho5vBcFWAwUmYckekUV3r
kRsLQ4+twJnHo34qRPgFgV+2MOGTmn8zj0eaAYHXmw8G6kCxjbhUPwY9nUpKoa+4EmJbJyK/Bc1a
59bKLhsD0LRG2KN8kae7asDWpU7CTqdHktkrYHQL6IjZrV5Wu/U5P6KZZwwYVPOYbcozF4AcWSHS
ljyX4rcC9WE3WNuFZ7lv0AwptVNhYFescLr66czHILSGfNbKSOHxzY4zC2MoIPhpRHx6Dcacf2jm
wp7glFCdf3S5yZS01T+RtClnyLeIw9FDMG9mROrmvHWmlMXNAiVw/6O6mD14zIdvQIl2M5OkGR+H
dYGWHylZtdKNGkBfREQHEV40NqoIKCtcN6B4ge0S8dGHcP02MDnuSPNel6u3mbP9DiM+kmJfyDq6
YaLMBM4w7JwSiUkk4Vw4Oo2V/nGOMJnOitjJGPx8LbOuYQGE/MKbrnlGcOZ/QRH5vkbYxHF6B9d7
MbspDKM65RgNzATTqy0ps8WrdGHCaUF7q6EJqR0HAKhoR1zLmfiYsCyt0Wg55ZL5v6kL3LRrkhIm
Q/PVZVBAOFZ7GLHCxNmoemSgYtBvf7E/JS1zvvF3iMzB2LntNQNxm1QPATag83rEBFIuBSuO5OP/
vSR9jhjehOs8ZS6CYcfTPjWrXNPm8D4eUE4ob163Os/njlkh+QUjhDFeuxEXNHgKysMiIi4RoH2/
EjtqdqgcapWzR67obZdsggnGdBd5pflkrN+h2VUbta7/+jtIHbiOcybORKtlG9bwDEqO0hnlGIXL
b0HgzAVfFJP2ZOLfQ5Ed345Ko5QxyH4xHYAlDM+jWeZJnAPFRVhP1lghtaHjhsDTG4Jh1xw5fy91
LJt5U4NOen39ACrHFBvj8DtsHXusOAqqw9YAv5oltDWLHxlVpYnSiTgqrBbfolqDYaTRfElJcqzI
00yscI51ITu1Kviq2pK3j0T/XPhn56A4GBrVv9D2NxVg31lu71dkLGQhFYSojE0cn9DwQj81bAEh
GW7NZBQfzf3sFpOGsvsJ2nrMZ8WjnjHKF2hAcymMAjWbSibAkGv3zMQyJDlX/bcr89E/ty6duXEx
XbfMZvZFiFSTmLwF0ccIixDJTa4Y7scNIA6Fe5/ijHT+OGQa1sgIEpr5dJIFBQAijZ5ai0GZn+Cz
pecGKO4XYWf6k0SWUIVFWbwAuyGQDKZ1BU3TQYgGCh/YwgGp4uHPP3/78/Hc3m0T54HrEC7sCqa9
UuVLKlUR4v/Sv0iosrLlKUxwW5focphNjOm0iB7Ne78TcJ8OijGc1nrgcA0enj1lnxfC9PfwxiSW
REn6phD1iS/+4IdDVG/UI4zDP81szpN0NWpSBZYU8dGh70QQYVtbLYVIDbnF2VFg4BdPe8V734hq
XNQNZjx4MppoLcuItZXPXMPWTchXX4DAYCJ6yErz9ypvNWePXJbQQYuGSawvPiGzLnqok5UbcDF+
4w/qNjKR/9nxXC1FF4NueVqLMqqR7wL9yyz+uwdLKQTd8ehV8wAMKUQO0WhXxzOFgV45Zu+whoAP
862FmEQTkoRNcwvGQP0gkBwNSbfjArrLbMnvNSGFX1ArTQaRk096o9VjKWAsaNfvPAnPv3hZiUQV
54OJKTZbL/xp78NKnvS3+ON8bVRyVMPg4dnLKt5U388tjRBxYgCng7uJrOTwmIF5Jud1h2wNmpmE
DWcTyBBoIwsmvmsHp3Gr6DM0l4RCF4eMGbEmAVnaySxEeE1KB2DYD+a1Fnpu1mSEVlwHeZAdLfYC
LrxK75y4m5ZRXEDvEyTisPgxyJLidXLeIPETg/1cJOHTCJVOX3VHyCh+q0Fb6YX7kBGLB6Mhktho
atd16i70gdMdXJmawj0fR3Xl4gcQWAT2Ew8bcPB0Qv2dGWSeW6ZGZeDfifJ7XLKcyQumqkouL7dt
P9qobe4QV9E4AOYziiXAiOE0IYLKhVIc4sQDSMUvDMNBI8tx1YTHbIJMZhTXAXhRGKTsmmSMLCOQ
IQbT7BiWD0+AuN6Jvy896GcnMgKuoyNCHyqeqADhJMrixSWvdgfs8dSzP3egilsP7WkPADWzL+wK
3rM/VB2J/76eFR2QppoR3mrRv2Z366qdMGko8defjXDOgI1qirriVq61iFFeXzuOocg0VRbU4ySN
Hsfb0gttBy6VXoUnPwYOYn2d4czmuusX8u1b2eNj7ft8u4tUvPf1P2KLGS9XuZAKhGnvRunpvj9R
zJKexJn1U/h2kop1yt+/BT35M47KtQa83N+h/1G/5dMLylTEV8RBt21FdicVbbYHJikkS8PzDaBC
twBmOkBnYty0fXBjWRfKi5NFGTzgteFRsRCUgP/P8Thu8utQibI0Wmb8PD8ir6/cL2CBUga2tIsu
zRqJOhwGIbfvjuyLxyoF+SLiP+u2FPQ9ThhFERyToDUnWfcD7lyBDta68BVqRaF4O6oy9b6qwSqy
NEHJjE50aq/9b6yMFJvCeyK5F22gE1fn8Ot1212p5VOyGFhgLPEQFzG2r1rfPNzPo9J9BOaf86A2
md9O079RhhQtr4lHrAc2YpLL/XYT9HD2u13noo8nWriiOUz4ngKOWG4huX25jLB4uBjkS2rLENAm
hsN0xW6jeerZ7mCKalvpPLsNjqNeW/+49kI2cGJZuz8bi3jq/CxcdXECSu2MVLhlDIAeeu3bO6QB
b/yeU/SDClhCE7pX17T2V2nnUSeaqxlE15Xg3yr9nYnN6NWGPhXuFTFHruCOQtbDyZc/ssuBXGaf
iKpCWAkz7TH0iiYEHEGFfFxgJZ0OK3Ww0k64+n4ITeTTOW7NF/JjgU6ANMbb8pbWHspAQ43Ipt57
raJuCJC4Idjn/nqbSBFt1QsXS7QgIH3jSeRxEIgoaYyg6Xy2xYNLmvDw0MqZhySlbT/HhHJXRk4u
qbS9Qz3KtMdvZ/M0o9Lf2YS6oEMm9xrB/0xC1rqTCTLhEm+B7wCqy1PSOMhx1Ysin07v6/7RrS72
smoz+di3BTprIct8lsN80PoQWOZQ1ItM9Eqa9Yfp7Dy88GPu50T3klP6pRYXaHcySZfqp0XnqFzO
WmG//hHEcq6jNbGi7twEsfHF4AVxRA/OoowgMXuakWk7rVzHSAu5FnrdTv58OMt+a2pRijv71MB5
Mdn33l7CtQmoZowMqo5+Y0h371auArJZWP1eOSNT0n3D+ScX6Qy+MYvoq1fiwb9VTAW+fPW3AlJ/
uIASMZBfnnpCY0p0PybzJZHlBDv2tS7/uZNa2HQTyVs2+nKbn2Sh+YmjbGVlD39UCEFGx+ClJ1oq
CMD+lKijnCOxOitcoBPOVH/M4b1QFOpOwA8s1IC3CCbUt5JSieF7075cty/WPUA01j6oIut5nuFW
xzulqJ4aIleXbD3a6JsrIUWHL3X3GGWzSqF0dh8JNM/9gOQgPJvt3d3uWZnbKcIcEFZJEg8q0miM
Whb9jNFrbu9/BTohYxGVSjQkBqQ4IsNbECbY+n9DcL9zQBZTqUEFWabzcu18aVMoD011W9VPxZCc
eOJOgZ5CgnlwCp+tXCB4mnslM2KbMWCAfw1ryB76gfUG6LkhXb8vShtkpEi8I6BG0elJdR3+PqAo
iCwcFeGVqqTJXZZtykCY6BEZCmO8GdhbeEpP6MJuj/IpNBBZ3hImcSg4sYn+gtxE9IT0gQcUArbx
VJfM0fJ4eLldf2jCykTrxNrimemBGf14oGMrCGTlJ2irYzo13sKWWxDjg4gxkUTwjCy81gIdprh0
exj4rWWHXWm43azIkeg6TtdYP+dwXm8/XSNfkJCIrWo57SZfXm+pp3rQMgdIvGUwNdgQRj8agftB
DEEIq0Fkt9ghUs4h87obCp6eKGOfewccHSNWDNIQAgTt8UiMp1yNdTycFwy7z8d+L4rwy2iTw8ml
mL1GO7uN0qBLbPIMlNSqxiM3gOY/QnOqLjqdN+zcalE8ZeLke5TvwueUT6XByvfd19B7q9fiiehg
PaXFFvxFkOCjMW48JgT0JCr6SQ0Eg/N8miug2mOYhT83WDsLrLTaL6nStBWwvJoCf/bG+AJLiBW5
PFfwjhuRAmS9milM2Bzyq1QjWbsI2Jy6/IcRxQsKrRQ/XX5JdzO74oq4tXHd7mvTUb8Tc15kL3wQ
SoBLttCaOgStJ99/9IeSakGvQR+YjwLIk9jqn8fgiFrGKLCdTRRTuOY1+ISXHxiK8uOlNP5Ar7WA
gKCUTCaBJLQIyZsNmiETuNmd9whyVf/KtpHL0q2npKqU5HU7WenRSK1tyrQgvnUqYLxzWMr6LWLy
Lhgm8GVhtldoDQhid96vxTvhSMoqZuG/sYEJKyl3AiyxD1nqn0Xdy3jjiivLYnsFwptdTHLBT+Rw
fCj0HaSDpHDmVYYTbQGDnUN8pXLhOZhQKk2o4/auKI8cZkkwdtWfhg6GqGN5UPCAZ2TUAo14lKR1
M/owa9r2V99l0cFo44kUTSLQETh3OJQ2RhqxBd9dP3SnrGoVGQTkoPz56OwRYwLELtL4oENVziZ5
cv8wbT1dOw7YuF7Biuuqo/1z3RLnATNXtfSWMSgtw22VAMyjQgZfKNNVK2olyu1WNhaK/jM2Ax3i
e/gUwaw149JldL6mr88NCDRgx2JT7HchDDwaUoEXHVb1IjfaWFv7bM6eeEAqA6fnuakWEEoSg4Kv
HZJyNZf5T7O4Y7B+CLqKJPhbHc27nAD2i9JqGwQRqxSzyn6duq3mPrVIj7zWmf8+XxeX2Q2y5IiO
kggfCGi8E9YLGfUw6jMuGyIhVE3jRu5t7pYs5E3tu6/DUzabpYVbIfBdj7y1MZH+rXJCrLCJPyK8
HzHErVnFpRjldXOQaRbFfjEixcmqBD/e1EEBjUh1/AOkCjD8jJVaOCHSXM9+BniVSO5Ad63lNa0H
jouWwohPl6cM3i4VY565GoxrNaUL22qlvQms6o6OeLLC5ApGR7MLKym7ISF5XohvbG/OVW4mPmKQ
2VMcVwNhIXoTO8DrQDtha2sUtj/4sC1YQ1sVLR7NrMbPFruR4VDqgUzmNScGGoC1MeMdwV2irAIg
sqdupl6D9CXkILKvppxc80ZH0JW8/5hO8GaNq+v1dqEoUzX4ZDxujczfkdCGAUhk+LV0RMdGNKDV
zX+7M+YNqAyg74idv9mXry246hhig5lbNo4IvybLrApvtcyT9f/9BEmYnf1zwUwzoSlE14X8Wx/5
gY4jKQDygTS7CuaG4Q7WfraKPJzs6RtNiwf4YGqyWpIEfM6RKSWCwnyS1EqvQK5dbzz8618lYi3j
7olK3stL8lktD2WxEpjsfBNspJBGv5iqbWzVkphIuGzuiOrnTvjmu9zHiGiaduy6IBhYZeAMQbtY
kWdvDxVdRhi9mKFdOv4Glb5RUUNg2e4Cb9wfdIZnNsTfcf4Rkm7DHEol8BWT/60oz6aD3Rgk/lT1
qYIAofNjc6x9vvv2MyZlLM09tvVYEyTex/GQCytdcw1t7OqOTFD8smCfZp7n61hlRCyQjvksAWbd
ybKAVX1BH8fy5NniQBLmNmg/+kByrYf8CYnL/0z8D/0TS4fzDXX8hMCJ+fKc256AH697ZIpiI6Uz
okgZhLQUmCrKD3M7AkwJFcXQ8w5pXn2dVn/jYHn6Zqy+LDnzEEZsB9jxzswhWb46H6gqa/gjZ5r0
2fQvnsKsph34iaFAlk7DX+Xio4mbaNjIpQBMYTL70RXO74bZXhvSHNikZrAUwk9eC1IvuVXQ2Wv1
awDYXI9RUuxEHWdPp2vvcCZEcKQsWr6dICgwNKoESHiLmWOgY3ASdEqMxOx4yPpABamTCIPu9i1q
gY3V8YubYS1vF57mgx27K/gOcHszwuvAlBX5tMCqf8AOQ3bK31QGn4yUQNee1Q8e+quKi+y8ixmY
5sehD2I8Er219wKFSOnVSt+r3ZaN2LOH70YJ7UuRi+1JmnMFKMS0WVyFS5mfwZ5s4sLX7+q/6UxI
OovCNbgX5HaWDxwZjzJebwMlGw9VQHcYj/cIO1qqNevtt4hmSLynp6ktqHI2hLyo5ea1nuMtzIyS
kQK9uqrsUmbR/f2xQJtezAHqVpD9sbP9HXC5yZnmxUIJGforSRm4a6TgzhLh5REks6E7a+airi/m
qSCdS5MDy59lT/Cat6UML1u+k4VLQ1TePKHX1b7n+ZER8v36YWWT0aX0yh+w7lrAmur2HsCtW5VZ
wUtvJ2uD2Yqsvxs9t8MZ8PIE8opx4xPxN5OUQXZ3KHvcGchHzbHxIr9VtZxugT+XXCAgI7rR4gdQ
NXOSy5uk/cUDHjGCktrs5ErF2YpTVYEkWySc/XVuRorO8Qw7hYePrD7QpItSLZkFN/ZNP4ysyUKZ
Zmrnp56UO/vOlQBUzjlZGo0vl5Jtxec+UX1WYQyCXmwaK0+XWJoeagXlByLe0V57SyP3q3JEKJPJ
hsvV8wJKDg3IDGzYg7Wg17LgLRtZaGSpPVp3dmimzYkW1WDIR2G3J/PdcICtYzzq925itU3SD6Bg
LHfhCp7cNqiYwwAahXySXLS3iI5eyiN3UTdaIUgi0XFzV83f0Njc8UIEGwVM6yJ+VAic2Xq2s9Z5
jE9v56KsoXRYWNkAaJg28fsFEALEUQd9XVKIR9MeUOtyUq879vFkrNyP3/2onN7b8enIxGG8GCyx
VnaBRzPp0rOMJQigj4q/begUB1pc1G19jA0fhMi8VWTu058S3FZl+ZhscTTJZABTV06ckoM4CHaY
IP+kymPeS2sBSXShxqJBRTt2a+qCiSG4LkixH2+L598gNK2j0EpJcuivVASR/C0ALlHS3AlIyygZ
dWbLWCMsWIi4PbGc+wJBSMHMT2EodCOUNGp3gTc4JJDPycTrOYhYd3wGepFjYB1aL4mCO+zkrsfr
v1+gq7+rw1Wq0T1S8P8w4kIa/R2v4GGvTqL5kdUFOwZvdXLQaSzx6RY1EpOZEfCiB3JY2IOeuHii
eUvsxU3x0xjQ+LhN3ZZ2RgLwb/lf0ECKI2VZ6hOdyVXYb7vSt47ZJuwO/5SE1/OVkRkeZFcVRbUe
QQBf9ftrdlumrUF7XIH70fV8rCp4NzC0k195xsz1bmWf+YuaUhND6+KiABnbKAnpmXdqDOAbnhSa
HofWYeMSoVJUZY7YY2Bn5hPtTFtMwhcGND/RNDO7KlmOtgw4M4A6Pjl0Oqx1Lzfu11+Iz0mLmPFp
Mly0EfqvpR1U2D3bs+b+kV4rcw/oyI44XawdKyZdyR1iSSTGjDjM1barbY8Dw0DFPEPyPswJRHEh
KJzuHkHATKRI0laiVGHstymR0Ln9vDGxlv3UiLSy68B9o/h+E4c0Rcd4BDb5JMPhmhTbN8/xZSFX
0jV7a5KutsrM/jujApAQKnz/HNJK7aOMH/RL44eeBZsrGxcGEF4jw7vq1cCVKc853gqx2rn8fxgN
dRXa0TbjKsOuoFXrh0XqTNhcMmi/xs+WiHGVTDN9a21jmSd1krJcluU9jrIIfzONWVA2N+Pt5gA4
h++7yTeJgBH2HUHqONl4tFIYFbMAZb7DFYcbm1VdmNF5jX5qGgoM2jDfPJdbd/ZsGJ9RUfe/AwIZ
r9U2AKbO3WXT7vV47KXCHYWlvMGhyQlrsSNGaOelyNTvlhBp8NDbvW/QcKi9UUJiXUwpsK4+SA4L
GULNKqrEL+vLHZWls1hgSvwNO3aDmoQUDNwBkDKpl1jCzie1jw5MChNTiccQnmFs9Iy9qGG8qjmK
n/FGPF3bUxNPoQS7Ut6t78BqK8ooJYYeQ6uMnRVtMbT07u6PnKNi2ygJM3+secGzJbNQ7seF2YEN
vE8hqUghK9bxP6w5o6gQArD7Z2UIpNvbmnGCTmeinicYuaPGZmSLRsHJIZtlkoLyzqBvtju1bIwP
UzOUbe+AMbl2j6M1BnZRA33+Y+oz27u2aWznG/Y7R292u1cqqeKVdrr9hpn0Rw5X1MVSsN4/KuPm
1e2PubAbpjm14mMV1GxBJklEPKmyfZknnOAINzRjRuot41TMK8fsHvw2ICSCv3jG4U3CwLup3pQn
sFuaEhNp6ptA0vykbVTbdNSkVNBFs9cpPnnXjoUtFWrbkTd9OoZwWoCiWROFl4oIvt3U2dNw9plK
58Qs4I+jcHkm5jV2KMOHT56TJoi/KXvjbHLjoHKEr/5LyWt1B2SkXDPeRBlFsPycQrMUyfdJXQbg
4ZEyeJ7s+CWSirDcD2B2TLg0WItV/IUKZUTXXbH9Dv/pGTkODGYo9OZ0852VVynYsRcGPq6WpFR0
YwinpVTfWHvdn29hi8UeH7CPcS8Z3DzTXAuic+Jay3OETXyYE+FUQGe5fJr8RlvufAqu8vetSNpM
8wIvn+toL+dYIPNlBzq/vm7kcBoRthCagKw92l0YTbNBOhfD11I+VX/xr5Ni8/6xz1Or+s3mA7kZ
+MWU6pLhPGN4TBytPASgX3vlinBsR9LDi23oGQXuQd4U28Fo+KVWDdCDBcARr4unxgrIaTsIa/ES
FyxlddrjJG9Q6lekZsdwXvpuQUldIfBteyBexVd2qIs279ph8aE46NQw7OUHdlIQoXn2/CtZqBfR
RDfzeoADp5vWo5D28a7pHDH3XAwt4uM9FrsrIEaX1Tg7DX2InHCbZWDjbvSFu9UtBR2hiq3zjsNR
nwBXiMlfRv2J8mOiYp7mV321WWsPC8YLXNmsMcmi2uL0KmeWi+vqdQJquWdS6Es/JOeeubh2qx6L
kbTg66HokHLSokxtlM6DR4agB+MFYw7UAMpikquDO+uBCI8wpSu4alllwBiPBP+AC+Lyg+S9LMN1
j95AUt58oJh93nzS3fPnI4N5bRLprmqlO+DJ+PVfZcsRwnM2m750VH3j6BdspPUIFVbLJLEt07Ds
3RuclaDF6RzcbI/2b0CkVyljSR/Bzn3epqPlHrqjVk2XSvzhP09djtVT7xJqWbsV7LXJGw1y/ufq
fbRBOhsRy/hDhYQryRCCj1jv2M/ncTvfDaCTQjvfsyNKg3ZOTjyVQqW30FwdYF1MvYvPtRcdZ3x0
rVOhTf30qfRWtW4sl/j49lmzaDbgOL/mpMXPQ2mW5/B6F9u8dz/6KmsJq2zhK5RxBbxQ53sfu74W
CfaZHlOb8vj+U64uZL/jtxAY3MzttcrNgyqWdfB6YI6KP88yFTsx+T+MDnzU7w1XQ848GXuP3ruc
mBbgZqT7AeE/wGVKXbWFvrZqOl72daWKHunJA4C52925GalYi5ZQTrUqAKf/Nlq1s8QT/c3I+8fU
X5L3vnigjrRD3upNwb49E25nwp0QmljqVAAou71kg28OncnfNYJJDS6N64O68I8x7iJaIaZsZRX4
8BDPfQBf9kXV0o1rvsIhLcL4TwkXBscyiIjtESBYuP04BVNYOO3GgyfR5U0bB+Bgxf5Pddyycj8a
JPAYiVhMweifhbvopbLLvnQarcex48yHG8az9lMmvGzCM5vdGd+dQ6zf5mves6CI/NQFpo0DlNfm
O6EtGIUmZWKKbd0j/93Aa6PxOO5oXJmBaVnBdXP8hJHT5Ofq+ylwSPUFaFhsFFw4zfUAF43ME8nX
19wuNGqqM/jwdcaVRyxlTBxjLi4cuWgaCafYwzkfrYTfs/aa1m1MUWJi2UeXG29wPB0L0gaMzVKQ
mZCZgF2tqWNF8vK6RG/zIMWgRcD3JS4BA/5rngM0NztYNnpBstHuO0GVtRms00PSLWQZHEBnYkI7
tEmNyi2kzH7juEcsZgvm+DaYmKKR2MOsnKuGIrconFjxAqwcfUneej5blFKgxs4LOSb9mLKms8we
F1EBu4gnrQc5ARc6lxrDEqND0upqZ3ekjkP/l6xTQyRzvT/GGmuMThzVfa+NbqcSWu7X2Z8m6Spy
tTUMFWyEPCTFJ/gSlmmmPbmJaJqU/QumX0LZ4Qao/9EGuAXrMeSEuXAc4er5DL7hKIYgm5fNRaDT
y0e1TwZQKUGo/AKjL/pnqbrryNd8IKgosPZOqw9JVXZbGl6HIf7hkxuIOmZh8u+OVVG7KoWmF/ri
0ycRg9gvnGGwGEOZ67Jboa+onFP1xbH7Ow5ehhwoBQrzg1Z6OQx/qwrY4qqp4MlJfm/PC4exQuIq
+QmlCD6Cx+Az1WFpITX3OEF28pItL8vnsYzXFbKjcJRfyOGpNqEEEZRNW898JlnSn8wcvl1shJN8
BKWxO9aGXmdSru4k8J0SW8nQNhA655aymALOqd54i7Mlw0oWSaewCjfqCxjaL/Q5EzRSnlweXp1S
6Xfo4Yfnv/RXaKtiNzqEprSc2XukMG2hok1Y5OVblOjLIo0zVnRUBApVTAXvvOOUptY4c8214oeQ
IPKeZ8hamNZvV36UE7oMsNl6gjZx0dZdlMW4v14YnhCmFVGEvCf3eFvNQTyGMkBFq5ob0iTuzL10
w2BI6UvknBDta1NDSlkLnyUFI6LT0vcIgTRjw2sx7SCAlRNfseupDrSocKWR6zzGU7dS+d1+9XJE
OC6cUxbFQErZAtKKkq1mgnCE8TwYMsJYRDfilZAD3SUBpZMW1Zole42R9w8OYc78Chf79buSoib5
IaV0JCZBVt91S85GNGyDlc2ZTpeaRnpwJsLOJ2/Gr2RZzJpgXjJPiEVFDmIBmItBO0USeOqBVjPn
kr8hPleGhPYbM+QreNjNjIO9abT90QG1tMknnc3MANE8GPzH7MZiXW11vyrbb7Oni3ipJs164YDi
tj180rpjmIAuv26OL1a3dR126UofI6aIzxjvg+S8F/5pFlQEdqkGZLrNkefzo05PveeyDqpJ6RJ8
0JgfRcCgLGyzVHS6qScTd4depMnpG+kH3G3FqvUORiCoCWfkF8EGvXvJ0RCHHzh4AXU7jI9mHsF4
jPCii0KBsR4uA6eKcQdI3gIpC232EFjf/MVelehmmAL4CjJrPV0NMT9tD4+vh6HA5TKPQXqDzRJu
dgxMwjNIlT7eeUp7H6pfMy2mcCvEYUunp7yZk0AcCz8LLYd4rB1nzLlZSKZ0tmbfznIueMZdmbUr
65FNP2nRCvirp6OnkFZ+Pj8BKyOb9bb8w9aT5NmhWGNzncNZm0pgBGwf/iq9RAmTxNafEO/Xu+gd
SqyKaMfAbkbalR9VoMZvETcXa1+Bs6DvsBf/IoWXhx5alkI+5IOQJhNb9eom33CuByjLAvclF6ma
pRPIggEaIWczAiNwc/NjhJL/MHTXU/q6qlXvmdmJzGm0dAheZy1z/spLBV8aoj5cVnlrDE0l313V
l1KZtpK0chAXNRk6wR51eul3eO0ZvFlK7eG58g80FLeA/ovTNqTLidW4IxXSnNo/ZInzUuQSqWr7
TqDePIFKWbArsBumhEwIcbJ3ldRuhzBAIcNODVwxTWSNG/ubkv9t2drjG84x93kgVkorPRb8qt6v
uWo+AKZEVCNZ3BvAIh50g6juCcGOQCm7M6av55KssrSqlP/YFGWauEISyKPpl/18enkQVXGPoGep
msRUpj/qysQDJYtJebQ6PE+nN/gPTWBxCiX4WkO0bQfZX7ZtzWeNKwE694In0tSPcEKSb0KDYLLH
pKGg+u0P4h3qrlvMkyzPbOBFXzabBGC2HtQzzq0OnHsSyiMnoJcioqZNfMn2X4nvH2uP80x+onss
tCmfrTJY6CCE8yNjMWA77PZ3/JY+MoaL7O0Vv4IydrKjTCsd4YYHO0eIG9VKVvFqbu5QbTrG36kI
ju5gbA68/xMUhrGTruMIIYA9zhrodwC+YPKgdb+4HMVp6NiBbIknduxt3UAIZHfiJpROzliW1ymo
G3DapfansOfAIbczl9S5Y3tTNfSIGjJLt2Q9blAVqtitZk4HJ29+3ag/qGtgA+t1On03Quvo6OHT
k0usKMQWcJWk85NlRyYQg2RAtPS+3J0M8SOVh29wV0O0YC0U4B2gmIE/DjTGZ8bFRGAIas0a0AJK
uwbH4fH4thVsHy0dQhnNW4TlvoBrOWEOJ7fE/y7vVVpxObpGPUktuL4N4O1q5lbmKeO127xPcmvr
mRgNn7z5FnApYASNB8MZwmpQGH4Rf6wOmvEYpWChuQCiAYmJQCTvYwpTdURZdL0dbGFZt9XaybIw
OGLCdec09+dISN7yqYTdNaiyd6djMbLxBDGcV34PQYe92j7Xfh2Pw/Z5grdz20i4zJio62HoHwsM
grYKBLN9sTfhIQ0tBoNAmuPsozgmpJLc1s3XFEja0psEnWlzPxcszEaPw4xzpnbStRMC5iFIZt9b
vmQu2DaCsOt04uQghfIQj9moNWNvStu7NmANF3DU4Ec5x1NpvbtXcwrMM1M7rBbcpkTjToXtvLNl
lEjvl9D9MVN0RBSEHLTwxOT633YyXwrhTs1RvHJZEHKXgL/x7DQ9IykxoWv3GzzPisC1dHLmKxdp
DK5hxtmZizoAzTZFtTKrjoWkQkOWrC2SjoXCcn64uP2266gmq6+WZomTzgg4ZXn+VWunsvHMc+rS
+qrOui6iP641ESmACj0tyZctgfUmBKjq+qxkEtJwKu8zMKIbR4jeKYXOoiRML8Iu7E/0++y12stM
livdXn5MbtHDxSLgxk4KDVoqPiMEOTPiozw2+F7Pd+F+7GImUdDb6faucQdSXNQeI3ybsOHMhpKc
gErCWAldnfqmMrWg0PoRYnts6huqyzLGsp4cNNCtAyd4CjBhxY9oUCt2VOx9vFyed8HvNxRrh0gU
haLhbKflJ6Duv+YtfKmntJR9vPR3ViNWpyPJX1Y0kOBfMMROK/aXqYl3UrOHb+I/3RaPHEvezI/q
EYBi13utbTBRen0BFbRDdnDZjPYMETYTCVCfUVbmpQNWOV5b65O/4I/ABcx4tcmxHCIfxeTwOPH3
F5RGByNYIamEMLRyi5XOdQpk+7NZ17ATH1QqgFtvR5WSdvaQV+xweBAiyOQVl2rsU5iiKdVCMd4w
w7cRynB7nz6KdndhN7G1Lpkvlk1TJH4GmMoLB1WV/gFkWDwdp3sUYEShqgUN0vqQSJU6RFyJ1JDf
V9WNQZotfgAexoBqqhyZBW0VQHrEbKZ3f2mOt++oJKwF8Z4UMbMXpjrJLZcBYSY2XhdEN+EtadvP
CGLTu10SsG1ICf5cQyWF5bHQBrIiJP+O7CuwUhaAEt+JaawHxa4tRnF4Z/yqGTw3Ie/ZMar8rY9p
/yWgMhO60VW85WnLst/sQwIq3ltL73d5SnYwnxpklV2BLYCohT5O3aqKZVQjoBqmQmTFrGezW405
/Nt2ruC/xnhCRjw13Yu5NqKGg1WkPHg+ks87IpHbXGUMT5GOZH30DDqM4fmVRF9rMKh/5/rIjzH6
LYDLd9fZEgX6rY1+zwESILofcr5YN2Kt9z5zxGgl/t3vYcxH4srXhJTN/S74gnNxlAsKV7Giy2aY
85pQQBQUSUmWdaY55n/dgBSiB/NdO+aGEZV2zl4/X9veq9Nupz+q9QDe3hzNNVRh6356FCBofZMj
GbKVFRdrt7W3QbAntKT3EIQmPpTlohaCNMml05c0SOcz4ebbc2JfU2j28Zgx//DOpO45uqoNXkFj
hkMJ6Z6my4RRaeNjEB97qe09rshRdHMd7BP8wG7qZEbSM4GkPo/HXgqn/nNeN+lTNbMWsC6lpdqK
4I3Y+peScj+Psb6KAlJAzFWBFU4By3kPCFYwrZGKnShP475/Qxgy0LRv6H6j/S+0Zijrnq2/Azqh
yni9CKSJfiOzFBpXb/fB8Oeg/XeLVyvJZl1PxDc5to+kKtOrVq0SYz/Wy7qT4axjetRKgqRFkCV3
xDcVj6MYRn1lK3THs2qY2+W1suc7YGUYSnRZEMcb6rqVISX2q+qzNwMExm+Nm/u5LkRcS6UudYME
xGyne/TiLh9Q2qYIkCBs9rK6nqYyvsIRJ+KKvjG1ZJ1YvCDFJuWavyStTNIYImEVitaVdBx8cB4U
ZiD1DaCWxhwTZ5Euwy3ysI4YDsueQXQ+qUMygdKfN/Pl28omobnnl9nsRM2MiVLHKdhW7GwX3B0X
DyT+/plcTtIlfthjXfeNQWQcj8YRLnEYAyRQHFudbYbvZJbXMrR33/2rH7eqmmbQdkuiJJn8L/NZ
EZFVxrVBVZLmxUjAfyM3hdD4P0gexQIueOBj7rslOvKaIIk3TUzTxZGNRM5t4IdzCOCF3X84nuYp
YR1H03Jv6PyNDdXb6XipXiOVOMy39qkMAfA838L+G2t3K4u4FbK6NvDzFQW0uCLoPz4KOR8P4a+A
BnauvBv7AgIB9mGD+cXwabDwgExx1eV4gE2UqFb+u+HZdnYz6cW0631dYFwVyDXEiKxVBICM+mBT
AnL2jO3NhdYPSo539/J1TOmGhLNbBgSEckIX8f39S8HABCW5bsXTM2bTq59/w0g4fV0V7KF09QcV
C4JeaTNkKquaYb5Rn3MBSPtJ9kQdg+Ie5rXpB1RpuVxcx9m8JVJ8pcltvTXMe1qWfYjMYuQooA+2
7D1s9nPY8UjjlrsjF1CecbgTwdRq2AJC/AdNjTZzVt993IzfoEGp49C3KdGZh8rZf+dyQXweOMpM
We0MLNQ+thN+W1i20j1RPM05DWOEt3vhQtdyUrNxXWUg/W3J7vsLdV3O30NOj3kL+AwgSIdqZygv
xnI4SP1NL2Stg+fSsGbGNahu5Mj83BQbbRXMLZ0iKKV35S3xTAWrcP97UwGdSGg7OUSbkUUaF6kF
+BOWiy8PDpOVgpFSW6346rOAQY57ITz5s9l9e5Av/mVgCST2048iQkD9NcmrSH/xL3DCi6kTxRN/
pjWdyWY/8nJCLzyVMKgOrPF1ayMc0CB10x7iEoYkst4nUnEWWybLkNzai37fUuDQ1ewv/t9T3ejN
0QZITr0OSmoVeLp+fqnkOZZzTgWZwUqZ95gVoy2bNro8n/E7eETZpjRvbUYDmTj1XSlmfKEKuKHg
3FnNeoN/dAQVl9tYnkuxowBv0a3cQMG3wCeFOO5gpKb9JBm0Ejv3HG7t4vaL/cySNNNm7hTl1lXW
3OrRGb6kuJznD6XewhSc1BFrUvhdcy4sZWKbi4Y3cpRyNtNxI2IRZYZqrpNCE4cT4HCVHwRNrsxZ
IMTUYZN7aadOPo4nmNijm7Lhf5GVnryAj8LxOio6OtQx3kwOaGFyy1mbxdqnsDjhAnTGidxOPDLg
JHSZRSbsIC/cEwfWdL87VpmccVG+21xnZ8zGXwxRxotkNa5hmo8NruTTCUKHw1XBA+bLejquHtD0
YfAHX/Opt/izdBefGuHfytJMCSMVAwew77bsS/v3YZf/PknjXwZT/DaMUK0xjzqBKZMeua5KmD/7
luk9K1LpMrXWpWWMdRNXOF+BXu7Z+codsphMTcEMLik+7MpLKXojhOf4QZCILA7JosK4pKRejOCq
Qc35M4U9k20Tr41k7z6yForGsrNJ1nQLhdhyn44lraIIk0mvqd68hCvKqoxnQ5SstXOAnnFVbBpy
0f4ZgKC3gx1RAps/zuoI+NvAZZZdCkCrAgNJ2ri96l4REtIwak2D+rf5ic5GH5+CHt4XdxBMxVY/
VoYZmi+0BSisXaq90ppALAqFjCzDZ54huV40oFb+xwdESkF+GyGKUS7+DndKMC1rQW4YdhPGKN+5
ATJovG/I/v+U8VNVVN2JAgzTJFnhQn//1V2Ia3QCK7t4N7n79XHMWJw8K6gPewZ/XcXo6TmqVxiI
YAF33hoKYq+Hifn66TUvsujVFmk08xecDkuvsFrHoS2R4z0alCkNZkwLsshGTf0WhON9hw+logch
XTFatGSFtV9Q4R030hBxEKy0CdYTcFro2CM7x36Ai8G2Yyv1OyMu+Kbwp9hK9c6qM4pjQlw4MenC
pBGChIOkgbdTYLaO7N2I4r3C8VtaWj+cErLKpGlRocdn2+gtFfYUI9hN3RF0KreXJDmen3l69S3D
cuCdcihDPLL0psGk+jsSJT2OZIei9NNCri+JJxYwixE2i9HkHw9rFUVfwRky+gZKAhg/UZ1c6fU9
s5BhYbd80pFKYdcu6n1kk/D3dDk+46sNVew/3wxckXjJ9gJki/S2hFcJj+SjJpJFUApeErumZXui
S7Vf2fL7ME4HVKh+RoANsGTwcNBI8vw1lhHzqRQtRT8sgBqNxqMRvclv6bAeXtnifPR+6nWVcouR
eMELDJJTW1Is5NzGCwGx/ZbHLGa6Zl90zpzebrYGuQ80wIBfgipso465JW2lENoJuh2f9Ha9JJkm
Wf+3OGmY0NdXqkuwZNsByAKLjj2azT1L02koqR953iYpluI0crWbNtvEvJhcOOGsSb/SO0GdKtpQ
oJ+GxDuOPEfLT4Fd02nkQGERF5sqcN/qTUS5NVs0rKzrwlC6g0K27znKFZQ4nznssstYraq/1/cA
otcwrGNmKmV/gSFZcs/JD01psngfhu64hz/O0/PrH4Oplahioh2hSNzNVsafFwTzy7+erY9PoYcf
CZJFDjCS0E8u7rtWyX41BDPu1KEfpfwwXte8d26RTAURJco6H+/qX8lOLgGghLfW0KssXu46Dstx
ZhyCOZtxEMIXVZVcIkb8VWrVch2bNmxm5kpOKrl1GjNqGVIZeOLtLLdU0eoTMQefuiY44HyYk36e
AgyDxRuyvAnglHOZza3WsEkXWFHBzQ4A4zU3hcucZuw7kRkE1WAkcU6Z4TDl5lTE9wpDDPWJmO28
HjNXvoA4zNP3P70/KVCdZgXaRqkT1W6EuOhZpBecm4pStA2IffC/kLk02kePoK6mNB4BEy0w5K1w
RtFYa5GhixjBbki4XTmzI+2ja6A8U9NGIvaYGwoF0HgC/ofqJhKMudG6tttFuYIIV4p86V+5xsGP
NHJMztjlHYmVHfoZChB6ndj7qgthdp2kZCYCMAxUXjBTkM97rP7w/cbyrIPgc2It/unet3xUkPf+
zW3Bu7AKGfV4VhEVzHwTBttZ2RBnADiZtBR0NphVeUpUViwrWl7Tj1bXBvuzoX4nLpI1i4NAqXbZ
DLJCqo4bLj7DzhKOf0MsolYm4NKe4ea/iJDJC1JkOQa9P4nLC02WJy29w/cc7NL1Tbrj3BTKbAwE
NeDAnxDU/XJw3NXuaN1L7xTQE69bEISqxfgIF7EBsaTLJAVPL+ojE2XcYDtk1wYS6kdcDIDzfIDT
ItK8LV13Zeihf8imT+YqEMxwk3aYdL3+K98YtFmjsWdpPP2bOc6nHeYd46+OaRSjbFUfz81R0xUD
atyPXOAteoB500scs3Z+pHZmAFqeieXRrM3dQXFV8GEZX4oF1GcYWJY7BszdTjRWau3NcV9Gn+lR
4Zjy+TJNtZyQNkAUBxvsENYc4vOEM3zw1smS3WnzIpQ+sREe5kQCwY+aOVS436whQ45HvcLGecvY
H+fFRUs1Qfavqg2rhsZmCOyZvQhdUJPrStgIxiROOczXOTvK1v/Ly/u715rJrcZR4hYtrlq5wDj8
xoBgPxewv12Y6Nft7mqh1Uv0UjfK1iP0b+q+TmtcSmmPk3AZR5lxheBZmEJ9fDh0/BO/598MREFN
iXvZS+DGWN2PMEZomMu1+CS0dtUknoRhqJsQEQObxepM6qSirfOeKphHbN/svRhV8syDdnO6bWW4
BwVoFfJqHL0J2OHTdumhR3LFmCE45xeY6UgjLQl8a2hMzuyScHeCN30zoT1hwRCQ/WWn668dab58
VhXtSas2KCqnm8BbwBC71H502ROaCjlaSFSTsd8r02zJFa/3R9xRbklA+qywBLqNG670fnzNQJw4
9ZxnjpgXzjniaA7u8bjrgYsJgvoFj+1pANy32VJBiTs16J1begvQoBIspZ01u1HRvBRkbBrllqfP
JHfxwYVIfisqBv06/7JgRbq2G0US3HdFWGnrLV++I/dTWFhZbNVTnIGLQEoQlN3sK58BoLqMKv2F
ECKJGXYEXoATmde0p1xVfcj1IwXErzVsTeDyn848CoH6S3qHSNgBgIzNmQ9J67ySdnfXwH0suZXL
P49Rh2Vc2GxNree6zKS/zCWDXdz1UyPkM6dCYL8soCe/6oJbz9s9SIs8v3HwsFK6znvztwvPY6Qo
gpwQTs3pfrBUUuw2zbAGChpMgHdQif1dxIKFtfxH2hhsHyN/pgsEqocpdbJ5+NnaqFi6Vtoanjio
ZmEiJk0FvO7M6X0D6p05CWkIVFXr3CSKxKCuzmTn91EdHknzAwy0D9SmUUXThW1PKGipUgHEv7E+
sjUdpElLcczVSi9GqjA3V+1/86Vpjx1XpRD5ZYWeFJ15dEW7C02v0pLFK1p62rWE3yuezjBiQQ1v
k2ZfhxNsg+CMZIkl3QWuCixYLz5WdZ6y90dRa08TAOGXFANVEjxmVA+u/CQk5pm+vUi37Ef3e9TX
ybdvDI+H6xEM8BLYszeKHbwdRx66iYeUMI1HRB6ZWFMQC+WhQn4vUoj0RWyVmS1bIEni8IprGKPk
ZXl1DyMKvgaJi9jterwQcpdb/3vcOt/bKFy0GVD4xgagTnQnjZnpW2hQR0jUMNj65qD3IBpR9Xgw
JCofaVqOt+ptnyE4Sdnjaun+xBNBOaMLz/v18fSRFT4YELndee8oD6wkvmZ8MKKYL9qqYP5UodIf
APjGH6CfkYx/E27JX01QOU83xfe9yk1OmW30gSq30jdFd0+67ppxz6lzwqLF1mxj8tt39JVOP6RR
4KHFn1VZ4QwZNzzpXWKpKSuRwSM49WVDvbIMC0jvXYLHklKz0hnaI3mMtXSHI7LPazepB+pfgWge
VnaRVvzqqPSZbAkSMBrCMXNJOQnSnuvO4nRK38tu7x9zgXBVZiZo2dRGBdKzktTj8K5HR1YyZE2X
JTzIEedR3g7CGDwy4xPQiKsMz6WInDrrFcotP8/+1gGSTUNrSdZc7HNm5fcDNiW40b2B4xMSvTj2
k47BB4FNAp0RZjRD0RlVJLNv0O9LMiul3Yv8MZb9EfDKk+LqgSmb6ra7eSzvM6brnNkvpiltQ0qL
ygX2CEM4nfjaYClBjkEezSjJhGbxduFGnwDxgcBd2s9dZ0zCUPt9dJvOCztNucADO1AfURMzGa2J
7AX7OYwvEzaVV2z5bvUJNsPnEHYlO4Kh2Ozwgqb2wNrloeVShwIdKkZc3WpFUGe925+qIoB32wWW
jTsy9hmK/Xns08MsecRl3FAHP891sXYc+imktNQTwT5kuL6pFD9/ywVS4tl0Ga+uHoWi1UwnwG2q
9k9ovYrROidn2UdU2tCWwg+WVIRWbbTBtAjXCttx/hyh6KZxOdU5Wi3Hmzv0JFmXARLYZqyH+7mz
MGP63VVOriV95HyyrG+aL/YmEqyR1QuFHS2lxnTwX+mPEkDU/1ZltmTPZfSUQiQXFJ8ZS0MXhPM9
fQw9jZqyYMlkUjllRM8qryYn0fwNtyWzR4pZEZaZ3Q3ceSlxuzsLzC1wBuj1zS003TfCNqW930Pm
amL13/QYCC1KLLDfrxCl/ZZH8HJYLK5zMum0e1AP61KCp7qRRBvU4ZS158frXbyK6JDDKSFi9Fsr
OklzK1As/8tKAPHVhrBitvJnwsGSQeTDeElXIVF10+8qZM8gH80w9erPi9k/JrCG52cf3WiXQbNT
BteIaYdaorqinUdFFOWs31S5uxh7DiSOD/6c09qJkwfCpjBgsPxVrqmxY2S1o4TdHj7+78yM/LQK
vqX9w5mrjGtw/w1OCTLhUYqv9hn5h8yM5qk7moy8GXcLPCQilznCNlGqUbSZAKDl7SSF+ElcqW2/
mWjQeWI0dk9ll/8872uqoY+Lr76ODMdG3Md6XOC2oKt0uiSnFP3Rn0ahRYWM3Yz4Epwu1IBOLBd8
WH+Vibe61THJjaW7srJmLdMjV+zlNkg3IiaCFlUtofOTK2AJCqSDazGKsevFOgrpR+tNssXzyunL
cm3ZxjfqpDA9dXPCrbFkvBEzAyOos7qgMS3PDA5UPbQ0sAdahybsMevHjujd4uF04PJHDd1aRHs0
Yv5QTfcXLDRYz6W+Dwq93Iq+2iLZ0QFJD+8Jb+Vm+Bn9OiYm/8c+zf0UVJFohQgFk/u3NHMoewEb
dqmerQf8up1beAibsJsBghW5SO5Ryo0GE9MJOFSFZv0xXT+l9xBM2NP14QUpo8x9sw/yemr50Nwl
0cye0Yh3G9CnAMHWCMiK5NPuFecnefgwjlpuSxTUHnP/kksIAkMe1L22w63ZcDjc7/Avmsg/W7iv
AwCuzUqGzyFg/U2O4oxqB0xWEf1trxQdLB18QBPRqEVx+9lCqBBpCH9IyyL53UC67woWXHKengUt
yhtcWu29AUazs8n+//1s6VzOtRgvVowGVVJ2DCNpIHTPop2ue93+IByiaUPI0A3usKVPQBNtIhgo
Adq7PTcCNYKS2hII9bP7Akbk7gx8LXv2UNSu/f25kwMNM0X2+FP+lwY9Wuj6Gc+fbk0qJGQ3JWQh
AQOUyd9v5d6CVeVbYAQUW/C0ULws4oBpBboLFiiaVYly7YR7A+GmujK7yzU82eCgSoUcu55bc/VV
ffnjxP+UscpsV5JEYQm1DQXN2oy8u1uD4+neDRGyXx5cS2G580DkCxc4eqASVJ6XeZzyb6CaYOx2
Pm0pLyYiWqxOCVxo0DbyhCny5h+ShPQjuBW1DilNsc+xqILrqAwPCLDziZpincZgmB0oNHp8tf2q
C/Uf3D1Dwxky4H0sA1UWXJ3nbhHv1tkX8y0NSbrvA6Ct05Kz46181WTp5nv4cTbAe6B7+0ZYtDF0
0cff9ZOBsKndA5xUowS0Z1xHSpsXwXyI+PCG/tvMnrnKQ+lQ58CH6r0YXAQop4tfYKn7sUI6g6xf
GisjW5qCs6R99AEF2+6IxBQq+O/DcFjLEOsYewQoVAM1RRFCHMolJGGL4jKyA5JEZ1apWQ/coUUh
8RMoa5LnCZcyXkIiIjlfq1pnNrSLvu9uucvux6nM3oTIf7y1lR2FTe4XnMdJVUkBxKMvL7Zp7lRa
sHvGleZ3zFQhiVlUdhm9eaO+N2KAo+Q16YnxnxQ9wJi7DcQIG8u3WRLHLP6K0RmyeLK+mKiAntoV
ctE5gXxwfg8+X46U+O/sFBGxpbthSB+hSfJ21tWN9BY+7HphIpw3nzbYjY4d5sa0N0mdD3Xtkcq2
hGMYMAI1Yso5IJnXZGZ5nkGaB10jAEd30wSLGVd7aC/UkN07PcFUbwaMKoOkvygJDzDtOXoMeBY7
ArAVgtVXaXL89VQj3RZ2xKpVZSQvQ4fvUI9qLY7NZM/NvAt3Y2KzYflhpRGJ6932fMWxt8rVfmG3
8IjABezbfnco5azkQuQV6vkew7hpx+02NON75Jxu24FEaQuuSv2x2emguGb5zD6GalBg6ikMZdDE
pYQEvWRGEorsxrUiukrZiDhld7nzj1Gv5FX0zylUs38k232pHxuTCPrv1NSZlovtF2+ht2v2IdE7
d4z/Vo0DDR15U96DKzMImctMmCltymgsXwJ9xSecVqSNfwvpFlsO+N6C5ex0J7tUsBphumT4TPkF
rRSX8zsVcGM3wlQe7d1LrokXUB+ilVeEWovrSdux+jPs7+gYd8iEphrdpso3p4gTfUfzMlmCJmw6
Z2vDe1a395k6NOMmgIkYDGkau0QoFJHfVr2xwZKnMsAib9M75wteJIk802lvJzmHLC6d8pJom6o9
4cRP4cTjs0dIHg3666Mz7QV1SBhHieQfbZeEHOQrUzOGhfhisaWTkkxUpGP7+8gmrvTJI5Seg7wh
O8HccbQzSkOHVsGk0Wq59YO9suKZJT+8jzpLAmmreMnmpjNiGB0oNJ6jWSAsTwkyKcpukBpUtfQA
ksBSj9EtuGrvE06WLK9eSn7utEm70ffEBQz5LH45p23cGlTW/b56T1JKm/C/fzp8TeiiWsBXVW1L
0s/I3TkBHHC1JCrVjcaTDJs8QLY82GYIAA1P5W/pzAfRKamH4whcP04tbw5OdpHdF+JjTpGWBPzq
vCsjonhhwtjpmtrCQozv9mtIgizf9numZ7SjbiERPGduHRPAQmgvaRVSCqvpvMfbkU9GxRLvk3+C
OF0SJ+vdRBoCKcfGbC32cxN6ut7zsHtNngC+Vn+4aeQWq4y8oD94LOSkA/t4km8VVRduHQtpXEyR
eDlYprhL4DpqqLzaPj9YQVMoHGsBQ9iU/tcqfm1vGB8xhbMjtjkLCZkgYtcs+x3CGJpCxdjIU9ch
a/Qr+k4GA9tp4kfZL6nL6kwPpXH7t5mPFOZxnp9oMWB5EbAzsDNbEMcGm2ID3gcff75nx27QX+2k
cdAnUv0MY2b17g4c5qdipDxJu9G+Vcb9arAtaMJYRfSV2jAElBolsFI86++rJq+jOP3lLcERdPGV
xIOi7eqBG06uab7NlgOwM3ZnRK9+lHaoSZyhS8zUE2PO4yXp2rvk0rIjD+wksh+e4/DpFMmYDzeY
0ZSWfrO5hXNaCUB5pJTHUscjGtvB2sJSQW0bqgXTgqvxhZ1rAa3xyYYNtJyp87pcLBi67Bq7wg7c
bDxzz6INdszsjbiHZbBwbOGHnLbEnRbN75iwuVDBQbCXXzif2v6ZNi0PghMFDswNavfxW966Jr7i
CadvYrdLLfgn3jFxyd1q1eCuZjP6m4syspJ3rU5VovJESPOU6vxcm2ub9Oo6y9zhjk9+D8+JoUNJ
SHJ/AjmUBvWD7/cb+RNZGqqRfZ+rr/k7TFl5icOvPx6N+F7j3Z8SczQ8IoWIhsf1afS1Y3iKa0Fg
U7hl81ri01oEuzzgwbjiRfuDXOI46dVXEHOH/Vw4kBsb3tQulao6WZ546mq/HWLZgtO8JkNvIt+P
il9UX0NWdU0JIr9i9iqSRA63vNGxohrVIuD3U1MQ7h4LTyu3cejBdHixoVbDCFau5lYPy226+N33
1n53ztA/DRr1Xop5fLTuCfud64OyRHwbXILBOHCBaKo6+5pT2/piSXgRPXBIyndAwq/42b3rfF7w
J4wqYsRJ05S1BsxcuZY5FYuWu6D66ra+iY+elKkjL6w3AFtYl3alCW2+gO2ug/3wNXeYbvReu8dF
GJBuuD5HkKvN2PFykG8sLdfXqhIKedHjpB/r6q65AZDPw+UlEKGK8hIWRJ0dd9+QSUfL3IN0i3zL
UlyJu9AOZ7/tGXQWpI0CZUJL4XJvTAFKD/kt3bzFaIq4iXHTQfBLQduDU4bdAlKjz9oY57t90nVo
add0m+wF+Vq8HZMkClUoIJGcvMVZPn+zDNCUtukYjH18OzRGkE6S5MwT+O5mimVh2brLIDmuTb08
D03pTuVZftTsTgjyDK+r2N1BPzMkKX0BkHuScvq70X4ZkNROCBn97ADtqIPY86tUm6+MYuDvWRIT
9BxQv5e9gLVCUahencbY1o8EndGUBP4QU/V9Onxxp3pQ1zzmkfWO/iLzSoNR2WMsgYqq3iOPHDIu
Pxau8QBaqnyFiecb59k9I7qaQeZ+hnEIM+9+CParfHokbyshtpg2Om25b9BgqQaaNrmIrCMQFQfP
b6offl37WWwuZ6IlivdkZgV0uyiRobWZy4/RbRENETbJ6LvVoc8VwQm27F4JgPK6xVbgM/P8loPk
iuDGmyrA/ogiS6I5MmmbEl2chvPMvW0RIBRy6CFdqCUOCyVA3B8bU3sHglY/e6CX3O/JWDJdNHGZ
YfD4QLSFYWZSvDJRdeO4FiSvlDKv1NFI/PWyThSiMyWmBNppgB8SCjVUgU9ZYGwhDh7pukSAm8ie
/RCyK83P/f8VjxvC8aH/ypUDV4lxu3/v7jk33/rAhA5neb4k1E0RwwAYveMv8FjSQWl3dLYyxhvL
FzbQhbok3n/mq45HqNmtTDIDER3vqdc2EAZbeujtnMKy8RJ4CU0BQZ/dyxPI3OTdqhck2ont3rYg
7+0TwwUfjwg8fMoB9G/Y8He9CKynkwsOYR5tev1I6kN9JeDWAMJ9HoLffGLC/kaV9uwCjm5SO3pR
q61h/B21rIuZNJXNYYBiyNk8oOh81fogwSilUL3Qo9NabN5XzEy3dWn790F0AF/k4viO1g00i2f8
MCMGB0Di3DL3mpnvAyHWJh34CZqbaLZPEXAcLl80f/0097ViBYb35Pz3YlAWGqd5BpVLQNvlGQMy
mNL4lW8BpYi4zd/zkej9VcBHxRigXh4YXoGUP+R4Z3FYaT/LJP7bBh37rdlTpHInO8YP9rfVDrA5
ibtO8P2fN+GcVwCrX7lAGb6jnv8U9qEEbhxPpBvTw+N4J70pH7x/LZKy7UUO4jPxrpCS9TmyPkTW
01cwSBiEd37OhSfEkH4Kums7hMXVm9dMUhxTHF11DJk8fLa+rKkjDPnSKf2yAaPk9wjB0nQqZxVt
ILIK+gvb/gNN8r2MzzpnkBKz7AQ/Md/9YGMZ90SqmjHOQ0/6Vy1eP9SZYsSgETcQLTF7wHAga7Yz
Y8xdF3FaFq/2zKd5OsvbXccniGnvI1h8MHaECC884WUbFGl1D53mi+4/QobU53Go1olPCkfe5N0o
tJqs6UsVWOBqeHsq36hRGqfdjeEfAgnWUtGP6rQAYhPphuGoCTjr/GALFwXYoSuQTFPHKJrBHaUA
IEmaHG03FsqaOYQxblQJ1aTHB+CmHlvpmQ3oQbCklh1YV+OF3ZfE8bCVtgWNVL8HpB4sYxN+ahvE
MXrYW8gwyNSVSVlpXTYd7F4yV9gbIA9oUtf66jhMghJloCzKKLg4cbnBTMr3D/t0dkU+iUuuE8tq
BHabbOJPFjUXO3K8ZPdb0EWAG+fLc5KVE2xII8UkwHB4eXIC1bkLjTHgtmH+vFF2FnFIzq30Jdu4
HvmsEnDA6ibHziqvAE9jkd7pzKpqIMOZQN6Zvs85GLASwaW5AF79eEkBxH00dyZcssLHvfrq+M+X
4HArAiHPG0rnlBCHq2VQKQLCd0VM1sSanQJYq4GUl+MrlC7xanRvpp5QyXk9PR5pv6TI91PPWO5D
NBds+02r2Nobo0DeN5ddrUAZEolCLSwh3ZFbF2p4BFrftojXGJ9FtBggUKizCnfEZjrqgzySBADU
WEGjBoeMSo6p2SLnAopf8mgL8Ffzjzmpv5UZhgJycNAfsG4AARP4rcObhk3JhLTkhi+6Hbp2WtI1
f6PAUe2IlROte0nLA3taPD47yrVNmlD0X03qid0cBy0h80f2Vl/Esd8riGndqE3yHJLJmGJAGRuD
kjKnY8VuflydNoDdg/2TxXOcWzI4idFA3xZSeS0scqDBsXE+gj+VsCV07rzGXWO3nE8tddrhx7/X
KsMNXdwWCVknGafwVmzWdwaHK2x+aaqmYq6txMst+zfeAUm6uqy+skWiSzjm+Fny1AiXXOxiuXWJ
RKGnXgy7ZpENQkvz2fKNyx/9XPrQOY+dnShdEcboqMSgjlXiJSSbQiB8Mb8AAosmf7Xy98p9uY1Q
il3YyvyskB6tq1au0BTXP/oZSUR3VuSBbBYJXGj146hS7ybM1JNGIeSQZWM/QezjyrXXfNtnC3Q8
77yfUouPnPNnzDgduqcWoeX0ctiJLpBe6n43z70CTrSAWKShi1heIsQCjnuPKIzCW/oTltzVFdS9
/OBv9ervPHJDjfMfPWjZ6uWVsQmy90Pk43HFLHlJqwMYVr0X6/gLDp1YOrYQYait6Uc/7MCdoYYF
JrF9/RJbiUC1tTvGHqvouZYUkAWt+qmfbR50ivrMvy2j/pwId+d4GnLZFD4Aq+/5fz4QdqeSCadW
kpTepje8I0fjYiKOA0UVEdn7lkGxsMNZnEltLmTGIc5pRo8YsJ9OnMO4bXWIBXII1FJN4teS3I5r
sbiX/ZUQZ0JCAnTZR43gMxsJyi2wqaoIrlk8X3eIrB3cT9LyborcuQ8AS9GKfk2/9ceCEZGia0IJ
Q4dNmXBgAV4VPaiaT3xCwsxtpTCmHrD91dBfXo2mQCfpazmpGvxbtWGhJhkLecFpkazQ0o87ESLC
91LK2wT/2xhvbPKW2CPgdzOwSd5hsVzDStgfePWlWKEZKXi9URtvO4zbst7eEz+gse6q46jHzjCp
ry3oBRlVAtHp1N04MNzGP+KUz0+nVZ51bFK7bniFNk6NPG4PmMxIzNenq/7wfK9WKDcpPhhX0BQP
LruR03YQbxDZ2nbfGIkyypOJ3R4RZ5kzc68O3j+5Kp1uXUHPdNEYb2pM+Qg5QZl5HUDOqkvv4AiS
azCj+vzgdoCC8hx8YlrVHezunZZvDNL0UOdjK1q/DlWGHf3DKnYUc2ine/EsZQ6c6DmyTdLt7rbf
AawhQFeq/dYC+uL952JwaXLqJwFG0z6Yd+RrRvDrT/P8WC5yZ4nTQafB3FdQVWij6WCQB7JwIm1G
g5SQj3rVZFbVaGiJdszi6V1S5pGDROkB/6HIu18acnnKBAjdYDXF2ZaGR8Kc74rUoRNfE6jsaaqH
GUGOd412Iro/scnHeZLnS7F2TKfg0z+PJBVNOF9/sr9iOKwg+2oOOhO/ABGy/CAFGNKkpnPfUUPJ
lLuP4XbOPbXFmu8qMIJ3EwGj4k5MMeQ2W7DizNxu+NJLGS3Wk2IntOgrlFbYn/rf/YQL/L/DlItI
3BHHznaWZKrlW1tOQ9JyA4jT8BuvuNsKcH0yeI4Il0KgJOX2iTg1UmmSA1LVd+ew79Zi4Inam4cT
9c0I36b7FHabdCu2VpnvKCgCGfhqPiK7BcQz+gHOq+1h019Ew1RCNmAlg6uUdlo0nsecFVQfKTrc
gH5/RS9ncgxZpEzrmq9JaB6V4Yn/z+YPBxSePQRSKOqBHC9rU8NMyiCa8l+j+nb5NStiYP1/YRh1
zI3iZr9OSxbiwNpM2p+9IWYZU8tNfEFjc45QpSwlucq6KXldd9pKwqPZMFWz16WrYFgsh+TTiWf0
Ekg0rdcbp1ULujljHQIuC1uFmniRePdv0EIdaEih3OcpcoMRGPfNdpMsVoXu1HGoTNjo1EyzDF62
/UwZxdxYHI6+vRIvhTB6Mkg3RKJpk4xTWNfnbNREvTZjPwRePpVD7y15Yigu2GgWFj3//Itx63xb
K8dlHSiFdl3tCGiLbGbrYLMArKsmprigtZGJNTljmkgPOYxHU/IFBVKpESQrgGa6/560Z7BUSLLD
wLyN8qgY9Rgw2PIzdAshf0bLY2FNr9/RXP6cTPg6hej6xjpLnbu/kYbWFmmfnFm1lt6DKupfb4mc
q8JMC0T1YVFyWNcnQtT2qQqmQr9SFrxuRlUyHeY4UTz9cC8NURHV8XycCd1Y4yRLJgsnAmea7O+7
ag/kaJfgdZeVipvLmVt3lFTsIxRfAG/wNl659ll9Mo39ZJjdeEcagmeXnleGlVekSRpxG+Ta6mja
oajhexXOpALn/ZR0457nm9hI+eMy7R1znh6haEOE/wLj8jFZmmCvwgXyLh49XI2I3Di/EhbVwKo1
vE/xUxD6u5gg5VZqkMzwLpCa0OnEsmKOulOa57VFLkFfr1L7hJAgnwxeDGp5yQA+dC5NBbCDh9ir
ddYUSDGHVUGX6kwIvHv0kkeG4GsX+Y6XsP6qtv063v97qYAMfDt8cu+R8scbHpk2NzSwRDqlP/nm
hXH2hwc9P6f5ZTBuyr9sAedlXDKdIcikM5qD3CK7vonv2EKmFI8lkkdMgL5ZnX9LpTtJvx30xiCR
FZzbMbxVTxhuZge+9wMN8BtsryV7Tb6YysEp4OVIvcpxn3r87Ge9KPGVEezEVkfxeV/bdh/LqziQ
Fmq4SRByLeZOEMEfy/ZehIHgOIa4QcXEDr6eUMlcff1XrN5ilhuwKsTlF4uGGO+/AEKtxFhjGg5f
upbJEuoyBKMOEZGd+biAGxI6yGhgJiHY1YlFqaIujCovKpVHHO/qAyY5jG06KuVgT6ShQN3FXiSY
z6GkAcO97Lg3Ql17rPCrX/PqzT4BeJL1PEr7gNooT0V31LfAYiOxCgobf0IuGGDQBhLjDXD9VfOJ
LDNJEEm7nmmygijMIDZT3dYTakUV7w0/3/z0Od2GOzb0U6ktwXDrEeg26Cu+uRQFXLNAoTk1KQJ8
3oBVL3B8gF3NT8jB1waGwg3A7istkxu5iwvbi8Q79VYfLfnhjze242T44ywFb30ZpTTFimpKraew
Bqiqahidb0ejaVsbJsDtHmM7q+R6w26aHPooHZRob6CYNwGE03uWBb5GKtPiiZHEnnmrKVpoyd+4
MXc0xSXP5ytffZZPGfxHyBAyWUO1vmMcaOCAVRR0yCceLIwAqrLi5FbJ254bcro0fa4eaorevjod
71AV/vDnCwjMbcSCLFjHydZy2PY7mUKoUoNtblfzBLYUxW1FuH1GMvshdN6uOPmmBMoW7k6D8n1m
yhHV3fLrwhwRE0jpXWgn5OvD4ELXCBFsAccCLlYO1gdhRiwWyKN9Z/uvv0RSoIut/HHriDWMSLlR
pPbreKDzx14Ji+6sTKCyYz54dt20J38USCqoNBijkNC0KQ+GhKTTbCIJzryBUF+Cyci/HmiFybEP
DcWukunri0MJ9N8TKCyrWFOcm5zwxk0cq1Yr05Klsixjczpp4PveftM5uSfUtrCo+wLcdpZ/ckzW
OFTbdMR/xXVio6ofmVab2Ddx3S9shF2kuhjBY2SzfswGu/fpn4+6JEw6wvpiM8Psa7x1+O+FaZlD
SCn1KbgBNH4W2+qbSQ3gdkMjbNbEJ2dUxXoGjmGyAQ89H/23xNsMI3nz6L/PjJ/rhCeSL5+AtdXb
VHGhKpGV6agvca8NPTWAtO92CqHIpOM1F1Yw4hr3T6sKZEKLBqO72HLBsFxNtmHa5gU1BqF7+XdE
HZHPhcq0coPaaTkTZDhCVuYXIRDwT3iBu8Nip05v78jc3ONIqeuChdnJbPeqwhrkbZPz/prsl811
A1m1jRP6y+WamY9jvFgRkKJkcHr2ufaWxULpMNxB0K05YIIlON1/V4xyHJU5Rpf6oISfgsQqsJWu
/LDkUk93eEjkb23ESsUTmgFU06C2tmOLEK2r6nC7bpuM0mGBBBeUl/koR0pLJGQD1sgYO67t6ErF
nNd2MsY5z9m759tZ6jFxsD8jyeEqGVsq5IUh7IkRJFnH90MR6tZWxlulrS+rqFDiwf8w3/vqFg8B
JkWensXdjF2T0o5mFkur6crVaBmsIfgDW3ApoVNSXmJ0DfuPFWiM4dXsVVQ/7Xx3TRxGVvblyIFw
D4avXqrcJZC/oqJGAcFcZq3Qbka/SA6/Hus5Sk75vz1HpAGMseOOILf/0BCHqBsZ+Ar5AcfK5zY+
ThwYbzh/TN/lrubKFZ0DlISmGgS7Q+BbYGk1mqaB/7MIwE6M2WYwBeqAz1XY0oIT+9fSto+JEGvt
Dxu1mN7NNo+HVCsSOOy+tNw+I+/3uct4MNWBj8onvH5FNgcZew5Nynaj4Qt/+ea6IjRv5ObGqrY3
IXF4E7Zvy3lveuASwlQiBAeVdyA2JQWCNRPNr2I4OmV7b+7sL2F5YcGfeEuyrch5i4qx9eniZ8el
zHDWMgGtWvctPg1E2gxtqgengCUtGOl89QE2wF6FM2aznNO5a7gHDfLkwNPMzOs16pRbdQtTSBl3
fQR/M0BcuAFfikNbsdoOoDzLF/8ojkSzSfH9FT0jaUM38EeAgzhtY9iJz5guATLfQCm1hCyHIdFL
wWvsxSxrnXL2eoLq+haYAVUzBaPo4m1jXG+Xw0CgWzk1BKqzL9tOQROEwa2o8hr6VbvfpUWNnygD
jgyz//BeInjCb9+N4Udgm0bLe6lvLUQ3k+SeSzCbfjcyEeF7Q/PmoZYYLC2GI5NKEFblh6XqPkSU
p16pBc/EfTdW/QhrDj2es6GIUfDN+RfQXt2g8WqUNGMxm7dcUcqv4IPxY0/uLFAVHONJ7sV9mWWO
S4+Kqf3CBUWXpIB6MXwWgnmiitx9eg98HMEB2P9eK59iUQjCb00T5fHwkFgq1Ph6kaGsmqMHLzuZ
K1JsOftENwA1bUGbPI0AAQH2Z2vnLq4UTJkw12nOOG+xKopP+cTk2kXDOCisALsVCZHSDvDiAbUh
8FRsilQBkSObwSNh0eKNgvXVuCjvdqeztTVxboX3py00AU9+k3EpatvSNv/EcNQA/adYc9nz0Su0
pIDWKf3mw/GtT7C0kUBfrYixlZ3HFRHa88Q9H8qCzylVERawBhcXI8fqlsyZ3eA+4pvuRTsuh0fA
6BbGGgdXZYDKb52srkAcM2lA+0DITTiOTZ5G856jguWzvvWkMZuAJVgCpd9mjIGpL+11T2ei/cW2
RJ5duiwreQkwd5SDOmiKjQLvNqhnAH/bvJVeVVWY4xGD1cFY3U/9TJId2ZJzskNTJZ7JT9a1hNIY
t8QAeDeg7WFJdtB9r6wEpR17AFmImFlnlRF6+lggLMU10OnxI/s8DQrkxQaTCMhVVenDcYGVd+mn
53ywrM25FuoDtZScrJ37NpKjMhMpVYnXqL7AaKyn2YmoRUUEhDIkQI0R1EcZF0lrAA4/4XQFqA2y
pUEjWQWlpBmgo7bX7ZE9aOUankpKn5YNhhnxXvqMn4hlkA5QUJ838QNBwTyjgxOv9nZ3nzIImb7A
0KHamlltarn5iqe5+o+uDnI1j8KXNAWL5fufdrkkJf9uZVJt8C48fkOexKvwo0GXNVO76OpGrRvJ
c/+4W36Ao6fiATlQrCV+dkaZJWm4ei4cdiJXQ/4iaaNnbsS4DPFLIBoo0QV2wozNViFad+DeKgWM
0HlS+wrOlGTEhGLxPg270QqVYZunm53jvttKBRr+PMxh6Ls+uyvk9eyqeBKS+Ba8uoRpAobA3/9Y
+OfeICd0qZypUVSyYL4goeW6LAY5OSJq/Rl12Dc62AXqtqgZPs/r1x1jEn0779dtokQNAeC6ViUi
mvjrJPoKAZ+l1Ep3p6EqU8fRhHIRYWcszXhD3jDknm9shk1hZ2XThBl/poiVROAq2Gy0Jn4tE2MR
e6b7T67WnIn/gDm02Zhc7nAj1q9E469V3onT/GcuHzaOqJSHKJBbCX4QLqSPWp5HOy+7IUb2RhIe
F9jGuDF4xQdxf1yn7aklnZF43vJMtsJ2zBRqF/zL+LgLhIN6kD+Pemg3FIeZkoXmJCUsM38hXkZY
i0SavPW4O4ON9C8eylJTtAQs8W6ifTZRyvK94MzISs3EQlSNw5MroXSn8jQORWk13IACmkXsbX1R
ThvK8XKEA0nP8OBdYqnaJocTh1bAF/1kuNm0EIHsGUVWkUT2PGyUjwnBrTlca8MmkwPBhbZKSH5b
VADiene9zGhz11LckQ+2lNvb/0OZgKOdvnVCB+46VCMHY9T8gTNTF1uwqSPiCX87rtYlJ/ebs661
kOtQhxs3YR9YBti/p5k6bTAGXzRCKQVv35D6TemUhnAzi/2Qm/iybH7PDiKmAAuImSYnE/aXs1Ms
iXurOOlXvX+kHHedMhHrGxzq8T56Y1aLR+6kHY4h8RCp2Mf+Eai/G+VA1S9CtVjk/d5YHA0L+Fgt
nU5JArXsmYEk3yvlMxOy20pDzGN7+bs6/6vPjbg3fTp2XqRopZe/4nXgOdAQhSDPNVCrnuo3DawL
tcNHB4gIKgAOPL8PxUnXLInJRzBkPDs+otoU2RAiNNO8zKYfTueGlxBiJYIw2pgiL/DUMb0qX/Pa
pi/nDun5vkPFy68zfVAW/eyOoQZEraUY842jOR5mMuXjBsIQ1kgKd75Ab6eqCweIdlk+Fk9VqpYS
01HVNFeNLWiZS28RUrIsGEXyGWA78VOqR5mvdf1xN9yaqa7KnQxQuZJeUmmPI/h+xhEVsY7aTTFg
9WAieOqKKve2eVhUqt3Gua8a97drTk03OidMu7+MTfIAk3S2UXe969gi0z6XztWhhmyPDm6Tvlbq
iJol7NzLxXuy5EWr85bvJJnIfp8t0hz3Y2tGkE0W224dUeAI2FRlt/RxfpU4+EoTggMwYMMeKjfG
7pmIvT0OMzkGO+dsaLcRw40lSM+VIw1Vk4kysj0W7u06pWtcsefTOaa3ZAsxXbXN7uGAIPaaxKbu
GFBko70w29b7sQlG6h+H/dIqw17nxbM2zFiSnFJ0t34nui1XdGbV5g6y1IVzp++1JADNF02NR/j/
LQqVogK6NwCufJ1Z82daEAkvRprsAjPsRmf6ll6rujti5iF2QbrHFA8+IsdA8lIirSZ77lA4HH4x
am/o7eH2KfJDO7xwfm2itFzw71hdnGHLLMKn39oOpPd7NM9v/GUIzipx/EpkOWBhV36io/UsA7u+
jf2ZZ6yef5jSbJOQQzOyPuiUJOsfJVdamJO4x/h+egfW9fOJ/LucAdKHhmGCnR49dqaWHLUUDFcH
rl0bdCG3eFd+ptRhB1rG8iaG7qX3IxQO6Au5/Z1gmtjkTXXN5aUtgejxAF9Fjfht2tRQ0C8ofQB4
s/FuAhazqU7nsoJ3y6wTyigix88T8bJueez6DX7fmSj8UkCrjgY4FZ045HZ6t40IcdaUqEm3OxPZ
21fAr1HwsBcU7m7lgR3fEdsMXl40y/EIPrS9yT4qsbZlStFhDc73ewPJo5Mq2Ag1ZtzW6XyaS49W
UfeiceCkf8Qm2XWzSXfHyUSKfUcOElHkAjXPooNXTbpIcCfSLIksxbhKhDBJETexBmvm9th8Mil7
YDW4KPVgIAU8xc9qWHLMPR3WiyJnYgPQ99QzHzjms2vJoXmtYf3SzRXbcvUpEUqw3AwB75XQW4ox
Wal/W8KDNuU7GijovObsfVsFLZ44P5dTGKEQJfwJAbLu4vGztGszchhN7VGopHGZf2/Ba6yKYrwc
ydMxzrOPklAGrBOccfrjUBPytWBLLVdB5/w9ljFVNk/gG+O28So/YUGA79tDpyb+IEmzn9QrPhbC
lxWO7fjEjaNLNcZ8S/D/mGKht3OowkCHfqKRK6Z4qT3y3PICdotXVVZApdkBR6OCgNF2Qgw3Imw6
EmByPnUgyWWYzV/NS+smhZjIPMxK19Yq5tlVd91xV4cegminLXpnxfjmD5Ycuq5J8qKSm/KLLyHg
mLclYoTh/5pejX2+coI8A0wXZWPpn8WPtJeNgERZlv/oWwQF0LKbR+5n+M7OFj2XJb3qsd6fEDDL
yCJVrtVNrxWrJdwRr5WUwedlIaGfa5ol8LNrXotsl00ZOYVTauoYlnuyNDp1FvNqlkUisaqXAaff
lOUwwmSBo8z+6iBBE6/uUa5oAaUCyzZo+CJrwsgbwTIW9hw6K9oadW8DAFmFNZs20IXg95GWak1n
UMlcg7RH4ill0R53V80baGxIDLiUcqn3B4qis7qoYsQEWwDareMuWoys8/DU9QWp2I0G+xfvDu5V
Z77jYNMBRY2Xd2JCnCbpdYU5BP+ENFfj96GMOY9dSeRDkI9TLW+qE8aZqSjHbf95ozL2MZE66MJd
fwBizrCrlYLc/O3VJX626Lkc1j0x9ZV9t16wMY+LveCNnuFlFZnphjU7fpVaJSiTlJPhuN8ciIh8
Y0h3A2CJoW+vmlEs88vdxo/iiK9U1jFwqcU2URJqd+n00XyZ807hoBDHDFdd/aymqa/MJ2lvTk0z
5ZpHhKzdUy/WbPMyxtFon2e+w5kNgXZMGgxpFjtXPwgky90rU0WJlY8vFHWDHsrwCz36MBCaM8Xh
k9ORxdYPxJWBPd19WdP2POj7nRPk4ldeBx2gq7d+Za/O3V9ComPgx9CchV7uzaw3oio0cyOmRmpM
4KDYOacmBU+M0Gj5AFTP5gl2lGyJrA6fZINu7B7ZyBKxqdKatjmHRuGl7HPLhueOuwu/7ZKYL+pE
yutaqA+ZonoS6tjYjYJokhRsctE6wD9Oq/KvfW+aANBYTzPE3oPGk2wDWzdvbvZiPiU2Cz8oDspV
GHemjpK/SGJusgGfVx7ltinJPEPnfVRfusHJMGzvy/Cp/baDtdbp6bOBL5vEudT+Wi8xe2ByiSEM
bNpdk6WF0dQ61IIfpcgYh2NtMhUb4pSSZb91AIglua6yaS4M8sJJS9uQ6HYWK1Yk9GSiScANHZgt
8qQpA45M+Pi7sxCLHeo9vmM1+zKb6l1fmzo78t3ItDgyLMMmqx7X5r4TY+2uo1g6mVkb27+vTzNC
5UvsvC9bkb/2eV2DD2zO0RqnL8/1tZWJx1spWPwb8Iz7Qv1VAIRKgzhRdIMo7F5ZRWGmHycux0xJ
APbhyEnjh5ABRPULazWn1ffVBHadkHIgdDGJuOWxUtskZlAASZ6TMagt3ilDBzx4Ly5NScwZcumm
+R/cfE/88Vc+S87Le6bext41KSHkz6SuoK8mBBmeNiZFidPwmku2zSbaM3mzMLQ2ZQxHaWezszVO
4GSyqYPfYujKqUGYPlGs5FaPHYBwU5m1qoVILxHbeF51zK048XMlBAgB5PS31F9gl8WPJx+r3eCB
MeKmf4tyx04Dg6wPZgN6tF+Nt1ne205Zy/84XzyKnPkEk4BCKXEA9Vp/8VFNm5VX+egy2TOn7mbN
1f0qsv9L60K3uPZVjIKHTWmKEFp2wph2oyPRI7uO0lS6gdiZN2FXmJkC4uwYnJwKrSFRHKLN1sQj
xrUbcsvuXoYWx46mI+osyQYAWRpKdPVa8R+wZpO6/JFlPZUrGBqQdPGakLW8AfWq0lTx6UtaWsNi
4KhpzINK9npKA57gl77Lc/KMcvxMVHWXqXYnp/tHcFQuBOPgel4bKP0B1lY5OpNXz0UhAk37wVa1
Uxb+A/uQC6YCltB7orEZFaFDt9rCj0aTFhsPSHxozaUcdsNM/YiuVS/rH8qxb4e72jT4LuQhG/oX
UgR4yXo4n9PhxmRK4S4Ta2yFylJY1L7yI6ZRSxm9knVl6u0cJdHvuMP7/3Pi2Dr/Fr2dZg/8L+Ts
9eAHak+u5Lyt9f9JQ/Ls88WR6q5QxK2AP/vAsaosnXQPPN0/q5XJZZvWxxmhiFv/wdKt9a2V3jw3
e++7NbSQo0SO7LOpqymn3ihIolcpny5PhXw12WWoY+T6BoqaEVq9f6ajOPy5qCOdQWSe+hK4RRRj
NKLRF5hEMqkTEFIm5LiHTjr6f7LiivJVd3A3NMNc8JwMEAQ8AwsGrjlTT7Dfb62GOzZCk6zhwSi5
i96gcQZBp3QTm2U18rp/yeKmS6+xUXov6SLhaMXDl0t3hPukvEOI6a+tel/kbHQYOaXIjJXKVyDN
ROkqQl2EDu7jPkMZVlZ93drfS2OLjqMeIXenwLlDDwS/lhkDVfR5qKHxDp+objUU8Ut7rKd1FHvT
de0d77Yqg8faOd0Uy2gnVf0dfbrU6PFAa8DDCL8eP6wJvMZC7KcPvdKopRCc0hb5r6wA0QQR+oqY
c7OgppG1kEkcFRjNxMAQXudQDY+OuMokAOIKtIYJfKenHtHRwoG0DQch7S16BdrnIEp2LDDF0XGX
aJx6rdqfTsIRYzde9e/5ObWuhRp7woW+PfrK0hzr7rYyutzUnQXut0RyoV/tYoBkT/GjyE6BqEGh
5VM7JyCExBuyUe0glgi8w52U+a0N2WLEhQxa/c9vGjx7kceXxhT01XY+KDPLr7dZFH+KB2GparmO
BzmDWkTwggfCGD39+vRYMK36q04ulbkFeKPhzASseTlj8E4IxF6Aa38WJ9EfMjikx3150HX9fAkk
jSEV0mVOlKDsw9MEyMpEG6p043tQpOmOcjpVVQ7n2pru/dYD7lcuuu+RVd+4nNXOyOyX1VFe9pJW
s1CyEVQWZrlFTsW5jyrL0BqQ3/GCuk6dAAOTjZlqz5N2mHx1OPpyqUdiwom5U/t2ellUaCdThEim
seoT4TCGB06nLSIg1cQIdRTld/6E8+uJ2vLFjAcpPP5F7NMVoaGcRWbtuT5PkowMRRVETpehdums
G5SA3WJG+pbjNK7nywMw7c+n+DlozElOcmM7t05EYwm2eEPvmJXk+KjUpWo2m2C6C41jukaqS2Eg
KsF2bu3uDC40Qgzv/NEOOBATZXQHIhEKTX/WFJRW0Tv7FlOHSQSAZGgjxQ1YeSwzxOVT1TPbgr7t
XS3AKcEU+3lJW58ACaSF917Yf3EGzCgtsSx5bD5kSQzjrXfXm+zkkJhrq/7rDchoWzBiheKc01cZ
u35WtBjfUCRTWs6NeVBOpMejqGPHb2HOMY7eI11OVSfMPrznI1NYEqnkFBtFZYGyV9UGu89GeO7d
4Xpt/fCnBeO3hDCEw1/gZJqRX1KwMG1wov5qbOUka9S7nc/RsSFu5GWIhBxUMc+U8hGEJerysvbw
rHCAKkF2Il6wpyYGkDp7ixfXR+0KXtj7aDS1bo9i69MImvKBU4Q6h0Q2Np4GUuDwp0dz31Lxq/4F
xLzmgu29TalOTgaoPCkxm9z7VZ+NkJvR3KpNGqww2Er2pkImhXlBrGeb6vHzKzkv2lBM6zdaR7ws
Yb9knzV+8VaLVQVsxbuDe2eOgJscmPH1V+iGfIX6uuxUOQerMGK8+qwG+A5brM6jNsgCl5am/YDt
Z+Ce18IuJ5R20fwS2eFo896Mmogem/A5XoopclerZIMexMcHSbLMuDDaPFq/Owit4pohD7I2z8UC
7VD5zPX1sZ/6juu3n6ILfoPhvqLC30E4ZUmQX096bacHU0g4bW/B6iOD1v/jMyG5aAdS+h86Ci2f
urjAyZk5jClhGMHdUD+eszcg1RXjfM7lEL4oezKgDQ/HHplzF3IPuLh89FQPcborMiDFE7S+VLMc
p0P5VNzYIJ6JvU04YwaBViprMjUDqaDPWRFb2SYAzyzaSRRY4F1RuFBXLZIChBkqQ1AoJ4gFs8RW
+olgUHtJSVxqOUzRq2MoUtbcxekj0YbO8nlBkaE/xLLUTAU1TdCyv/RuXkJ+6Icofkb/b36qU+oE
D+UALina8FihiOm3zttTVWXfI9NlA5MRm5OUYRgeut9bcYmF+tEVlSW3fpGQmproNLMBhJgDpDH1
bvCX4rD45rDQPCiI5xSlhXDtG8ghUAnk8Ps7hIJ4QgN71+MbelhqcufDW5knIu1Z1Y3UIRBl3EYd
Z5Y0qrZzgdKYWTLm4ORd6aNRhdlTWpQ/2kXWm4mRKv2zzYk2f7jY/sffWYTpk2FzuE7FgTmvvWwm
N1LBlFfIS/WHyX6YPn9jvfEDUlrpMo608jkPJLwF1UgWgbJxCBgKJSCjgnBda7K199eXmaJeeVze
9zTTbidpuqMo5KHcGgq3OPIg/Ggk7AN1JnwzBgxtSXrLMR4X6RZzDN8rC3enxhx09WaPWmS+KGwY
yac7RK1UnyaCe7SD1AAdljqWKLdF7mBuvG/7BiiTb3R2HUPU9+3HuScphVsqGwt8UBGBlKf2dcfL
k9D6pA3Yx388IiWWeY23YS59Lrg9KD66+kHJrdxUj8Ipt1TCGgtexj2vLe5nUib1Lh/GiLyRwv06
T6klhPV/Nk/TBGmRCwBHI+ayZ/NFOEw7Vslsws5wGrUghLb4gThVL0wTvEgNIH9gwo2HNsZkEV5P
NRolCApNa79bHqn81gByjk+eJR2qFxQFsKj2boqe58p3DsqKIloD4IC1oKw9wVSmOO8/K7rFtdb0
Vk5y9Pt2yLFeoDw5VtMvcBlIcANhZqa7/Vj5AR1v9NtwUBRqe+KlaV6OAPKMcRkh+TYPHy1rZ3ET
lxF69xML+mvXeqHBEx1MmpIEwe8AvIIh3r+ni6m+QbRN5FI3Jb5hB+DH/vySIf/V1ig6+ma9ONBH
mAXC66OwxPu345vcObfOrJ/wLlwwtL1C33KmD9ZyhqY8AIH5S3sV3cNOoYV+se9SlUj1QgHKYDX0
6loYwJzuf97jMTsJKgRHZazsxWRyv9gggjQ012ITMRzFRqOxa8shnNZxFIOf99lpej+VYphrSeyC
i4rRTWOmnRnwaeFHpJuvNGYb/A6O9ILOl/HbIQ0UuHIWLUjXpq0cmYTcg0Egl2XCDy3yGFNK4ebM
rkPrpGP8dlgbSHZ22ElNlpy5r/XZ+n6Za2QlvpYWA/uwQHHbQt33sKLlIhs1oNgkq/sDyAMeSkV4
dxZZ3rgnbdFMtuSTsHkqegb+qFY0VjPcpP7YjiaLVzpsnIR3O6Kx9J1PhgGhUKyfsdhvhvdvQGm3
etA4ybKdZYi4UmEUT4/11gQxIgVX16pvBS3RyYvJMs+WXujjbEimhPY3DaMEQFtrItN6pXvb5uQH
b+C0L16HY6Nv7eAWdrXYrKbkCIrJ8+PSOwldy1sYGAT9sC96RIoYjFIAEF63DpUYbwA8I5uzmDwt
cd5srJ330vk8/ohy2Ch+PutMhU/KQbeVYN8/SWSFOCyNbaXAPJoRvCPcasJOKjzHgwW6qT05Qn8C
6iUQuDJYEZUNnjW3s++Y9TBfHVqFCMvyo2bD5iLc3SXczHsciueZVd+pA1kojpu4H/N8uhCde9c9
M15WTvZjILRKrFN3UnBY4I/S4wDivvC6xO4zMnSKsbCc0edyS6V44lnSeZ6vG4GQZDvRkN9GuQGi
d6jmsrSSOVVpL0pmN2UKK2n8gO3mmir0FJhykIocL5mfQkGfK5Wck5/PEZJE12gYR9GP2f8vqBwF
smb8SE/iuelBDublqxoLtVkikKmy+RfkmejM+IVDoegBXNA+kIo5439vaEVQ9x/5E68GNwlGhBX5
S0/QKUChm3wGPnoo9JfBCXgkNnw4mrIf4yvYTzZiR+xswsmUBCBQ6As9R5WO0bpz/B5+riKl6QcH
np9XeCR9z+q0QF1I1HaRCG5sFmh+ywR06K/LHVFGmHaUzLNl1TVWN9rvEcL+AuKhkTT3SFbg/mZ6
39kYf6gCyKnO3BTbitdJzTYsLosFErxu6qdbUSTMSkQev+9zSSz5b9UmtoogEFp/TLjmjeNYetkW
DHsciR4TUolqsHzFJGdF/JWBtZTZDEPGElOrOG0ROXllFnSe2uOis/SRTlqyp1oSX5NUgECCuWq8
yhGLCYdLOfNamHgm7HT7XL+R/Nvo8fmRoBSkqZ9KTSlb+EX7YcZO87KnAgHOgeP0XbhGQ7Wbk4hz
wDqx0v9mvZGy0muQVPKzh3YRJNNE/HUOyjGMNWQUVMxXzi3rjlpeB9kMOGyJrmn8PmiUrhGX2amW
7AIRljCqgCzYDPYbNv93pqNZRYHI7f2zQFwIMB2d7aU1RKzdyDhFnAIs+DWUlH/rjvXp8ZDvApIc
R51MYPEGGqc2mrH76Q00r5SoQglpO2//5Cyo20+NGi6VWIW3MwghznFSDJYJpzcgcOl8W06G6Wpd
XINwxvHksv2ocY0Zjvzpqnsji6o15myDqDQMXV0bT4J66CJ2MO6dY0b3Vd81tKW2XDI5tbNCr2vO
8rPE+++1uLGbOKEQq6Pxt9Lfq/Q+Ddn03MDF1YnNI2ZsAPESeSasqXRHgyl01TwuJElKBqFCn+5+
YhC3TOtxn8gP2ZGtaWD7PmvKVsx981/ldhKMiItuLPE0B/sa+GssSXKdP9WEweNn+ZXUb/kIQWxp
00CuZMCnAUZewyqlOgC1FPISMR4v0TTJ9jptzjwk/5MJGjIDfaLFu/aornRGvhTIvXNFCe/sRlfv
h7cW6DHhaAmSCj9RDm5ChEGEUtEVtsQ76MApxoKSfwVdpekzPqbe2dWg61ewt0Hrc4oyPhg0X6oc
jZ+mk30eXOQxpB9j0tUhTT4G2kNiOlYAaiETQYda/3BTmwzOR/B5m28Bv/meA/MWxozebpOHV5WG
v1/fNXgAb+lmuVM5XV90mEst1UqpZGLq5Ay/Y+NOwXpFocacIXJzPDosFOO2fJqnv3K7Ei7vi8dN
Uf74q2lvRAqiZvgYvmeRA93DQQetRG2ialjiCf3FRumJx5ulRw+IpL9fWp5kSdb9EfWzCV8V+geV
txEde+R6x+y4UCrEr5jbwDhX2J8PX/4hTpXpvh6EjVU0TQykEn1H/x5b1fFVNBNcvnb2Xb7nu572
BSB7yQQjPJ0qkgv9W29m5PaWJRBh49mXernDc+ihwrAyc05HKa8SsutWGulEcowFZ59xHEy72PcL
mAJUzVq5b5YrMVaacGE/Eh3dMD1X2mGjPuNMVa6J5WILf68kiCHIT9DUJPk0EZs7fpbK7z0rRBk8
fofaphDupzwIpv0UIv7PkFtvoiqsccrqMRj1vNLxkSlZcheG9Q8G5d51cTLZD/I+1IvPy0TUnxir
m2pzc5qYaytTBQawX/yGEzyYFSFaNBnLCDv0l3/EByuJnl0NbQa9TR9ZJNQJN0MZ5Kgd5FhvmDgh
eyJv/D186MrOk7S7+Y59x5N8sTy8bWsQWumnlIFY3gOOC4V5724xJjMfaJJjdAUqF6A9jO8Cfg1z
pDgznnz6V0Hie9pTEvn/WomD0Vl2hXdYhUE916z9ds5/j86dlBT0wshWImWjTZPlS1UbMjrMmQXY
pugrIWSIv/Pe0OuU/Vli1Bccb/aO9K0RgoQroZQw6yHbbG5mUyqmTWGKA1o/rlkYhAuKaOPW9iCe
AsR7QPWkNya/R9Ut4cVtCcyuWb7EQhBS6GASHsFmfAFgHi9VEr927+S3cRwVa1Ek1n1Qg+3O+IdL
Z5cM9O2fxKuoGaliu2UgrZv/pTDokW57f41sjKAeSLzR2mQRGfhdzlXQbp4BP2nTfv3TVQne9D/J
EZTyfOVogq/LddMuyx93dhOmjkESbUupYwy8RpEkds34jHlV40yRlLJeKcf1/pCDWN+/P1pK4dBE
iFUlC9yr3QqjVKJ4oVdfR9Rz4aqYZviW5pvExa8A+t6jNwNl7734MN9dk747kkz4rWZ85pfl0jk0
FtsPrya+OncKRbw9eaon/HzicAFBmvVuRqp7ymgJ9JWXRyW+MBsSLRrjYfeZD508oz2CHR25eITG
jD2ldyxJHClAichB1RVfcTzzV7Qx3fVT+cn7LJEddiCT33V1YONCjxk+X8JlwI8h0WBKkfhSo+5d
JQKrG7iH6gSR9lLoyqcCx775ewfBBxbCYeYLlcLzcayajerhY7OAP6Rhd994IMsIto+TMizb6ln0
+G8OwGkbcH0nNaHpidTUoyumM5tyfAkelFBktAfytgOFluxzyBY2Hj5a1uehRSH3oHWSCuxTRmCO
MLkcwhNCa/pWzfq1k0u0OM1YQmUYfNQ2Vq48n7fsgnj36J31mvSy9Dv0ZUEnV0HxMsoBIq3ozBbd
PVqYwfnrx05wCY7yMcc5/zXUbmNbGL9URGHgYiGNBCLsvE9doj1A9SBCuuJqF7SbFU+FRkH+2Uxs
oq+gjGLtPzGgjRF+shw0CMMDazhS7kWG//ps96sn1VB/BUXDpvPpcYaaIs+Tko0QfjCREFgNc4t7
AuGNL+HsmlxyCLgxZuLXPiMpOoKktc1pNZ1q0m21A4IWd5oxcCLjYsYN7OOpnvDiwgpO45kCl/gX
e8S2KdhY5K4rEXx4Xo3RsSUd/+mvIQqxy4ln5cui3MA8FFScpTzl6L1foIci45raVBtCk8EXMw8M
GaMH+4XeZRj4lQ6p8fPBBH57YT1w5NzsNdWqXPSrWt47r15bFG9fG7J9BMPyoPoxzqS9T4nV0RsH
uXjT1n2xwPx7AhJXtGJVkxGwKEkOW6VBYTp+ENRVw3Xmew+HyDxu/0LnzmaBhOeGx8kxkNDJQF7O
3f7yIU3WmNACykHwg0LNojTriDwtmt3G5HEUToA+m6vmy6XGxulAgjg1HaqfUDEOUo5aCIqtdWwu
DFHbrNLs9eSbw0sevYBxfJb2Pa0MrRMw2YkpiHlcPsp/JKEe6jtBRKysep8TawFAAM4mdDbRMuAq
HQrkIuVh5OQVyyzOCFPuTNQ+x12Jz4Nmqj0W7pYGRfJTKkSC1ydYGzJRK6MMftDO8NiN7gTnCbKi
AcMNZx9VkyGdf8e/hF7h1qPiC6j5A8KyiOhX8kimgv5RfpI/LUPWT1QBH7ud553nk/WC9ePqQPU6
AN0Vu4l0okmUlUvA7ebkp9IGUgbMjLDPolpkY1VS4SPRNE67pD9rc/Lw42vpgbGJQjz6vVLYEMhd
yQ3duw1Uqs9eoQekXD3pdg2JFOC2ipYV3oXey+uSfdd8cax9UQ1yFCwNH9yXavsxOemuwxaLzWFz
CeoV1DYNDvKi+AFaYQZi+hM88wCFh4qg9dYLuT7AYuQwEvRq3H1dIfEpTUckEEoqSphlA+LNikww
YU4MvkVKzRGWO9P1IILOTSNwxIGFDcrmJgsFYMcTRIVQB5YmzUjyKf7E1scLe9yH2vjR1eUz0hyN
u5pK0ho/gXOdG6yA6iC1gvCEjOtz6nf3hsT3I6ffAiVyTTzH+4AGzFez85l2+O9/x44Vw3oeuW6K
ZRiDxkgj7UKP/WRGp3+yax5fGUpmdY+zjiLRGEZVw3vcl9FJ9e9GucVKciaU3AGo12qZop6FYihN
N2Ei3/splsxHqRSOJjId5s0mhhdaTYg4bTs6no8X/rHVXXOpk18UZPYK1qxE+7NibUMy7DFZsvqk
upgMYFO35O5lJwfrQiruRo3N1mAjNxPsVUIZl3o/wQc+wBADcmYoVfcCXdPKIZJYtVLcy7fmPHZP
K3KvfMnckHbcqBbvBJCpzax+SmZ33VBE4WnHN+a4BrHdJBDvzHDsqnOA/0Pkm7YSCj2KIsgd7iP7
ZfaESobH7N4q4y4mNRCdobVux4/pJqX6fyJote6AXm/I9gw/T21NA7rhaM69+ULGh6kFAvJp9vaV
3UJMc04Xc3KbvMaof6J9fSS2ckYy9GT30qTS6qYgCRJRRE8N3rx61dMT/0IEVw8XB6XS9LD6AfB4
M2TDtmznmhfTN8LyKuIfJ/rusqArJ724CxfOEq1DZDTCM6LfZ5/0NyKYhid7szPOH24aorZip/E6
2wLGy0r+u1x2ZMPQOMbijRF/7eVTexRR53C2kd8oRk/ByJ6LO1pIB6h7/lW8nS0AQdSLitS1jh1h
b2l1UosTUoj3lCkPNMxLelS0wbpPdkUOCsl9jC+yQ/DRQJNXuNBJslMrtPu5C3rDiM8H6ZSF2ETm
esMTbs5pcp7RU+YQb8B+HcbtoHQHs0TRgICU3mXdKnL31FHdTTdEpXvQevu8TBdbcFB0CuHwi+WQ
T+kAQLtmrSyd0xqBJjFYcO/Nu+JkwDSo7Gg9LlAMQTBMDtfu6JzGca2GqJhh4GSVzsQgq8NiueRY
xEHdt7ori7OtXaIjsZ4PK0f6Oh72hQVnJzWpyz4MJxdkEFONdkBbICu/8eEDLwowkORcLaNglLkz
R00FsObW4rNV6fUlaePdVSsi452aZ+U9PcBgzQ2jkEX752sPmGG994ewZqVidEPLYpLjch17XEeU
CbH+zxw4A+1yb4bONnzk174T04TGocLSDVhMCNctqD5BNcBj4+bK2ZwNcTzUR1bcsmt4WZCdxfrI
ZLYLJAjUPpPkVZwSMY53FXz8vuKlWUQBLsYHquot38Kx46TDH6kGsEOfDXTV1Mo3E5OMki/sVHUj
nfyZK4iR+jOb+M08955AHmrHa0bGzXNvTceTxrDZTxK57GVbNZlnQ1hNd8+RZ66iFUtX8oWFwFLA
JAWWN7ip7uN8nzbym7rdx/8GiMWgN9zZ1xgHuSfWxwGq96lutQTGlLka68j3AV8kBJ+yI4mbs21f
ydppxZe1aryCeI3XARx98XZN4hTFb3ZvFNpRs1P80QY9cCfz4IhwOQ4W3XAi1m9G/77TPDfEbkhN
OSCP+14qssIt3PqP03/FBc9+8mT7Gno0teCvVKcAvqwF2bOZMXVStf9DMjb7u0jqLpi4wlE7VcsJ
LZqSJ0u9NOlJn7tOunApe5DI/7z4P5/yS+aGTO/3QtdvDedel4602/hVYGpR7btGb4ykcrzEYLIp
y2TvQpLGFBQDxtPI2mH7tP70w9JCBDF5zGxBMdsuydCKb4tCyce61FnIszf4HcgUuaCS5vbTLTN2
4aeG1l8Bvwy3GxPtqXK+h/Y+0m9XKcMb8BrYIsBHsQnpD3DN2sS6ux6aWqsQ/fS4RvhMtwPTHt/F
ecFNTmBOIhoe1eF4PhtYIowifW4jKyCwCjxgL8g6csotlcy5SXa5H+h2kM4Bl7ZYUvQ9DhNPH7qm
kKj9s/H4TyuABdLqDgwtqK6/QNlfF76GzWvCvfzoaoWhZgDnnAazybV+XElxGwrh7TBy2ydLBc0z
b3Us62/8YYV432onDqAfTK4E9FqGLrj6LVkSHI87iLVdAKkoIEv0ffPwno11GRG7ATtnZOl2xtKq
YRWp10XNUGcU8jBXeknmE9jFLYtKEmVBIBUwYSKzWiY83bjqdgw8CAbZUZ8LXAOnBjJVTLGjdrb/
0WIGbu2FTl+oPoui6yIKxf9usByuXM1ECArzc2A6449+Tms8Qwk2JNYrUKoua2vzHZUwa3wImE5X
BwPOr/vl9G+X0uekLo48IE8H4pUZR3JsfgMXerzy8HashBNnuAASrS9L51ZZ4OyHzmkKIDkoP2Y/
GzWZOsI2bHP7ICu4kb8fgqkCxLDpBkV3FkGP5AcElqdwjCWyr7FraciX0vuMUYo+3q8T4JhaaHR1
dQQ5vpleXBdAi9rP6WlXTOGc8gLU+bQKTU9YjanaMirqPZs1EfKvNs1RYVTU1vRUMt7jub9kVjDq
Q6CdjkNV+qie4Rllg1EU0UyTC6q99B7VDU6xq5UuTdVCNkrvFSOOu2OaVL8M3ym3CiFKBiM6zbSu
b0qdpd3zTGt/q5AXEBPMnECXGfpNj0Y9be9txJOnkaOitObX8OnxAD6AIsfWn1pXjo+UmXSvDVDw
EOaJBZjo3yqvvqYW7KJFXlziD8q5YtgMmmQPaNW6i2pxj1g8BQTRjDABubtJEox625migMTCBWRH
rq69OVaeAMkfALeLFBsRLg5ahYs/jvDyC4ItNBcaFZi5csHKqKQItdjWmpeufB4SOEWsE4OCKBVR
IR4eNsxm5lbpP+rsiBP4+qUAZmuK2vvHepOwccRllnbXQQLyAjWGH6X3uARvzOyYOXsfs4MqiTvC
WnZ4GgC6rvr53maomp7rzwX8B3aWDg8D3oMaZ4RcjL9UpRTpa+BdlcIuxxpRKiHgQvWDpZUpCQJE
s8egrPj7y6vOPtmlyHoVH6F2+VO/my2GU5/aWvsFI4K+g9Bs2SfxgvKc3/QrTUUxkYh856MZIomo
3y5NW6CcQ4sTxH++OebqkpjmjLibYOOh2LDoTCOkVWpE2/+V02F6Pm1F4XykCWMC6rJRqzGrPSRY
XXPKX6guWyVmgVeDChrBXF2VltmZoREadgkz75GjDAhjLTqJZuRdU6IWAKo3ZgnkKD2b77TFDH4y
Rd5h+1Jdqtjpj+47x9bW8bPa6wWlnNaYjYDMOXZkCyiRpeUxm19qnxjhvXSo2/DjavGjANpy6FJ9
oT3icFPcYD3EmV9USLt+b+XgD+wKCbDjotuyU8xSXswenN1v8UrMbgbY2xBW4HNbmLE9AXknBsCb
RAiisAaKRHu2GNnhxAu9wZ368hnajs6Usep3A8E++uHoMuaEEN38jLtH+5tqDPVMXYesVta/AgVx
jwvK2/FB8BC46o1pn4HUHG664TtU6QlU8d92+Mx4sUqxfHCTPamKaQOs6l2upM+DZWvst7CuUZV5
dknWteZSnObUczagH2dR4PzbXqvXKfCNbM/DxhSDdj7Kstk2NxeBC5VnKYNG5X7yM/Mf/Ide69jQ
I9AfAvWFXbiNg5fZ5Uqi4fdyikWB0b2U0dp9My3dGwRfHueb3Jj8ViacIw1UsVTUQ3j29tUmbVXF
POTs26v47XrRQ5Q41ZKaE3ghcViMS4cq19N74X3ORXIonwrXl5MaX0R5ZeGN/yT91gOF0/KbqFoL
h/aOmy+7bideBaAIi7RcaFXg/j0CuJrutGN1oERZLpp0IJlm4yLMcs5vMkWqe/1LFLXfBuxC/ADD
B3h/SZG8Oc25Gaenz/sDlvZ6HxIk4hG0b2Gd2d3iZf5B2SW1HtgOhZcfDVB1orl/V7lnkBKQsKtw
+/vNoNoi3VhSpuKBPS+FGJGjXI8yrK40eVEeXA+d2PgAPliozY+t2MHnatqM+YDvint4edSNl9Lp
+BGd9aE0dlsaDOrW7xfEX8TpXYhKPXinv3gUDhnIBV155dsJIKo+ESdCSpXgt4nJAC0eXCTnfxyo
lmHKfbjlzC4mlc1OwN4lyzYXVQmJoVWq5aqjiza9ouY/uL6Z00IsMLqgRNrOe7B9BOnoZGNM3y9x
Nf5ST4auoG1xzuKFKgV7zb+xXX6DpzBe3Wrl0vXgWEma0TmIXzbuqtCWBDKYTbpwrF7c6Em9wB2K
1y6rnveR3hB91YQdJwpxYnuNWyZNX7OAkJR/WgXvWnwdh0CAAAr84/Wu9Wxg7pCQwbQPhrYZI5SS
uFWEB6D4l+p3CaqSfJ7ogfc4y1vuc/bnaGr0iStAXn6NgAw3dHoFiRmbxzdkI1v2IDV1tNdd1Jh6
zlM3tkDICPtmD1nyAL5cqmm8fmdJsjRYB2IxuT3z8vMN4pmmcBeV7Uk1dTFG7ld01U2yDqamJ/93
l9jSWOsaRhXNZJyPKiqZ825Td1WrxatseNAgtu3118xTeS1LRaDvrRFzM0oz3FGjvAwxg46LqkVv
zSj2vLQ5T5X0R7pKq5jrOTo+tj1PNMSZkG7rnQHhXxeASfW60EYFTaha6AFP8jBKCHXjWeRm5TQ4
CLwtbfZbWybWrqAJWkATG+cRbsjo7KzJlPiFGD9IdfxM1s8pRTPBupBjfqBP3YTLWLLKfp+L/EL+
/2obQkyyotX0DfxE/uZKBc4GUk/dPdEFLz5JeSiu03mii2qpHkMTF0ZHJwkZ5KYFqOuZ2Ss5uOFa
lpxEAHlt2EdEopPyNi94CEn83lIuEheXvJYfWhr5j5AxqFXNKrQHWjwGTAs8mk9hwbSLyhGTeo6+
JoGVEGaTi/ah2tM8U2PTsWT9c/0BFqw6CxbuEJ+/HPL1OGy8bW7c0MuPAGbjQafSV0j1rDRfbrTR
MpUJefAYZ+30nHn3DAM6k36Mt6prBKXVcGSKYO1vZkJzI8zm6onyUMsX0uWQm1O7xQksySAhjBLH
Tz/Fz4GLHJkF3G04zqq0vK8xd4Yg+LoDzaLOnG7f1G8ldLvsL3AIZc2aFUvIhbld8MnKxRAjR5HJ
7RTxr0xtuyy4VQxUXWHw5ovF54L4ItCJdCQXf2upub3zPv5E66LuyJn9dSLdmeeRsdjUi6UOcFMd
mRKba82ao+PY1Ww0fLjvXtnFtmfHES1o8b9JuKQ+xUEfLr2Xx96eOcn/1+NFn1XV2TKCUg84De2B
zX/C5tMt8vnM9atRw76ba3wwnP31zx7vUSUW7bAoEAlMdLDuxW6SEh4ms4BlInTmhAGdSu5deaku
0OwTEXIEsVeHUihSCagwbgk5jHvoPDlgS/tqg7Ow8O58SQN0gVG/qdzvs0abuuznbdTFyad/BIg1
W98BV6dmKcse5LeDJT3oE/u0ldTVEPFWjsKR8EaCCreJv5uN+Mej3QTvZO2rXLkt5djdCLx4OT7J
vh5MW4MG6V1RVSVzpHJ7pNUK4KuDnB5CaQIwl0y7Fr4qK3cuGBMB/AKkHhHfWpBv0u3Xsb710xCS
zWObKto4InUZv0LIWqnNH2kN9oY5/xm3S0nGGcqVxSJzNVg4NDT9vKBI/RTmbek2+bx3RP4XmunL
qZo0POx6VJEZnXS2VBfKZlWbcUeXDt5GXebwJ7zwRGbmipAbNQC2JeeW/dCUBE97iI8QPDLlF6RE
BX4ptuFhr5sRy938dDOCUotIr3n8gB+ns8lsVd5DJWuMxYfILTwbqSQj7Z63RbWrPqMxW4mUKd5N
eBCg4JwkMMDSuBLDA708SWZrY5VWNlts6yNNjNIljojQVwu2Opqa4JjnnydV7TdKpdSPfshMnI0S
n9Bh88IJEaFBrGEwtWc3r0Fy5gkmeeMex+519ohke+NzT0m0MzK6cDcGUOPUgypl7F9/+p4fNnFy
Z153LudIPkzrl6lmO2Jtp9b0Q8LYN9EPeCoZ2+5vHRubOHJ4F1SoHGKWy7gvgefteu9F1WnnWoKG
brKm7rvv676NZA6TrhWZvWnQnh4wa8yvBnTTGwmZJeKOqKv1o93Q/suyno6fsjETZMUFcLltdqLS
u499zWeEgbIaM7IwjIEeX2xO/ALwSilR2ZN6ToImovF6XFFmCgY/cdPBkK51ymNOvoR8JYXrCXwQ
EUP62GZG173JDvZu8qdpoMM7xnHXqw2WbAXzA5Mj3/+8+KPvR+yLruFqkzSWBxPrOWEfIZQ37JcF
9SMx8Xrzy/p4m7fQmTQFN8u00kIbivRX2INJTpd1PKoSKdMXOTKPJ0WiGbxx9LSb6J5XjAGB8g4S
XvaLeTwQk2BJvtWAmh8B+X/3iPxDIdjzUZuf5Fn4dSBYTRmOyRKmcy0S1zsY9cHkJytMVFlyo1EL
S9789mQl4JGvoi/oSxBOPWbQqaUDaGVHPPKWrhoL1SzNy/vwVie31OcXDmKVEHBGpdM35T2b37cH
S/ZyVsSJ/coKYr7LHTSWw2CM9FcoZa3jPt+PR8OtXcnTKv9HMJTxgRPvxMjiU6+uuYo8WYOo6eju
s3prOqUhQlFjP+Y+oL6uGFlmwqMK0nTcAOytlKr+8iFGpIjzN8TGXmInaGJrUCuvzKEW2AGgrc9+
GF0qA3f5Vzx68fyRHcLwGQ3v9h8zu6kH4E9iazBLLCDOZTVInq0R404vv75NxL7Ciqq/MwFFLn41
ztfrui4WebI3baKOd8vhDGcrAthsbKXq/ScZ/RkPc4EUYVRWlhGeI59uLFy8YNbsN/XDHmSsGpl+
3KGWYiEfHQFOj8A82/RwXOsSbeMrlD24A+U+VxFiY+mYP1khbf9j62/fsOtp4FJHnMshdIPDOlXd
+vIVrPlKi4/wOBIj8vjsaN569LavuUozMhpeEgw90MrvWHstm6N++/Ws1w0eeUK2a6iA9l6TpeOo
7Q/r78s8EUviS6NJdVCDj6+WijDaIcGmaOjE8v9dmYrMsqQVg7A0kpLIL4CQgfzvK9zo0TCAPb4s
8yFOBipU9WZCR0/4eLrKpcyGrSH+Ccnpzv7CMSmxE7FWD9LF4h6/8jZiaPPXl2U32JkXx8UVEsyH
Yr1xBiI7jEBacA8rCd65EIPlIcLwc8Po1s9ex939w4eMjdc6xbv73T1kFWfo4aVUOttuLDhJFIb5
gOGHrwamzaHFh+iWZcYbI+U5mXUqLHDc6jtwM1MEEaKSWSr5tn02YYZHSKokhNE7Nuib1PiXOupi
xwVoPpWTBOLjGfi7VaLPSgLEWvhCmYHPySyHW/y+HdyGarHZKTek3bnmQ2Ve2FyvSpRaOHBvAhkL
xeL7upvKwBfqZOV9f6j1yThE1TEol5/Sz2VxhSbcIJlTjo+cq21kzD+5pL/7hHcySviGTmX3I43z
7H+d4VYN2vJRGbkah+Ub9rSryy7NF9L5BCekfwhEcodTiX/lwTgZa4VXP75aw7Gc200Rn0zynfMb
EBgO7HzD0JQqpmirBipzfE7c9BfU/QNau6wzlxogiCxl8C4glaD2xq6umBVy06QaBFfQujCzKeHL
OEa8dJKvY6Xgn6UFFhBfZBK9RrHq64dPg8lauInxhbRVUlWfZEvGAG+gaQlpEGhaOiI9BfrESDgk
ysDIeQ0BDPLtNXsp0G0Chq8bn4taMnZkF1K54jWkYvjfC8KCqB2NfRRMCpZ5W40RFFYBs2d4C8GQ
cNqKSE/ihjMVyyKdp7+pb1bYo2yAGvQ5xoliR+dssJp/CvKUN/UnUUuClbe26+OMBZgUn1/vgIsV
0jaEHlzwfvGEI05fcdR12LH4VsvwcoHlWMJ6XfpdZJxL+lp8BpdUr51QuzjeFa8eJC9uT0tC5ysO
usNI6M0R5q8BKr9zaIZwwjdxjeFp3eua+RAQgJ9A9PmkWtMs9tiKokRyO27wqoUWlgvBDhXr90Ek
7PSTb36jMymam0A9LMMoy7jxgs2Z6wiG7aS4LFyOHiMdjqU7+axM4+VNISlxFHLSdsUKJaxW30kq
AjrweoMxjhDakt1jyXmHvhiPO+vvPB9KKYdWURpIX0mi0cSw5gu7xVQO3t2NgMThUlSasTy/1lcN
F6RYxl6dtNi+MJ6axKIYcCWVCyZDc19uJvepmydBniNVGbQem9SwtrhmTiqIBicXyB0J9jUV1VDB
4hucmFKf7fShvcyiVmRAh7aZO6qMX4987vZzhHe8bizkWDfTtdML1GTTVAsusJiIwnL2E0wOvOtj
KIZbecZXDvOBI/a/SxIYZF5iHrnMJyzGF5cP6ubsjuSI+pqSpClvGkozqJDAeG7nmekPu4/4Kk7n
NjvE7q18x2+ZqnBazvdZiVGIh8Gspr5Aj39UaXcqzAcfXV/vVNq15m6PD8uSWE/8xmFQdGLIubzy
Q3nJQOdisCkVdU9LEzYeT+J2Inw/jXt0+Zsa5zQXXdd0ukN2eq9ruNuVd4WgLVhqjWsaNSoLb2Dw
I8r5RCe7VIHIrbTRiz07i6P9mICQiXGJW/kIGiyXQ8k1Iu2zThRvTKXpJNLewj7+q8eQ5oDgD2Hv
rawez6MQfvOxEoae5dwQKBCLg7ca2JxmXFLVNH89OLBi7xDSBMqazT0LFRKBHhTB8Ku9tfV/Ta16
KmMr67WiBDtg9ZT4CIShB+MZnRROeEdHaI1yhFkm2teMUknZgWk/BTk11GoE60VDaepNipF/zHvR
p0jNODqTC29A7NYR+P5YIi0LoK8DuTxnm/XCviZFXBxn2TetTVAne8eCOj4GkATFzpuEccLvt4Vi
IbjIdIzMUSdzio4gaKFbNNYRkNQK99e1c6W6sjCymSBWiRIgHFUa29oUI9C6NwfU4Ia+hnbja46F
qovAdsCUweZr/+d5c1uvv8CHnVX2fDQHMiOb4417DBM0+5AjcT+XXG0kf22qPxxLHRNpa8OYLwjS
QwKDQqWgogT4NM9+fP7xWJy251HI5kXfkQ8+F30amBcG86q2Z54qKI/Fo0MPfwQEjfYffcaqEN6B
S6tzJt/rUnLZvZIy+jzJ9+pNUEDpvTkNLysHjDAHPiJp6/U1r0LTpTBSRI3MHcG9DuZUhSPxrl+j
1rwGWBRf0+tSp5BhRJ5+IPVUTtBJ7qnDAEw8TebT2lD8Q+lm2kXMpGyA7lZx+H+B/H6Th5cP6vk7
hiqnjqNQdBhvf+olzDjlWIQnD7Ve7YOBpAA0vpBa4DuuyEqmx1Bj3P6pyLd6I0vES1FmlOoMQlU9
4nmpvRKT58+BXeFsMrw25O7eDB2hIazDew+ZFvGarxXy6XYK4uDQWfKBnNBzoPv0yfg+Khp8HO0g
6ZZ9gEiUbaMF6VMyuGxLOtZF+ThW6xiys8LkAC4KVLCBoMRdEBu2L6BkbKykYRyUnEtflSuZS/uX
9hWUOg3c0yIp00DnK+qf3YJen+3aMcMeIArez2PBSm7ChfB7elfftvEtEr8OvN3MFtHnEgObBbuA
yWjCe70FdDBROuqhwNHM/sscMRDyIgXjjWl2C2c92jnitbODTbtGHMdnYjo5xEaGOWMeo7EGXKEJ
ktrxi7Ic1GOKVXYjLZYwqsiXSGjuQ2GjCUHMATbHskQlng/Mr+uk+YhaPIhffmRGXDN0pGZcRkhj
Dr+UmGqeZP0D5BY1qtVdQBemdkofqUEEW9F4N7ENzaSy+6ZnI8l+yK+pS5MIX2WPVL9ZNmfVRAzx
omvCQcsGZ//b4Gwknt5kfz1hifOPe8XQxYjV3wiETf9DGQlXbk8RfUktRu7/icvgpuoVDwCemFT5
8EudDdEw9DzTJH0sYrYluEo1MV8SYbq9Nd006ECDTiIXo0tvMWI3FH6tBmUkknw0aH5CwV0k/zgX
jWJcBK7jPXEz4e41RdFRV5iex3G3Jk0CLu6rOd6Imotgd+IGcDwrCbQZNX0Oo3krWZkT5Rorr9Ws
i/RjndVHUryNLDXqHxjBbkYsJDGARKGys5R8/sVWfIbu2dD9N4WEkgGCM5lp4/nC8z/DPhk/OYjv
k6ntoBmhSi3GaYeJPPQ+19Fh72HDzew1DbfvMVWDOawWxd57XGX94GP4sMFPMGOvEJ5kYX+F4Ca9
DOCZEmuxm3EXlDSeR2Sui3giWY2z5zIT9D7PvQpd3wol2fVemUxbMKj6fRAac8EsZP9udKJDMVKx
VYaVRrKD60vToSYhCJPRihz2HVID7jJWI2+SAraVbhfSyGaHz+4c2u8GgGcqV1CmdUY0mPl1W3oP
OVDIluB9U15fvU5BVKZdUuXyRJ7FjOGpJTPidZdPhziWpjcsKrPv4VFQ9FU+AM6QrzOdjAl2FDVq
X93n/kqoRajL+agbXdFM6VH38jw0nX3Ii9/fLm9SX2W9bEPktNzp6oMBum0VtFPKGGZoRubSt3UK
bBwxQH34iFfA4oHbkH9wDj/2hNPZIVyMmTqsrt1UlcKxyRTC6CrNrEraHcP6CuEfu5Bnf3YfyEUu
Dw40qW9bnKem9Hni0mfJ60CMgmb4ZxS6NINyuYy1RtJAzkPLQSlEL2Yb5NjBqoJ0SfK1L11kePXP
TangZ3ChgSiRLPp/1z+yghhnmHqPCQ1b4lOGNrvHSenYH5aYKSo9KPuQjHXy1B66L4gppUyUGfI8
gEdVOkXKcPGdeg6qN/lyTqQ4x/J9hoFB/jQgjhGbOs6lv7GaFB3aQZC62Ll9DIW89VSnDhdwSB17
Nbugv1bBBLZ9itr5P8gHZi73fC7Wgn0O40GxFt4DYMsL2GTD6dvbf/zu2p7/C8460MNw/OGjDJlV
lcptWqsME7Uv666nm90hfXP3z6rL+EI3EIrzPtFr4Fugf8eVkDdrurQVwfmNAlXDqUUSA1dD85YF
BN4b6K1crIcZUPnr4hM4nOZTlYuWCYV4S7VH4pMohOgfPUtR9BdRF2VIXkJhoZClK4OPr0evtzvS
YgH3Rql8y173DCMfYDaS/mHh66p/e6Z0IklPIhDmS7uAPNBUuTXLwUOeK+QZRwdfIPmon2kOKiLk
TNJKMpl2cCA8871oH3ahJlovD2oMjz3CZ7EjlGr7IWMrm2pbnoYWc9tZSO67cSGv1VU3ZcekE6Al
AjGaxy26XfoDuIbpW+Mba0St1jBWeBPi2DwpQ7VmBmY+9K4xUVvgx0Rlzv7waC9rZy/sXXchZo7O
GJ05A5oJQ/e/C9mWORR9G646n3/AswK8wONzL2/j03onoylyL67hzKsbdCreySeae302OTArWEZA
KyoSwIpLitgHj+g7aXZrZ9DAeS3oHSGcX+sflZE64iBWp5pQSrWAf3Z1GKTKgpXdDtJ8F8YkKjb5
045AyGod2ibDWBuk6ps23NisKVbpAVy39xxuJLW8dw6BrruKjN969u6SrC5sbNN/FXTyebN4/M4X
8eDIYqxn4DcewnXaSby+r7IjwhWbmhwGOJM4Q6ZtdV2cuBKUJd5Ou2jmgwp5AFTb4lsKNi88wcXO
tvOlwoQcwVHWsy+haf1tqZspmsNvAdlNUyyx/YSUhYb1thXeejL5kIXb8xkNhhH5gvzqfcfj/unp
UPysH6DuXSIjCpWCMnVwzZiil8Hrfba1yWs4KmhxxlJybDc5qfDEg3pEBtJMUIo8t2l9Aa7UbVRd
3HIhL3ZFxPTVqNCwWe3SQ3MRae+XfGkaglZuOnLapfFfXPHPCkoyZiJzKhpLvfwExOu+LwW3v2tg
8e59GoWmCyThP4/SJ0G6dGMzrScOAjsEw4WXFpskyDbEqyQ12/4OQcQGoZbCAD6sAGYZdiiKhx2I
6IjwAHbHj3l3TkFltiS9bN4wl2d/eHbTgY3CBnK1aQC4EBcTmP8brG9xoyWzXdyYr+Aj9o7UjeyZ
bDDKG88FH/PTtDao3QSRuRY61Fa4WlvpzHbkosYAoRwH978BTNwnLsnIm4faDBPfOsUgTGOYZ5+Q
/cpgmFFxNSt0aMRsTeUFM8ih/9cr5L0w1f1mwR8m8/ALurAGcVaex98ZV4GyJftPDL03kXGBJZ6A
ukvH/3Has80xKybFtJVBPQ7KSFN3YLE8jTetzjw4BG9i8GhfVNq6zzabOAfqQmf9irfnKHCy6s/z
Al8+/+hYw/WYSBJX6mJl9WRIbYCQJxHdD4oEuyWa5gfuSSNx04W5rwC+Z7NHqbH+Zo6vltENohEu
UNzslaH0HTyqLVQ4rfbqsR1rgaUerSSvWHR7ZCm2w76s4lbBZOjHDVdgUf/TGENFdxsBngGfYZ0R
0lu/f7YKazwpBH8ebFf1KW/3FMAMuFN8f35A7A3LtyBAuEUeJ2XbQQdXijdhkzsZER6oddqQ2C/P
6jRbHJ9rjl/wwFve/zPMFbxIUO32nk2pAvRojBCmLvcCzO645nZ6OtabmNDOkghd0Q3xu0QmkDgt
2VjDgW7XN9i9KPCmN8hzOQP1+r/gYQl1AzkVBfWx7Dks1gTW/Yey99VCq9UwlrqZNEwL63jrtiIK
Lvxii299mKGxbWh3pssUd5JlWrZ+v9MdOCs7niN+rg39u1tC/TvobePlczsmW4SuTzL18TuG43o3
wm+HWrwdW3pDjnSccDKjArqhUGgXBtFNi/kIwz3bR7c8eCPPYXn+3072RUyF1nSOu4N4u6BbNjAH
Cw45OmxyAvVAFfpPcuBYsIUBsQrwrr9DRUxLDhA4V2NJI4hF0d2BPpglezRnWFmGMiZFnZiYaLMY
umOHe/EWgmrX7aE1+pRVYLRDuGS2vcXy/jJQ/3Axs4WMBZpzLEYYYBzbcu5NWynackGxsF5c50u2
4SIPGbJUpjq7JF7guLClkB0VoeFywY37VMD2jz3CT2xGmwIUWiNaz9Fn7rEGy3h1bnAwM9JT7uST
3BjgjJAlnD6HT4v1+8SBQBo54Xm1WqlZkgoiWlWP4slYPF0vkQvVs03sGV2wMO25u9jrkZIK17MT
8wkAlnpSwFvrs66lIy4f0JmZNa8xQBGxC2Clm0FyeLjMEoigVEtCMvhELHoiG4zrse0rteGA7Pbl
Hc4wWnRaE0GQvE09omN9suobKZb2VOBzm0O+wNHOlg/nZFetO24++TyTiHGhghSUXshicfGb0kr8
D9oLNq/WcJfMWFwzgdZtVH/U5SwhFECpjpCwwoG+dN93xSa8R17Qwg9A6+TPqiEhI3jWglJ86WO8
w9geJaFpVTABnYjLjgKVnpPfzHVnobEIBw8GfRIYi/o7nyHfAGo+QEqhe+FozpcGle1RDhc5gevk
LqPuhss0E4jky4aLBhxyJq7jf/IAdYbb/XkoyGrZpiAK0AyuBXHMwGP6aHa8FETZJfrzIV9hG8sK
rwcJ4K1ryUH+bmBCwCa1iVxXAVObvRjGsOoC02AM94pQ6RDeHvdJSgVu2uKEn5Y69Ij8O/OrCc6U
tEmIovB7QU1WSg53t/Apnw1fwT/h0ebUAVBBz5EkGESN6jaE6Yy3qJHbX5bs/Aus3sqdM+GpDyRr
RKyh9KXR7ug0bhdKESNhCxoeGp4Hjtb3MrPUn4zj2HaGgtg8DENkEwMvaFTO8KeBuOyk1gKnRnt6
sS9mJYA9YmDa11/9Dik4B1gwPTmkcY2WxsCdB6BHgTtNASUajqWj3p8sfZlYZURBe9w81iH1W2cm
FGIhJk1SWHTLUtY+E6xtPWLx1pb/C+R8Eo/f89ZByn8JunbZKmTs48aOhaHJyyx8MX74ntjgW0ie
1dGkd3gQVRlWJTkRMg+NwdG2QSN5IZy9zCgq5M8nNf8SJnO+rY+9DTFM0FFKjk3Yyjnwcl28Eiy6
3aMWY1Ie0sqZRjUWTinrGF6tBviuoTu1OC3Ex/LiyXqo3Li6QyJHYB1DAeJSQiKx9uWQKD2iBHp0
ETQrt/qN5SFe9o5cHhnT3ZRn+Kxdt19q+B2neT3+iX+tkaCotIID1FfVCewRJlmdG2KBKgr9lJBo
8xCbYsMGs36YQf1W5MJ9eleNLTQG98X8+H6zvj4L76Z2eB7tp2i+7fXEIKpEwmrH9+Ogk5+kdcpY
IrzfdWhDv6UyrABWQo2HG5ZBixx1BzH0XW77yWEUIE/iXh4HzBKzIc/akLAvzTCzQmVdNHvEv23y
kdOev6b8Kn17r3XXWHezaIZyz1cs0Hn43BPZ8ptcMuCQ9U5bm1Z9VD1dEhbjzZSyqKvJHxe9b8qg
tFdcVXHdjQAcUA0E3pS5ebytDztRqTsDTQnjn1XA9TC5YyxzEfsSxXHZs4D28B/3iquYAmnTE0pI
mhsQnOE1+2IGrJ6Yf22jzY2lQlZS2TnIIO3b1HiEqjGl+OAER1onrhBapbzPvcZEmObTm9WbnxPY
RXsofXEYQX9Ies9F2FzSzc9BRRKH6OZYt+Ce9FjfcdR/UJiSIc99YuTN8M8Ebud7E0h9PrAa9/CV
S4oEkfDhnh5OIA+UFCN0v1crsNwPfMl6EbVvDodlcwpjV376Wn4hKJ3zeuw/fJkZYIEDVnXF6OhT
hiEWxxDrg+bDeMuBb/hENDzKqJ/EFh407R+9JT09r+NOL3wSjcb6FS0e9zTxRVV5c0Ia2jcjlsfK
m6yTdUKp/1NC3Ufi+Etza/ttlTKSwPETkS9zIgN02eRE7k/xKrGF1/DiUkTkfQc3vHdWjgiMk4vb
0MgtmSOId0v2rVLTD6+H9ZyX8CC7Wmiw+CQmOqQ6/Uf8pOaZoK4EXVhBrM9JKlJYsi6BDQNTiYqM
jNUjWPYIX0xKaNem0HlV2w2imf4f45ZMoyW3vDzI7S03tyyBM2c85rT/Y1Sk9vP/vHaYxLtyH3wy
IRnYAR+RrRCkR/2SPNC/CDWtuRz23J5vcMDf2m6pF0hlkgki6JyA/cXgy8pCdZUNtk0LXQ/CNWG7
6xlRUTV5lsLSfwWrSVxSfpEVeU4YvtJZWzVDFtS1lIJndoAy0Hu+rNSpoWV27DJfu1QOWpqXiFd4
h+DJU31iU3lppRkOLqQFKKUGeDfZLUUdOeY5eiLsSo59qR1aElMgArTVyFhvxyOY61Km7gPQY9P5
FZ6g1Gdsqpwb7DzwazlS1hIAjKIxi3Hcc8flNgbaITeAQclcRHqJtxps76UNfx6lCOQxwhENi8DI
msFXt4LANdd8Eke5TizqeDAGDvRSmYL7LJtUQsgdeUIyATVWGZmplyn+MTfuXyQtsLnK6ltEdIUw
b3IoiRGm+QA3NO9FUe96ELtoFhg00v3+2cAEYu5X/6KAFrU8AIPDdQfo+ewieh/mk3WJdepM868W
54bFCvS76U0Jix3wuzuhH9LzyJHJTVLbtzfbCht32k+veZdaFwAQd3MO+xuOUjkJ9i3+xwnPLFPG
I/VAkMMxuXTWLnQlMEINZwL8GNB7834YP7+NNmk+Dlyo/b3bGPDJTISp9n60kbTNaWcAWE5nIEme
Vh6VGGW4J7guO0qumzH2FCfPime+ZlOxai15TXrsrCQD6bLpv5E/R60ipCpDoTlc3ofYhND4RERQ
jRpLA4Y1TN4IVTwwi8hUWo5WUyA4wd4J4SKlwxvceJ9He4GeDaUpw5DaFU2S7oeo9ESGwrorNGIB
11Wub1hY/e2Ow3EjzX1F9JjOIk8K+x0CbTGaGco73KiFsYLQZ6rEDUlkfFbuUVDVXCd30na2BCdL
KaIQnkE50wfher8/aTGgnfOPpvZ9TrgQJO5yZSQIMMZU4HvB+sLwiFcx/5t2cuGDP/RvOHpPRuUw
qR81UBGMgAjARy/syaHFaGDgjA3PsXWk3sja4jBfJo20g38SmZYddWWv0X4bbWfwelH5yVJZ5eeA
+I/04oD85xLkzqGEdRX3QV/sBlVhMFR0RBtC+BTcixKuvYc35vpC7UH3qwqd2qMkJlRsfHE4YXXH
N1kN4Azlsu2oyKnuD0j4fahEK2SKiWbS9Udwn8NDploKgoxybiPPoYX5FXCzRbwTK2TIhplJztJ3
0O1Yh2g4roMdB1JgMKjUq6Gq+zBxEKmbnc0NpCnj0GbU0zQmXrYB9EYg+JWp6No/NzyITLX+rM/E
pyGMT2yqlPlOdqcAJDIKW9ebO0VPpGI9WLZIw790DRJIRMUhrdeeafz5TfcsbaF+7qA0FoamDVhh
V54smGZrpLDvjNqCHU7R9sVUcRIJhKdpFpVSpJUCLboJiwdp88Et5dlGR42gs+eFJKvBXB0kYXzo
1jwcsiW4rlBApWORC5kqKRYIc8/sIsltbeouH+xfH8jpsrFsFnVULN16X/9Y/TWnnUP1rfpia0cK
vDy58P/cvB/cbc+BGzjTa3VVm/0GadrQb7v8alFjOWQTeB9QlSiGIRCzjq+ofzBi9TXNLyfeY12t
dqOtTOuaYCmGqPnghsOMMb433an7Xo5VaGAcEQnPvDqPzDBIgnsiHzVW+kWDfU0dL9M3/UjlWdBs
IFYPilX+IfCbeFpLnft8javrb/ggbUHWeCzCL+hNhJHXGzEIxo+twDZG3C/yOrZJIvTvpwj72sTh
49P5yhGDNdZ5mEkFmda3cNtcPkeKwWlUcZ2JGy1tPZdnMfWl3HGf7WmT0g10s9/ZorZjrFE+I5pi
vpAV9ZUIUe5xlrBeP27lCypCGTYkoeqBG1lU1IeMICpJEW8Tz3m/Lrnl1kBAkry5v0SYi9Zdspph
4Sllv9x+6lzghKFECF64m9mBdcPOT3w5pUQnySVBNvMrvhvQldbDpBCFfpr6TORoe3XMsJtG8WeW
Nyu8P/EThRqzHJAzFYK7gEklTPm2UZmkC5+UznL7DTJhyhys/slTLB12U3rQKPG8F5YhgPQwZvwR
TcgA/Iod3qTDhBad3SgSFv8D11Q9XVLJKsuHdbh4HFj5Dldt5i/yA/IGAoy6j0Yi3Elxzt1ucRq+
1TRgtHjvgvr6Y5IZF0Z4JrUhteyk83FD1shQXc9khyS33Dv5KN3V4MSz7+LlMbofLABdzr9TQAXg
49H2ZzeI2oii8md+WFXSbkOAVhNTG9x9drcDB5RHKyzVrdh9gJwaHZSyNb/BtvdZSri9RHlzsRDQ
TTkBNzdad10+6ExctvstL/4RAsDHZSzLNMPwpCUqvrA2ugIfoFkbnHfjrEZDGNc+A6+O31m/Zmvo
aFHr/UfceO6uvXau4VG88hcXIy8NZi0Any4HnfxonYdY2ra5ZIXaNU8LsKXLmwo2gdZcrO1WYjCa
DJwgkIqxH4+fCcI9PGcetFMwFODF5IMliuOuAX5kE9JpwxD3F7KQ4wS6DCgw4bUd0NQVdwfq72ht
Sr2/MVuV1DX+97qQGZ5Wmek0Y4CvKa+IDLNt1bYSBOXdRGspQ318KUU5u/SaWyvOA3Vd8RCdYYz/
IZ+daJVPYo33GfQxrZEirs7EKhffahO4Yybqvt8Ye8vcoN4v+b6oqETO3ySMa12gvCkNx9PlYCoV
N/xpAdLnbELmhmlZWXHrMXWXO0frIEXZ7t4hprtMVNjcA+a5eXj5PPivn2074c+HhzG9WZUGXdD4
7KmrWTJoq+dPjbU+9cZMd4jFl1tCt4YPrCQ0pSVVA6ccxs85wCnWv59zYckJ3owDE2DTMgEBHuZ6
M/k1XkcTs5i2WsKbNnS2NdgCWGZTjjp4n3toS2y6PpCUZSbxsZLyd/z5qye+fjZm6pR3ipZDtEaM
sAIwImFShqUiDlzxjzHKZ3qisLj/+/4lli3qLChiYO5uYGyZg0sPTvhRi2ut4yaorqcjR4GDPOiv
+kAcH+5pTAdMOnxFgTKBbo5+6L/d0eu1IGmTOOTBLJYSkKy9amCFLpJIzzOZ6sm9bMm/gVPjA0X4
KB1WS47TclUsjloW3KoLTw8mO1uz9sE6XG6h7Zko9FAfjhqizfeRo6fy4+xfGZ9J7ntbUYE9g7c+
KIyXnFOstfltPHTTvU3dG0Cs08diuEnLzTccwHv2Ssss7EEBAhf92DsacmAIi9DU/Y8wfdvrD162
LJM6P4DcS4PG7xjJ5iUKWxC0lFYF14c5FI5Olu+ns5vZnunvADAvLdJ/UUiSL5XjyiOyqQC5MhWS
6XpGnv8N6iO8rssotnsdP8yuAFv8cqlcj1oFjaelKiC4WZRu6qjqkr0E04kWZCfQtm4Xg3FYkmuk
HhWD3uOwXBgKE6SVvdGQ/lHDrNyFvr8EVUJXvelVj0aKeykhFqpCN8tl8ZxHEF0wa+bqDKXNJkND
THPpfbRTKmmJ6CmHzg1jXzUQg3gVJ8QrH/sq1jK+Nfd1SkxoelYgEeLH8bQTmB0wAXfZK9ATzugQ
yEnezKcdLlC7Q9E81/UC5v9wUz8KyC1tUVYiqJDRIkt3oMzh8Yh7v0fK6ntRh/b7AkAml9YvdsB6
6X7xPD4vh0BJS2PlxQ5mqamdze9SL55WqMe2XwcnR1QDdga0O58l72SQArP+HPF3oGOl37tMZr43
BLnE6ncIFMvzfW6h6v5S3DcI4LgCjsOkDUCLFZsrbtyoRgjWxTh2z2ZIDOHrYg1LcXBjK9ojrYQL
o6Zr+xmb68ImfKvv2Sew8uZvkDjDoxU6GVyCQVW8bSxzxwIEQifcJEF8bwcB9UyfgJCLaIn4C8Lo
6ycGWMirwEO0x+5H7GgP2sGt6IEqinfohURjOUozrN3/RNYBDooE6KRHt187d1Q0klZxN48DdoGt
tqbssK2n6HlcNbvANfqVnzXzFNuXuoLNJcDMFIdpC0oH8im3iAcMWi2gd5JyOEjuapOlVMbUhQXV
0htYINC4yW+VRNzQ9snk1z/7QnxieBK9wcvxo1Tz83H0AW/xYyhGgDY2Z2cnUY99RgavXtQVPYbD
VAKMAmHdO7CYWKi+cmW1sN1f+JmMFtvuP+efqkfydwX5pV/XlFUf8KZz1m/TzcvBFnxO58ZYe1xU
7YAfjQvXL7uB6LR2Ples8ow/m6BDcWuVaz6pvWj6HTKhkKL5vjrctzeHbTuLrbhsFCB3t+ipko/e
TUhRU8N32ub0XTdrS8OqEP9s4mOVO4yj6s/BPT92qGGreTJaTzyrhvL6T29v/VikkZ+BasVZ/Z3N
t9mm7hJoCV9uuc4RSXPEeMNFdm1X75OdGfWbPpECjSvwZkU62pYTXdfbV0q8JSXXlTedwXz7sDn7
EDZeDDNIf7Bcuf/q+DZDyfOtU1VaLLdLF7EkciDkfYvM2pgvK+ihA/8QkjZDiUGktVzjqReiGpVa
0uzaS+T6yGJrJQgs1k7zfeILjWWmmDbDb/nDN1QYE3+JUkVOqTtycBzyljCOcwAO/Bj/vhCdFvsX
G9oWFtppkb9V57ZACi9kHQs1EVHVGHTIx0D+ps8Yw1ew1Az5zTajHzuFQkNrRFyzKzrFSyVXFl5t
CC3XeTHrxx2TxGM9iuNKLPa1+d//Zucj5RTC0wDkIQG8VLbJyI69nUU0p7EZyNbjEydgVTYQWmMh
R9aqYJ7kTETGzBkDoXe4TIbGT7DZ6V6hBZwJk665Cg9KvvvO12aXV9YiFpEwBkLetDWyPNJ6JZN9
YMU+/2YqYbke3OHqsc7yjSO9bvILLCsZQq2Gb9pGwmASmOl7Q7Oe+qntNmkjBcxrsWxzBgJ1GmoT
TpESXhwAjqV2fC3Ru6+BRS/YPEetgOL8UHi9tvzcMNWKfQbGiLNx31CgN9u1mGmiv7dRySqYLyNk
+n7+Rn79jTmoKGxNTyeu3mvTow0Za5Ivth78LD76sywF6mG+rZfKOGvsX5Sse5I8AcbErSIgWtVq
SNr/cniGkK0MO3DVoEacY74a0xHxB6Yfp7znZHVB7+e3Wlzt5T10lMd0OSYdqbwCA8nS2CBeXquS
ja2QNu5ZlNPWal9MQR72r0wUBv/lmMT0gdn2Xip2qwgc7FMVeP6RlpWSqcLKZVA7Q3EO66xo/MrW
zJj0/zyuMc67Jy0NkEXs+iPVPm0rNMganDlsBJhh808SJdmTlYJi9Vai2DOS2B6noh6M5RybuT7w
z+E4OXHAWVlYCCCvrO/9+StOiC4ztdlIB0AQLdao0XlXrsYH+Jcu4ulu80KjIkCv37WDcXA9hZKU
DbVstCw87UsOiJEZP5W4SO1ySTwTJ6wkL84TJojt6bKA7J8alshZRn7XQaNld5TM+wXXzRt38+Az
1eijFvCb6Ov49ifPV2C9BPXqd2SWakqPFJsdWKw+G3VuFMt1F4njLXFXzZDjJs40OjT+BmjCQyTP
PYj1QW5vmOvjoARINPIBoBpkImsauGZ/fjLtENpOzhs2VdTZchRHBPWswP3ERjLBdBdxxmKjeg46
3o1NPJGWBTysfKc1FFb2+S9SGaAjOv5OtRAyCDeOXDwd3y4I9pZAbgevGn5tYK7MjhuJcmp7IrXp
JLdZx85qDfYa9gh5MNtGxCxIFLsGfTwhiLuRScUlelfTOXZ52l8G3qLJQ/fTbtd3oTIXQu7Xtcn9
OwvP/5H8JHoeVyGp09jnXplNbklhsot6dX6/gBM5ud3NabQY8xAKQzJVegERDLdfzLsQBXIs1wKs
xBDFbgqQKJu07KQyAU7bgJ3GzJTKy+nv6byX3BpOr3toNoKgrRNAFWHBzHSBOqwJ/aIYwasB93uz
iQGjsKw/1/mc+aUethjj0L4YY9dOhWdpzFW+4KDRpbTRuWVadnTrMLOUCLsFvA0hayyDO4LF8tx3
PXkO56N0lFllbkZYvRg8HM4vyxi6iOFnAFyFoWoE9lrZjXEzzJnLVIojqOWOwD/f0wOzWpxis956
1Vvr82cHgDx0rjMhLdMlpCzp9fGnjgnrOLYzW8XlsYB2cKuZ6/ymqDnZk8ytmPs4qNGPz4yvspJo
bRlR0khkEo+6BySwLX3aH6uMunsC3uU2vHAKit7vMRsm9cn5lZBNvU5sDXe2zRALDcrlolfqeLFl
ocImRM/eOqAet2ZNd2ZQi1Des/TvF4LWFuuxhgxt3Ml04GQg9GpPO6fZriS6Ac6lcLdLfBwCgXg8
xME540E8ltoIHUfsgwYPU2L3FgsPntutyYHGMw3Rcp3X9E29UZfWdpogcIL/mO0vtznUJkdBze7A
qz4TJFd+KQFoSALdb7UgzUX9Ct88vwNMT2owPkDQYoiqO6iSS4emuEDDZFSSAPdy3vqoVcyQ7bwP
doMTIAV2q17vqe0fVjpDiMSKiQ3cZf7c4vPl+kAHLuDAcpbS8YLeSInykxMCZXnLvmXmr6a2kDts
WTAUkl4c6o8FTsV3Dok92R2vT1jrSoKP6JMAx/wDyN6A0UkMFtQR2ZJkHwUdikgiETSwIwCTMHzy
Wxw/uHnRu9QQRVfw4xNz+IkC5zgWqq23DOkpjKQs660M4nvoSa0wuGi06Az+bvYzpRsTYHZw4Lny
LNJP8BvBWE2PbNFc7JrrAPOYKJkfIw2vIBesnnIAnQl8jGu0XoEcRRilJcchtCZgLL6pEMSwDuHd
N9RznnbBmUkn/e1WoZbH5MzY5YXRa++XCuJSRW7NSftvFnuoyoX7hWnc+bu8PYtFATJjlIu7gUje
3VzNgvNAO8h00OYr63dBhfUWjrh0+O1cSYsFEhaLU6hfih+o0qtNsIJqzVaPLcl7qSJYvURUptT9
gYom+fI347ObAlswn5VkTq5Mb0XUgldFJo2LGAOmx+lr+QFkeY6P9ZjsDaACnsarIS18LIq7YKN0
RSt4oiB4eeOwqSiK9zDwwX1WjbS8WfkoVSPTHajwLbo8YjjgLL/8VjXaHzdGxyvBGgYY6vkQSxqK
qNAjGJyRJRKNV/vC8Zl1q/x2AAE/4diVo+bXFMhIkTgg4UrzlF2t+FqTnocsPAyKYa3C6gfagOuG
GHrmyHf3VKLYlaAuY1rcjafJoxjHhaySRUqX4UkaiXHZTtZl4X0YfsKmcwoSUxQkfVZOTX78PTMg
EU73lX2imKBCM24DxEtmzsM+vJGxPZVCBidc+GHr3Oar6Df3rLMdXxG+kvvbkjNhfa/Yh1nVgqyq
xNXt0MRnSrfIscN5jV8YkaTApGk5yKWev5JRkrRnBBwMqWm+t27N5laHt/2somOTmTVwlxKspqrv
Jz3XUX+iD3ds1mxhFALqrRnO91mKjRE2Kew3MHPdUgylE08kc7Om1W1xuFSm32EDSsRBB3Sn6yAJ
NnrkOsKnNE8urC03yHd7eOdJL1L2qqvDbfznjeOE8Woz/rDV3g2AvWWX4zQlPa02AgfzI0QZlknK
Qg+VAoKA7mvK6bv2HVdQf/+Mn3wiYSrphcBfRop6xehkv+OK6rqgVstram0Ac6NZ/A9NOBuuIsBi
lRLWEtH1IOkzUL5Fkm4YwnCbZVqI6oe30CRTUwDsNxu+I502X20XHoGdLAos1CENJca/tMVgAEbP
zOCo4OAA9b22om5hh3eN7D7LLLdDueWjcF+/o2ScQ6uwWA+O14u5dHvPbUzZkw37x0dTxX9atX14
UZZ8iLxYv1jnOMcJecZhod9SE5O+kAaLaylrmGvPDw3kAt2Z7QqYlo+6nh0Ss3pjI8N9Hv7E6dI4
/eEO4X5NhKbWTQGylsi5I8AFywraSQ5EbiK8j3mvdLdSaiJUXIHclKBWbtYqd7A5OtU4/ftv1GMm
IqLqtf3/yQUXqoGTjxlCk3ATyDH+cpcaXkUkATFvNphluO/aYlEtK0AhK2uIwUjc98Kfl9tAp4US
LW2HioO/mQ+clxLFXGxRqA7DSMNE8uH+t+uRVTEqD6pDpb7qE/aKO8ue91O2nhkNmyB71Oh77EUS
mAsJTKRJwHQuWu7nY9POI6t6sV350Rffoj/eZd+lDv8/ISWHmE3EB7BTN7LVKQYW+SXzj4NBewBa
tnZhXCAoFL2a9cfTjOpsdbfg8Fo2+sNU3+u4oO11sOT7xqvmOdowjB6La10NRU+ngwuI19epXjhR
SLCz5h4OIuWHZZ9wwgImyRTH2wLt0uUmKl87k+/a0Rxyjniqd4f1vZOmM91QWW04zKpT0lffUKdi
IwdJ8OFD4r/iJgh3sEaZAGf19K9kOGILIgLSIOYyxoqk9ILHg0ajfOHh5mu7ftleY0Hn2mXJehBT
14i6/zGCT5FtUaPkP8ne6dQN0cDTtxv7RTxYhcX+qIdVnLwSkLG/uXC0hklxoOr77ylV8OFGTYAS
nQsIN+VJIYU/3soPezlAXHspyzgBQZaMZZFLg+Gmn5ZyThj7odlpkY0mV44rsydZYpK/fNRI6CJw
xiVXvtvx1pEgenpYOLO3SQ3Kg8YUi4+ezxvHx95d7KlKzaKhW7OFEpoKnrRcTAiZVu1sRk+gYUhU
6QcM8aaCnxFJYcOgzr3Op/InG5jW+v0/wuPpGqu2eqRAAmLU8fLHnUWKbsglyxoyO659DGjuyCPn
1NxdV7WfM44UwztkDZ2T/Pew8oUvvdpA/8/GxpejHaYL9dLAH+qxH03rydvCvxspiDXGaZ0m1mJX
TtnLj90Wrj6a/FMkKkuSTAwh1SLP1R0zpWEvnF6f/JE919zQeSl26Q/3t5ZdpJMvmEK9iEvOw43m
HDxONjYpiFpzoaSdigOXSmyHhHpmx6awh+ADZMxatbJUu9ln+T16TLUkBlHSOVXnXIvUWwT/8hsI
9d/Ame0LSTXyAs8HN3b/0loVKfm3esgQWihuVG5DdWK8pNiIpsZNYNavWwvHRO+Ofq9dUiNqPr6T
LcO5M6zVWOlLEvqC1Wkn/TfdRFm21J+oHwlDmaOdUJyN3+kxmcJzff7HnyyR3WWm0Amd2XVSOmNK
En0W7U7qZhORC+3tRJOfw1i1uHSIraj4mwSOSnN6xhXE6E7DtRkDV0lydtA1CD0AHhMEZFjOY2fR
U5fRkjQNdsAckMbTGbBA19XI7p7fnL96kd+W07hYHQKaJIb7xfFcZkjQ+9PohVK+c2ACLonFV8GX
0XeSXBXSi48fBW7KgE9T6OZiSBs2u2xd62yKNK7d75pds5YL7Z3t8vF7WEDqx9zOTPhJ/yARmeOm
xeoEx9Acvz5YiOswphJzBnscGjSe6nntaNp049O5b7mNpiQfbFmmnHPU3av6VSdS1QF/IxF4Z9WQ
Ok5WTLKuTpngAxeCdcbwkmm+5GwexK6EGOD7S2fGfUO2Ci3CWNGboMdNgUZ0INKlqrHI1TeogOpB
Auk3YN37NwYI7zB19TC9FgE12dRuq38AlFpBFINl5Qtk5GXgfd9jprlOpJewLh0vPVVEY5eURmoL
7V6oqeT0BbGJA3mC1CqUVRtEjgMO5SWOGQzLzNh7t1aFzjlF5QSVqeL99QkdZoHciex4Cjtnw40v
zIDIVpHu9ppt3bTVUI6gebluTDozUfKuRznGPWLLOxqyqfxugmFT5Kif/Z5pZWpSf7lEGLxqGaT7
F/ykKdmQmcTGbbAE91MCn9BhN3D+H2RTLl+2L2AFtj21VIU175TGeY7P9Vn7Upa/TNqu5tU5KHQU
gOvFEIATdlxkr5pl72EfBtQpcWbdJ8XOrwRO8kfXuAjrWBGA38WJbyPxvGCJf6cS+ziEaPSHweum
JofVrhS+R/guuwVH2uoWh6bK3DSr2drfo3Tw1c4j9jgp0WJivzXRMgw571GUI2OGXfOEq3Wc2hiE
YOz/78wSxID+axMt6j3rKc/sL34fXp5OeUl3psw2HRUwEHaikACkCE+RUUB42TRIe2odK1oqu+u7
Zj0m6nwmwIHRipukjuu/c0EkmKOqC46bxzFvtznGMH0FmrKLHB4ZtXjhHSraAAfhtY9VpdzILEV3
0KV1fAO1Zz1P4WnngD0duGxF4aHekk47a9oWn3Qf5fuZdW+U+QZ5JqWy2EybFezsHRXbl2aH7UnB
2tQvszjk/OQgNZkRxjSmDeGvQTSKk6YDjs4xCAAL3EmvspaC1CwJgQZh7ZFKMWjDZ8GAwVD64OEF
KjxCfIjXIk7q1C62XTiGHhlOvbEXTCRHjC+GpAqpogfHKcdkges0coH5WqCI/f/diaABHGBUCChI
rZC3oQxfiIC0P3LmYx3wbSqoQ6BHH6Q1zyaxxGfr99b2yeRauLIkBGrB7BL1j+nfZ6bUMbPH3Yo4
ze824ddMZZ5huoiBADIEnJxS2bA7O0mEPi/LCdlSn3FTgRvaxI6VaJcKVLtmnE95dVUHEfvC+8E6
dv1QmXcfkn1z4RI2DZH9ZbpOf9XkBpG1rDSFja/i7HS8dVisuAs1x9Am1nSyOHIqJQfRTOG70ud1
HRs7HD8EgsEncM/EU7JDulVYFxaK/ew5QwITqGx90yBc0ik0f7ybTMl2KxjscLIouMg+fgNCzGA3
uNv4Ie8xTIk9goCuj+fojTg8nnQxtglm90vT9+YeyGKbEij/kjUhtUPfGYPKCbsQAObzQVQpR+i7
lJhne3UUaA7tqp/w32xVxpl3ljdGUBd+ZoV60b+ydnAxsVhp3gpxMBuabtM6PfhtpbKDEUU8vRHf
yFE0BKq7Bs8y7+9Qptil10eBV5jsouVMQuIh893nLlSYr/Tu3QKL4vnNvp903ovWd28Y9ouhENFJ
0W1ZDRRXzCDHSnq1OJl+iXRGtFrtKetSkGjgP2IuJGU+g5f6zRQBAsLyjN+lfsxAmc5vpoz7rOM4
lztk4L6nGxfkr4Bvpr3IFV5YIE7EZIFzn2K8xc74x6c3wsam9brPYCH64Dydms1HINKJ6Y033yUG
/epA+VuTVavlvNUE+0atoX0DV9sWW4dHOqZXAqyI1iCK3QndVVpdM0aBroiNWaKBLFDJ4ayLubfY
rbKRPhMQZBZ02c3quHIktD46cCoVtWZFyV+ZASKbadrNuQB6MzMUKFvc2W8fgsZBarlykKstLAlK
siNDd50Akj7TOcZZl7NyCJP3qt76pQIXgJsf1FNV0tcpkxc7s6mJ2cDlKSmjCbEUqxHmTJXih0Ti
zOAS2gHYVjepDnIYVOM1fgUO9AhjsEQ/Oo3djHq2cUhHppgb2n9oJD2c66KNY7W00U73oPTuWY/u
JJ9fjyhyD+8P2CllZs1Z7Kyac84FXemqMDxpPYEg+zLj8j3yz7iSwJMG2SNNTurCITsypFiA+ZDb
S6qm58Hp6z7G+JoiIEaCFCyKWOHVr0A3KJto/pBLBgtnr/jQqHwoUhW05V5B2ANvUr1zwYiVW4mS
sbL2sL7/sSOfSyxpkjzqXW+fOdqsaHRPrzTfToXMdxR/W65pcSpEXwC7MiEHi9naFYSuBmvPAD1Z
e7C9hgHuSssnmfyDT/5jsP0hOIVvLzeE2mNepDv4rrgEntNpmbFnR2G9LW0jptjl4FXAt8Ud+9ff
Vztzs8phD+Xwj6F58w7vQ/nj1mOQlxMimkn+w5drPRjTQUb16duVynhWUWALOPDz+edVZyLKDAYV
eoiQRYrtqhjgfb3Z880H+dyt8K3ijdIDdNlPViXAY3sZf8pl1wHco5a8AJwMk1tL1pncGLhSeZhU
njwJKQscsRN7n0I6nmqvbwzXkbzYCj98Es7Hl5zxz8oi7tjfOWFZWP88lDV34XmOPvpseMCWsrkE
m3ppiK1GWRm6Y7fsEg67i2cPydaEeSiMz86jxKjAG2SCKamP8Fjol+dnY/M0eJ4kqimdCa18QseP
K3J7THgrIKkGbyptcr/3VoDmsXrsvYANldFwjKDGI2w6Id0Y5F6gWR/OgSKQB/0WyKDePEpCHiIQ
Sk/r0EbjwvlrjnaJoJMiPSN9lhALKg/qtshEvDFKYCoJaxiIpFD2uY1438xb5K6CjCLr9wGCR78L
Z9rpBF3f52TeO1QtH1YIJY7CP46OMhb0owa31ffXSo3nS1Tx8OG1kSrp4rhYRp6HprpE26/APgHR
KdAOTAhLQhAlQHR4VMwMClnHtlKHqMGXqCglhMZuL7xisYAU4YqDTA7bArgc98xqS1wfqMWX9yjy
4OTN39yUaPiNG+TJ586SO6jsrVwWOnSGpPkJRB0/6YVH1WY2FjziGAZ6gfuItmEsMVcbCqZT/+z7
iCzggLcYcvg3RPBhddqi459sYA08Pok7r9EjMgmcViPXrw/wv1kks5+SQ2Z8xtpaqVNKz9YWpsEy
0upr0bOwXHR8L1CEq2lDVtM4VFwlWYTEK3gmSw0D46W3A16HPUmU81f1X1BvPyd1SGYxw20Ug9KR
WHFLaINEp1MxuOLYXxF/+/jiQVtsNCh32xzzvSAMlF5kqLX5/Jz+a57cpxVa1kuwu3R2pOnEfCue
7XGsUiSuJCFxbS2mOr5lNwDGcoF1BDfnGyHVgDcR+fcc2KrhonchCizR0PSk9gVFraMbgMbiOYoq
ZDYYKwJiyprvNRzfpVoiEWXbVFrmI6++Exii6SebR39z0vJLSVvk5ClitvAqZKSdWoPI13bgzSZ+
rp1atfsrWJ6SSITLHXmWlQ5mdNSPZhFB/51qiz7kwATiR9LTeSsfCFwQtM57nlo3ABCh29CzfuWB
L5O9yqSyrccJ0BIA7p53Vs2/tjMS4aCLrn/TAdrmmxFeZEuJhWqlztlS2Cnd6QZxnItn4K/YSq/I
w0PiBzfFx4TqoulWUSJYwM6fVCfeOn7pa2kBNaiso0ubPLUAzrFmNvoLmXAMVzXZik4/TJFbsCrp
wljSc2WflxZk+a6u3mg5UcgCKiA61B48/j8LmuhixgRBsK7+W/L9tS/qqXL4qnln7OZD+pOM+Io0
hXw58/TTS+R8N8NA4uRKh+Z5jTQxdTaGWuQTeyY2JU9Y736GPLM4gXzea2cONaob1R1OlsSTZX85
RVMeijsuIRLFBEuHgGgr4UM40f6E1LEqHKh23JwfTre8wjvWuWBe4zE1l3cXbprCJyoIw/tZwzJP
pGb4TUq+uAW73MGSCmuorrrZBabiqBmWurSYzWjHACZfCeMw3+2p0XQXm6Hz/I7eSkvazymFm4R5
3ftH/SLIrYDyHnl3gj0irPpSArJJVVbUNzu2xD1tx8wdZuSe1hbjWCuxd8D5U8clr9b0j3Co8LYG
D/R5FigpkgooaPqFqqVIfmDVtFXk8gp56II/4v5sZSz0nstIvLgI1Tp7I0yFoI6h76MFfL4VNw4b
fcogF9dsDnsPGPFsp7YJFVlRF/PRqK4VKLPg+XT3J3zXLxwp3ADZT40/WlgK9fuhdF+GsfEEtuc7
Xahikf4uUS6U2Exx2Ke328D/rXdGe1nPgyhbXIqXItBV8R+IysF/8EXaaY4v0BTfhytT8uZcQ3Dy
Q/5ZxahT6Aq+fU5JHq5XP51HCu6exahavKU4fzgB36gk//eu7+8rccNRQXYtcjnEx3Ycx1iqS2l/
B1YlsMvgnqiNjKhXXKCNU8kYrzKnk9EbeQ1K+AshIpnZoSBC1ef1bYNn1vgzEO/5ZTo8ZS9CELZS
8jhZwU/FPNJmbso25oKtycpsRhzKzTPNKpdJQeGZ/P6uXiWKJXJG0skWYLeupMIlh5qfHlVZUik4
TwFVU/zQ2ZVwSPE1QIWlMpVUsPwO2S8krD/i05UYaDkRfTVt9Pj8ISctPEcRJqxC6zApqBuuCf7/
G2+oTMaL1CysEOyIVWC/z3kUc1Ykccjevs/GcNH1ouUEPPt7WD56ij/Lui/S4WLovQVjnS3j+qBc
KMPZ8qQwiolEdyTuWBYEAT+Jf/Pv5HF33q5k9yE6AqANHrn6h0KH0ZavEIOYZlvq+7hsnxbCQPOh
kNMBI5EQtRBjSaqc94G615iJV2O1KK4+TyQczv7GwF4YMq+EwVaXDwqfk2f9vW3NoYhiuq8LrPZu
aRFw2/6fyOELvskf/YFYurpHTpf8crd4HScpk/44bTeWJ5KjcsBT2fjyLlROJshJqHle0yMuWOZT
WfMqw4q2BkBenQCg+xnDqOHl0kkR1ldktfZVa66WC9KSfe+89E3iwMBchWUOAC6NROXEItCAfbBI
0E1ZtBxZ3xkQpshU68WnA2bFO4BVGUJ++F9HJerq8GIkhlHaMZ6oWnrBI+de5R8Q2jOD2N0smj8B
u4hVxFacWmZsn3JhM4hUfsI9WN1s2SdNzPVu80N3uPyJ9YM9rBUtrR6zxcg8D8qng1tcj2fCOOd7
7boj7DOb5dkzICN5tTa+MUFLMs7HREZA7Q/OFVPEUUy69zqJECE+twlh0HmZlYu0V6V6hZc2+QGW
yG/vAdcyPt+AEhfTKB4O9CcRJPjK62ttNeZIzO0MrRBfl4USrpr/1vAavAOLtIDluKrF/ZS+i5o7
D5ftvVWvE8o2s5uZuzGkz/+22QSiUmZUZ34arIv2XxrjQozzml5ZQPsaDLuii7x7JRS+Sd27Mcr1
Wz+6soae8G0HRd9wvxF51s801R7cAm+1OxYZAI8C/etNfkj4XB/Ndbx9tjqX1WUT0YxYzxzFM3WZ
K1+OfDbe9Fba24ELgdft35Jeoy+HLQ7qsjvPZybz8Bcf7yn+aSVnk4+lwfiNV7f9qjLKSijVEMKO
wHTfdj4thDXfVEA9X92NonpMqlvif3PG6nXn/IgQ1V7ve30lRkLs74i3oq2mt+qsbiFZjaJtYDR7
uwuxIOyH/wkTjeDtyk97Z7eeV9r9rHMzjMoPc6QFp9N1WdI1r3hwPUNVyA3wJZ8czto3NPbObH1P
XjM13yW5+3cbhW/qHTFI2Q9UYgOVcgEq8VIEpibxCm8txJN8YQIEXWr6FbdUK/wSrVASKmfV+jCz
2SQToXDct/x/DxZOYpnZdjf5hW/iUFMRSTDcrEbsAuLjiZMmLO0brnLyuHhRDCFOnvI2jsyYHPZm
uFgSDQITk/zsIwv6r6W7H1Oy0vIwQh+AvLxQgCWZmYzypmy8tSkJ+EPJctHqMeuC6BeKiBscb2Q7
lpsb+JiKQXMnwZneEV8nAuMDAgswq0BgbzmEj/ERSYexs9PN1fIC9jlcdDbJpVf6TvmyHnp9uLSJ
OyzLXbV2lfnMvN+MgGikd43txfviM+SQts3M3QnRP1xe3nAPNPWR4S5zJlfjuzQy8elYP/ZYlskR
N6Gn1XICS09t+4QBUkTE0CDGJbPvuk4i0vCS+eE1C6fWwxJaA/U41UsqGyGhXy+P5OmcRFcukJuV
iiPOXek7iNd1Vv2F+PXBeEsgzwbzADFTSpkRwtLJgZJ42QC+ZgSWZCxXRHFxsnArKBjRPFq/LIVK
3qfZAx1SBgeOJp+JcNlRu+9SVKAqc+OFJH28kzG4n9laCZn2zbRxu7+qPC4UEL66dGilPQ5jBMxb
WnRMYpdGB+LfTk1cjn3eEcP0HNYNscIVyDC+q73mPU/jtdVhVisDxWBLTpOYBsoI8+SqzR1ruHBL
WrngtR6rGJzavRPGgDRQmsYTFlNQt3W3Ojkf4Zig24u1pEoGCGJzjK5dcmsTtUCiNcY2rEPpDUdl
ik85DhS43RebE4KC25Z7wzYZ0LzAIyMpV6PDzmAhVFNsOrLdMYtXVSHz8jx1bMXl7pZYJC3Rq9Sp
IQCFfF6bo8UCxa7WdHapxLIDCefIScVGr/AaAeGcgfauJUr4yBP4+7nz0gkHUzmOKM5tbuz8WRj7
DuicSBIqDxA4/VGQ0jVDUup2ZNvZZclxlWvMqWS8RITDgoaj77rUAZAh3ObM2scVMot9n5I1LvJP
7PStCkqtanYkF5ZNT5ybmODXuXMYeohlIQXH8j0GFp5VQHkt01LPkpHmWaK34AiTxGrhfaSSfIRk
kOWGeRhEiM1QIG/c7GX84ispsIhnBrDhRrJWfPDm+27arFwkXh7S81j0qik9PloKRSgXPKPJreR+
OMEGXjX97Gjn0anhksMT2bOsYeS4cygGmJ6bhJKVFX1MFNTnNTteXNGsFhu3/U00faDXkEbi7zhO
juvAaREDa10HJzPv8tQC8ArxyEF1sNYzq7Xl9nuiuu6xgpTH26TePsPKARZrIaqWJeP2Cj7/j1/I
oYUBE/tVKHp7y0cOXaUTas8wqoyPuVSA51VcTLND/C1Zo5gUm8HCg2aGp3BvOpcLEINnPfZsFcqU
Mcfmntm+hmo82Gpa+TFt9RLFtTEV+fBbsQ0BK7GzAKO89oemYHS7S3e6G9K6L+ArvgzeqD/ct27R
rqLFixUjC/5IYL/HwoyJd2S9UkbM0Rf4CmS/ofNBHpV+KDZh9CQ/XNQCPqU8ajiRvcV8QfG09jfa
XWKy7c73CTDjUaEVWhO3bP3vqDrIeQEzMTmZ0+4y6+/RFna74MZrPwgwEVBODj18w8yCL3xPw1Q3
VWHDox9zR5/Voz1aVVYXcPmo69BFOVe/dsdSBU8Y5wONx13EfrgzvzmawF9KBy4BQgMhHDWqWf6D
OlnDjEFOOl3WeCjCu2m6G4WFxlRjMYAIP5t5gnc3qq3QITA4U1AdN0cz6PycLLIoYHWo6sDH28jk
GolZl4npiMd0byKzQYPBEiQCn71xTpbv5tXzS26REmNCHeezh7v1I1a0GHJ1MNR5CTps340u8gY8
vL7l8uchDqC9p54fTt3V5/we3MlJwMQsiAXXkri3p7mtmQ2JEMI+R5HGbcJEDpIGSCyqRmiX68Iy
e18aF+iKfiX2Hz3dzb0FuCgkjuU/Z5f8LSdt9l7Xfvvls/3Jr3H/Pt0GiLWxvXdG05BPYfaAn6ER
Chjy87oduXVlX6NQ6eKoNTPoC2t9XiwoEYjETl06qn9EmLEtl1f5FcDu56cqvNmZHxZ02idmQS5D
QkdQqIBEmZbDVB7iDPbbJzyfsMOQMoIfPMd7d7QNNe4Cln+GpWxTUng+FJCTO8ithxgAzfNXfhrX
UTESeppGzGCiFMvM98ed+rpNXxbyOQa+RbyyxI07LFO+3vnUb43rQDfqzKaAyA0LYofe9jOrpFVY
WJKlMupewLzR8uJbxuky9EmocHPIM141HfnskFSfhv3NQ1535X0MyvJJx9QadDovi2zdZ+9CiwXe
elVQgzXMrVTqqfGicoDsrUkBu4c+NTcq5pVYvdQGNIaIIZAcE0fQjCd6hg+7P5FThR2TQeukuJfQ
B3xaRvREy+QWiuVPWU5j7UuOhO9SaDCJX0rzT5uiSAbGrRDXVpyQ/h9dA6PyNJs2c/yfIG0aHOVm
Au0yHm2h60o3rv9ef7DNbZDdo/MxGU9UHNHKkJRYbuyZ7RHYgy5QgWTALHMTJZBhjOuLSpUmcVWd
ZvQoi8GX4nwV+/Pykj2vI9a+I/oZfE+IS+TRZvgnud0TVXmaeYL8DqfoWjbbIa672vqI5K9LPurk
ywi1szONHvd/4q0yUzNlyIEh9LQ7PRpfuJNtlVnrsZLdtne4wdpNbGFXBcrk5xGpSpdjt0JIh2ES
h/dfSzCQwm50ayqZCbbhuSqsGlmJEeBGvdol6roi6JUHb18NHn1prC8FH04rUpE2pErZHZBk/tIS
hBsWyrI43Y9cyTB+c1KxTINj5VEBNLJ84Q+/f4dQ10C2/A0fs8Umid2NSkj7L0uqPeJNsta/G1S9
C0gCpAU7+j0FtAATpgmiumUBPwQgib+XavyYXUykjWIv8TMCTPIuETBM6M6oLFy8fJtODHUIhpO7
aaRDeQFJ6NPEUNRHqEk8VIVJpOn/IsUKHql+UZMLAqmtA5uVhVgoDENUvdDcWT7+TasgRtHULUk2
WCnnVdgOimD+mmP59yjfritWPbEx2WjHHeave9BxEL3GmAOBjrzcs/Stg6uTRjf/3qaGA8kGwPcD
OQfunQp2SrdaRP6o7seHQwWTUgv9zl0uKDmBiwEcMb1ebAGjkbzuVs+AD9zXrKLeMNgPol87H6DV
nKnUuRbR/w2+kQX2YaaM/5GMNnFEzgg8ovlza0Qmg6jiqFCRMh6JIBUDIB+c6aoPg4rwqSSgLt69
DwNlb0oirDwCViF+ELnXqVBepfnjjXwCezXWcbwIkuAophLfV5iMZsiC9+4w1UtaOUrPa0SuGvp8
jHJ1Eh2XxETqz3RcJcQnZx8MFM2GzfNGuxSDVYuZdUcWqnBKMHf5FfsMx6ztz8t9JHCF4UE/r/ww
9p2fpu8hR7jwcxJgXqr99H+cIRlt0L47QZcrGLXVljxwuYJ2xaKNtWnkli8Yc3DWDT8k5Pfqo+f2
aAgn4v0XhMi3PlyZPHGdVdHAcSLd7EzE6rKNOlzZ+s763N7OmFO+CRE3LWQviQk01jCXhhr4LX4J
pTnmnV5trBsRwBlRJlmgMD2hJOOOxmVai9vf/QQxunw0Ern2vCQBM/KPltLTvQCtTSd0udt7h0WQ
o6Z4j6nmLy3H0tAKaL/KJuT1EIVeaGf7CkyK55qMw60Taw2DL2Stw8VOWjQgLo4hoz96waVKtIIV
mNCLrYUHvMDE2iHaXrUmMbez2rKvgd01k9lw+uVVZmI6l0tkcu04s1pL4LEAMIWnuwM0Bi3RREbX
k216t7eVJSCWPSv+DnN8/DMcbBP9d4uT9DCV4xWcW4NJ1LSFMvZy1U0wyN1XsmUZ+QpFc4DwYDi+
4bkEaE7vtvS+tY3cjAjvFhpAzm/tQdSORDql7ISn2+zPlhNu+b4EfdDkciLqbEVPJQNtVu53udmC
UXuSZNM3SmSrVVPEzBXRwqZ3ScD0XDmVtYKYk8qYaZliG971xhhC/UKsKFaHym3zgiCwtCSLgGXL
H+412LZPy+cJ0VMspLog14CGMZ+4g9rG8s4Z/80C3xtyJ4fGjPZUVn+1nHE3xTtqJKItT9NcWa/g
DKOhtGpmL1wMzLFhAft75cqXGB7braERppcZ0Pnyz+lshJJHBltb4mGGL+Nh5TrWUQII7MBgUzxH
m5kF6uQUCwCdRk6aCWzS/Gtb4i9g0lNJWbbIeLQ9yN2P8N+j4OwXtbqjQqOzywOcnFgbN8EHuzvY
FlY5UUTLftetxYkL1Kn6umMW/ttjQeyNjKrOPvVf19vY8ilWlzivUb7d2BtlHy090TxkvBwvtdwb
pEbCUCNU3O/ccwmQQNTDs3M0E7h6E6ZvdQvqZANceMJ4xxsddU71lXF4nRvDLSvrIILEVINoT6Wc
T88epiuuIxIQ6VcXIBd+X331RcBqX6kUQlm47B7CAbwIAc+rJJu5gY5bzcYm1R4D9QG8Gxply3Uj
bZ2e9IB2bXsYOVE0WrmfD8ShqT60R9YLOU3lf11e6c974HEWO4JkX9Z1rT2IHg64z2IKPoNbur7O
guC7cm1pdBgFdpuGaV22v3yGcNjwvxXqKeUlj1To0nudc1EKfyKrJCCEnYvS7+kCtPHBhg3/GjjG
cOfmrR7WvZWdQxQhyHV1DkapyQBL4XzAf6DoQ3P2oA5q+xQQiTl3+7CzxzHyi1QdYR1RbBpPeu6K
5DtHmVML+MBCDoQ9HQ60xC7dBfctPUzFak1lM2eodElrmxRyKyRFon5TYCDprR0+ui3WjDjMldct
mx/YA3RdDRWnhnq8OWahZK6POMe7W/xl45Vye9pBfnV1eA3+2Q5VFUt9KWrrtmjQ5D1TO+Q+C8gJ
7mRiLuzYwydhSn84gItopr9/fX/TJQA+YRl6M7kV734dYDzTelsnV1i1bPnW2VaY0fE55NhNdZCE
zKFV3gJ4Vd/yFs3p7zcA8tLzOPuqhTtwQY1Pw4XzgnAqKDYnfLJofTOJYhbsr83rvs5lnZ3XrRBL
zruFODES6BFcx9wrgTRhyZMkoYsWGXn3qzf6VvIYuhYk6gqmDZ5dC9Er5hJcBFymUDsyw/8h6rN+
iLNCgYKgMGC0iNumdpSY8qfFreXrTdsyZ7dLKQC5BnkI77B6oYRFDmDtcyPgZo26wSdmrRDU7wu7
PShUO1y47iDbSAaQzb56x+dCUmJJEeFYQViWzXfDiuQcW3Qv834WVu5vDLLNoVzRJe3wfbJRvHk8
gTpOwDK4es/0tyWW2SlmwjHtax08YprPzexk6FqTbyg0bu0Ld6qGBWnzr1tuXn0ODplL+qGpponh
3b9mgZKnN3YCEE7lgE2/LbKGkPF+7DKq8Hzkpqk9snGFg9kLRIreLHF4OB0VlLG3ujgUzKC9c824
L2Fp8hi789MFGqs2JwhSa55cnUl4B5Z6xMks2ihEHc6GzwtKAldReXz7DASCI41fCR7foXteDOn0
XouogtwNAPwvCbXpNe9BLCxq/hKyFsFDgbwwUEMxU/LQKEqhUIVVxQWSPcQJki9n3y4qjQdBSyJr
pDxfG1rzeW/9Ul39QHWSljssCCQFQCyUg39flbGvtDmC3e4qzmdhMhtpMFFsBrZkbaKjgDolFs2C
qXNAYcO2x9k9ABRdaeLjmqqaOcPDtams/p2dnPAYaUuYAQgrjfOV0ZAseJdY42U8gg1Sh4BW6C6n
/KiRTSi4sgAEs9Tqp5TavV9PNtCZGKDg3v2it1tI2xycbiEBx1PR30Nk1AGOYSAJKZH9Rerte5hq
W4gPR+z/sBStfhb0ParQ3wxPcictWfgWB3GL8IN8ZAFnXbl1bBofw1QVPRAEW/mGbL25v5wFUv9p
iml/JCquQQSWuSm17U5idUDHOKOME8wX7kqZqgD2WFLV8fHzsx3J9eofxbhHYqwX/YuAfcILJiKx
ukHUTv/lrYkIJvMecYYamZ/GRaILlXrNnoQWQExvdFAaEYNYgEsp2gWJibSkaYRp5/kofW/FOoaX
oUR6KiQm8Vls0WudiUJe0bRlO5mF+SDYIvfuz7D4Vid54u0lpDmjK+oeKNZqfhVSTYAh4WEMI5pz
/mr/urKmzzauNRtdLN/57M1itvsfdOhxlm174ZZ+gSWr2wAi7eYsxnvCIrKrPkhtFyz+JBtHAyIQ
w73KePAUIvBGuy0StXMrnOMdeoCnIpaCu5sA70JnpCA1wudPCMFq98M1DeoZs3V3Qkdh6bWuaB0i
pjHF47aomoCSjThE5yPlWhOdf14eZrw8XPnczXS0YSsTOi/QSN3g5M4xg6aHVBQh6f3+9/h1MjCt
ihsKINJ58dqeUWYD+qe7RQvnyq3KIJlrNMJN6pN/oUexYbVCWxWz3TozWWLM/qI+eedpcMfy6BDQ
gnawANNK2DCQ7sQ4jZoqcCYLRl4B/GS8u5DIDPsSiVUmrdoXvt5Yn2vT/ozWt8RZX6RG9OV2DnKR
3FrWY/9yXgiYZxit0tI+7A1Tj2+/BCA7vr7du6xaHVJ+tWUfFvXaX6JsHJsS+mcUCAjc/VZqqJks
9jY5j7HKkxMNcCbMhapGpCdn/WzLzyxyA/6KaMxdfb+tPwel1+C3BqvNbC08L+hCzGaysKGao39B
/o6t1QI+NfAvA6zu4RnkGfkR/kD0PfEkm18Ct1bv/D0BwVGCqVQ4FWrdd62XlLdqdGHp6ruxZH+8
6/3K2sKcTFHx/oV4xftOvB8tVhqsU8UcowU63hdP4zfJ3nBEYnLMqxzcLAoaqchcc4V+0mMgL9Bi
fXn5EEKB4pM3GmdhxmdUttbZIgzHwnmG/gjUO4Jh2Gjd+LJorQ3lfxnHazqZPa48zEslXgSq5rTG
r0lHYKLbytDWBfRWZsSyrRh0iOXJkSKCYJKyxO4JCbLUvn9XzCt5Ges9s1bafKBUFBsdWjVkcnRp
L3Own/HyVKVS2beSPMV/o2ZFinUSTXhy1eTRhbKiPwQcdRvjISVF4P37bfQ6cItRrIr8RR85Uvqh
6ZpJFa5T/AhUYd7WqCp/v0zm6XPgTfECUibu/siMERLGM6r8C8PVKpwmkrLLyGO+nqZyMKFHYn3r
NvhZkI/99ejRbu0WRoKltZ/V+beqRSOvXYxdX4UX4tv6E/nrOkdac12vOnrI+JHzsUkbCCby/uX3
1Dw+VEAz43pjHPjV23Ck4wt2tRXs7rf1bMXvtcNYFMCkMkG29k3CB3TsDX1h7cM164sTonvZjxp4
7Y8gya0S4lRr6TrvG9C6CNAerS6JSEStngWJk7YlYTQi/r6XDTRVpfX4Bqsz9nsrppofYj1ht+1v
9JGSNBF9kt7J1dIbrVSRyDkxlQWxciKq+y87dSSqzpPYF+34EEYnsMMGPn8ViiMu/5piyVgXi5n3
7bE6O+H3yOUHn4cmvfTFXSHhCZRTWhjDqVbOYnSUBA7iU+dNiTu6dNVQqsB8VZwh8/F13fToXvj8
VmmU2VZnCuTkEiSsneDaPeTX2SUJA3SlpyNoSTo7YkPO0HjQdA5xZtvdJ+AzzId/YHy+wYnlXw69
uE7X4Oax5r1/In52C5cHNshTb1OIvwFf8FKKsjW/WEa1b188rgNMW30jxrSuFZ8EKWzrtA40EtvW
/fpRPGBkBZpzjdy3SGixMyoBfgnCh4RTRKKf0qahpSkGryyYtmbIFe9TDwSwfaY2m5WzmjfBN/L4
VWTm2qoyL/Rz90kn2W7YlanNTkMGv2i7S+8SMb5WHN0+e78bFkb6KOcHQN2bpdv9UPPYCBTXhjrR
Er3WvWWgxJViqksgyWvsETqSuxygTj7tQlC3nU+EqY31oXmwK79Vi6PAySN6WCUqXOJLTpFagr/j
n1jmkuJmn7B1zcLy8xrX/xMRZqYqDS4XJ3GUF5sSJWL0U4l9Q/L/SYXmJ89BdcmRyxsx0uBhtfi0
tS6S0H3h5AF1dpbflViW6BAw5p+TupomauYaJ5zPmjtsdXLglYLJ/zUznSXI8AB3D3BHTi33NiSf
27qVNgvgg4gc0vsRo4OJ4ScDViLn8G6N8jVR9rytmdud/E31RAJrXGPsCJ9Q0DalqYxtubVWxYv8
htu8JUYXeRHfdJ1wTVx4rlR7yAA6LNahHPpCHlz1Y/kTgEJjrKGmq8Q3N41upIsLQKyIs/h0Q/i6
3O7dhVUGjfw9uKX9uV71V2rHrb5n8hcesy/QKcT9m1mUiAu2n1byLlCRvEqWFUNG4NPRfRGQPLtb
I4SnsgH5GSCTZ36ORygcJgJm77nMusxAZrNiV74CDMrtRISkfCEprkn7Xe6k6FtJY3FTjWJ4eVBs
/ZHvg4tr2IanyErtnuNLMZX80CH+29MDHIF05CcG7pmqjz+Q5QBoJIQvWzs4fHpZWfPw7KfS4ye7
CRXYl0XjFRYAkujv60e9k5lf6u5DeMqw2cY+cx5FXp9Hrid3nxcJr6YCMYzZNF83DZS2+1fnvd88
LyfB6hHeK1pyJDZVBabFe5rbSfciqabN+qPQu/irlkNskbMHxhB2L9RAsC6pnM3Weiz1XN6fi977
1XrVefzXAXO4rTiCOQAI1kXykkHhZlSoOXBqq4MH8pHzc2Z6hfCU26i8yxIfb3/CIKNeexmj2hiz
ObpGKWi6MeUIKwx6xW/dXUEPYmHipgujPn/awlz6EWNP3wIrTpDEr9/P1DhvdvKWbXLIu6bRN8OR
ekXqDQdRgF4brXxkx0mqrC7RrFaol35badEO8qM2V+DCjweYb90o6gUy+MiHO3jFf8glcmPlUNW7
0nlL9Ncuggx2hq404sdETJO9j4elyDBxJuC7Ug0X2l70UB2Ig1+/Q3VS89I8VbGJWGh/zVuCAMBb
nD5xjcoqrStnOqHwcd9kJZYPnCkkWiLj87r+H916YexyyiAD44xG3/BYrAmvDM5JiTFOP4tzBgdh
SRaEwi3rLqgU2I5RTOQYLTKP4bLLyh1eK831IdKtj0gsnPNBqyprOgssTix9MgDUS5fvSzmaNuVB
lx0BiPsfFoEWjJHLtJMLEKNmrwdCS5E9vETty7F1sRYmiFZP45aAYzuw2U3GQXMBRt4Yyy3U4ItV
trdvgasySBwVEcyl8h86lNmo5/wr2mlSPPPtXEhkDPD/AYsg3Zh6hZA2gJlt0Unq1nl+KVm0icOd
2FigLgwX5aDmaKm59e0GLYJHS6/KYQrVMVH7GGiuod/+tiNjv91oizUUNy6s2e9T1z+wyEvd5Is7
yJ9jtr4X4dCY+5+x4cmM6+s4trbtqZfx6bmfw08BEyrVKuyWNo4Ar8gvkYAVtHIHfphPtXYy3XHI
Pih10nZwn3FeRsWaT101wUtuuizzoNtPhBKOZP1bpEtA39VMt3j45RMun4UFzuOG0idT4/o8qaJ4
hb2ckq1ROvNwS2JB1IGkxXlo7nsP1gvdlA5ufa1JVyieFfYXSHMmESpEFpGItDcKjlLQcvpkDdqN
hl/En+JX+Oy38X3/fRyDLILGDYC2QsOgPFDN0AdWQ3sRcrbbBANTgdDr+Ih/StUwcxphmCB1OsAr
OSD8sNKdoyJtmoU63dNjWw3tkrSGa7ST8ZxHmRba8pCLzMtriUYJEH44c3G0dFwg9Z3/eJkbAI/V
pKSt1qLrZjDVdhkvYvEqI6QjMOQZfbPnpJLmRsP0nUCfZmbK3/zmNOSk06sNTEU8Mm3z5ctx37TX
hpvOZzAdQDdJt3t6aHp7W784gHOrEjAVIkbbbAvmKC6HjOoQV1JBDhic/RCT3hZMxeghUGSYC2UY
BUzBRU8jVPnEZ1R1r5zbvJ9FifIXzDJnk/+IPJGE1EiMyOy0TvgxsQYJIlxP+my8xdp8Go+tymx8
8ZxJK9300lXszUVdry+N0aLU/QofG55JcRsV0hyGmtsrhDXzAsW6v/yw6VKLCHhBGct6MTHs46+q
lyEhOyjFX5pJNWcNnkggDrVgBaGvoW9VJqJnfsT5yyyqqD6KnyH1xjmMVgQJcFqekHyv+54Ffqft
aIsafjCzsz20yc0QQVIDWV1afDUDFnq4kqvJNlgdR2KnDjqPSiF57xWWx5I8h8DhfxRqckRTdIuX
XEt3HIJiSSgvFNuyJ36AInStZJBq7mwos39WTaEyvbQVIM+k5dCxpnKL4X7p0G3e/EKRzcIO4jIu
YU0LPCMpUP5I72XVfbCM7xkD1Uz3LMg2A1gw61SylbbAXYhUpBWFnmTJSpKAOsm8MPQHB/9DzI1X
RVRKO2II/Q6wmpWZvcn87gPKcjFyyXNcoDUOmvKGXEuR0mTJ3uKVZfaDtVJCBR1HgQmdOIWDD0uB
pw6ZwaPXs+MTvgCncAEGMnHPAwP+sqQUIKvPpNzIO2xemEJbrBIv0CQFJGnPKMKlr1T28FA9OiyP
WC429kkuBVa0GezownAtNZbfpVUJ2yGXzBoWRIkYpdzktgyxJfw2sYbIFZAykxP9eBSHzGTNgSN2
edHZfEFtR+M9gPS0H/O4M7qcsAMIKcjGFyJPDGCRcVKizbWQtj/Hhyv3Shxv2z0R5KvNpke6HDkY
gVuvEHLqh08Buj1T4eu6Aw0F5b6LqVVKW3ppXvwgr2oUXq7CtvnMyVoRzJFyxBfnA3pBR7hVrAzZ
LpKaNyfzFz/nUIO29pR+1iYGYMVWIoHL4xoyupAUENK1yFDFDx+Yr4rkV5S6QrFFVDWaHUM2+odm
4I3PV407ieaqLMu9jU5OW4Dkc4XGtpBirh47kD9PdcaUoLbX7qpfQ0jhtHjPzXqn2TJ9vkvZQVGy
rOOZNnmOagz9efYL9QRuV2hXf8aJJ2oKorgV+bszSbcfwQbqNmV99lDZQhe+J1608w8KZEkZrMWq
ufylt2ppGSFdxMhjLTVt6VwznDRhf3NIkqRy1GD/duRKTbQtoKh+1g78BBdF/wYZylo1NE+G1ONe
RGRwcq4BftVGAgPiWqOPfkyvTBb4v8LfVE2+aJnM5/34NOnSzyBWZdNAcRx838WTcLd0jdSgHkDC
v9duaDA8yGHyu1ijBrnOUpSoODlTJMnL76eoOY4ImLDd3lMjHlGHys7uLOQfqgC9+wSIBi66U6/Y
OHWQ0WY9jqxeCnvQg/5+zBpQJ+3P0moGEl80WoPoz8WMTL3nq2GwkZdyHIkc3pEam3l7b7N1MH1b
zzHwkBW7pbqXkfTPiEy/QY7WQeqdTzBU/cr11Z+9xU2q2sbDG5KywAh6R5gDtYJ0E6awD0SeXNvk
qA2acBX2SLpqCPkyJDGbT8SlLpTGUerSfVVdPc603q84dhMuyIrvTadAZxPoUsp1qlxQx4jTi8CQ
7PbPDdOp0upLyYWgbtxZbaqGvrAH+6RnalLarUuH9rQgWEk+f9ibWsRc5GtLoaE+vWN5Lw7RAUC2
Ua8Ty7YpXjcWDlrsI/VMDvxLgnP9k6i0J1H3hmNLizrPXoToUHK6mgsJjlq1YI1W683RHRG7pSVC
r60IVrFKQ2YGjafaD83khiEIudWhCCGQ5cjNTToJ+E4TS4Qk82Onpmqdjx+32Or13GQFqYm2rCUZ
qIBi5wRkf3ZFziux3qaJB+RanuCPbMplsvPQwl383Ho6A3SprhshGWGUJdt2g+bknbQ20+fU1aBH
3m+h431IsAb8ZTe2HQhl0yDRvcbarWZlFyy76D2fcf5PucuQ93LdFKmV+pZpE9BPZI+6O4FEZuCN
U5HwqkRo1HG0pimaFTYIH3XvYqawnZvIlZOWRSCM8wSE+kYRQrob816P39sDoHQna8czr/3KSePT
V5AJpizPaWkjvg257K0z4Njrk39G6jqsk2TrI326/7EXBQEvbttbsDFHh7lFmYTchQZebF2utMqb
neOLi6rZpV7g8czqgaEN1bqxSFxNxq6/EOAhLJHVGsMcJeZfxkO/n2NI4bhaJB7b0LI4rNelgDKK
UQuz3TUXVud5GG7zsgXF/UO6yXJLFp+/iDYgFZu64H+kzMnhXzk4Yi7OJ102LAHlghC2EaRyhM3V
aIrQU5M2O0KEh27LNT67BHBMrx0v9dbIjNaSvnokyRnazNgxtMttOpDupj2ks2BSmN3YCS1YXtoi
L/Tfl/ERB8pBGuOMBu9uSVcMfz36j5+BiNIuhpXc8gk6O5k+lmreZfkzinYjmzRFwaOUMWRETO28
yTtFl2jdbJSa50lf1EqQLk6DQUdCkxcPpl6dfr8fXoP91jUTnanX2Sp4mZWa57IOjG8A/Hr9EzHq
TFMP70vFaSe5bnTJSbIQIGqXGIXuBntCa5Dr7zo2dz1fnk9x9U3WfKuMjMxqVI5S6+CpmEXmoYrY
lIBxECW00p71ZRYyZDgE9fxgjXHRzqJmkBGjKpCLNjnxGrpF30n+uZUgx4QFQbOdHjbSEAXFlSgv
ufU9tWRAAJiLGLu/kKMbVlJovh/rF3wBKUlkBLv5ME2H2yEso6PNYegpmXtqO/I0EwLdmqQD9O99
9tfH7WFsWihMi/yzni5K+itGGRwOatlFJRtUh4DwwlpJ7HzTuU2Oa6RvOdxl1c9JQ70uZxH3IDxb
rQehncgtS49La5UCBXkYXmS1Os7KmNtKnzwaMTLlPdPz8FdHpzIHJuawWhshX8qefQtUTRJDhrSs
gVfvf7M9FQMEBrdsaGueSAnwuEdFGRWv6euqMVjp/zCuyAxSfX6Vnpukw6IyuO59MHosHEEygpmv
qjnYC0jhyOMrbgcq7vH/E7LrKsWfWhVp6P54DC+1ntzeENqL5OjuGPnJCyk2erzS5jhWr6nUYTmk
xUYQ1oyOS2BJ23MCZqU1JUbUn0xGKSwt/DzhZPhOtqyNvG+2RfX8+qJUiJk3ffGF9gr7foIVS6D7
VGne90QPVrkZmzdOp+twb9m4CQVSMlTw2gyBVcrGcpwdAqdM80rSW0kJi1Oi3yb5lN6UPRkRM3P1
TF2WktrUA/MuRm5msjZ518ZVyCMnr6vJcvsy+kdy9nMeA0iS8y2upr3vgcEPt+ye6w9/wBvlRVpd
8yXr0SaUDkI6CEaTrdhQH+yM4C85FBE3kQXIrvBBoC2NUr+OVbRG0J8YCogzV5o5ZhiUoqB9/dAG
LikecVjNgU/TO1ziG91xVZRE1n9JUssYXi/1E2y0Ej/MB1VuVGrQmUlsegcSCGJpwH90AoYyLT1N
n1XZzMqkSJUrTPb2nOgUCPbqX1dWq7vAsQqbsNSdBk9C+0AgACsNmmKKEYKLizz8Zjd4aHu+RsSz
FbKATPxO/aXFOvkdQ+DnYP0LjSmm2NKJEccWl4hdMXAQyu8ELcPystJ6rZKtULXeQw3wszJkujvu
fjMowiWYnSDpNil02xiCuxsD1zMk8wO/5rLNCF1K+6B0e8tQgahhYimsa2kS3L+PGa+ZYJM6KJ6f
S2KVECPhHa8DOG9ZtZvqA0rkQbRHKXAsJZ5XwNWQR5CaK9ErncRJauNhC05xaRNuomOoQPrnhENS
pXmTVdqmfibv2u9KfFn4sKqwpURzw+LQbkn2tRnwPLXJ36PV2MBD/2C199Ih+upI+M2PNCM+OfGx
PjrZ/nQeoXVa19IpBvKyTylTp/mvcFn12dXgZZ/GG7SHPGYm3YcuZr9fAS8Jm+bLUH6hJDa8FjNR
gCi6dWj4usVF8PHcaTvmWtbmawMVYq1hmQocT5YgXscSj82wghQeXmEbgyq1I3UfBkkwpjzAKo4i
bxiwqw/GO+pJu16y6NWOobjXjKFR3mssgdpeV7I7OIMyW0GFog92lYtc+/BvufJEJXp0fPpaLXxf
m+XTaKEav060ZBGb86Iwa2IYjxw0G4Jv52lDsxH4nJwYRY9QkF956+HcKK9e+ZVfx1pFxeuAwZj1
s1eaM8mufgpue0dtvantZCdND8lRVGd7pgGxRh6vlXUcyTVFyNicE1vEkAfWFHRmLCg06Jfy93b5
saWaBAONdNSof5TFvFh56FY+cftbQsI0FFwHjjC9MJTDms0z/ZqHaNtbb49YRLNCX1v6+IRUOcXq
eEgfT/BiNMVISuwNXcH07JTAsAtl63O8eFbWQLHWcFYEhy4HGCVWLFv1FRy/ll2pzGXRM6Wlzc8E
nxaFMJEylmRw9BkYmbr9f4Q1CuZpAocwCzG72uvA8Rwv15muXB7J7M9ojDEI2VkVSsWOiJix0kP2
FnrSCd8XRzkNAJ5ryiRKmiU0uO53cTFjEgmP5X5j6jAFl7tegWRBtH3lpicDVrQ4EcMy0sXmV2H4
WhdOjUBtQPMiT6q92QzQfb2UOMX74fLdDqTxKj8hnAx1b/TKf11ILPuPGbi5BL9A8ce1BReOojKd
oFQ1bQyq/QHIKi2tomztZTloYp/58CE6+0OP6An3z4P0ZcmUou7r+OclubWFDa90u95mTmvt1VqU
N1o9awOfG6Clhk0NaomKN+rZVIeItdMkMUw0EtvfhmQCABmw3ftmLInEL1r/JZA4osHDQLXPn8+f
oo9aypFTe4/7lBRIeULUgUjOnDw/AoLyFKj1j4B/zqa8J2HZC28IHTilNRWmQpeBOn/gNPZUKu9x
Og656Yhvm0jwnGl/Yw24agK4C3gfLmVGnPsP/t+7itWFCbsMH+hWw9HD/zcjdOSs5jSjauDzQ2aS
0+s/vDg/He81I7zZE7NImgugmJiLk0cpGO4Gi4b6bSO61dd13NxZKssg80ItOgu88c5d6Zbm5aR3
Keg374tDW6/+ccUY7FlCejhEJWDDG0vspJd/5AFzujv/j2lZd9mjC79WU+XNKErrx3M0YbDuD+X+
W8xr1VvubUI5Cw8HxQJqum49xM61+2zF2K7AD9K0fc0ruJeqVbWupzQp7TFjrYbjpkAJ1nM8E4Jy
cswwXKzffjU7YwDtHzQQ0HQWZ91JWF5+yDwsDmR4USP9af+1FkMTmAisoLhdeuFeQVX2KSXXgdFU
ZB1sSNIHRi7+E/9yE4V+/y9s0Ics03ChGA/N64zb13PDcjMWJdK4qWTatyPXXqlKP9RTvezzsZze
K/oTSjU1bEcF/mIatELAji5brFOiq+iILJF6CrofCS/DsK4UfGpt1sqKs2zAErVmxd9oMhbAcleZ
oa189Q1bSM3yKeqvZbuTdrxekl7MXAki8d1pnGBXBHcV3dRtM4z9PI9RzTHfpxrpNTGDizvJaAG9
sGbczgnS5obxI06rF8xUIUtFoyOk2zttfXbsQ/aUK3V9usR8BJoiJlB6fy9rGxKeD4NsxaOlHjKz
oZCocoxT1RJ1dDx4BYNX09KlZhGSKtwhkeLWk/xHjoxoc6PRuSiMlPPDm7I2fGCxCHMI7ieyfLT1
XK5t16GqgdfUNt10U8L7bIS0ulE4RAMCP/uR7mzNT93IyqdOg9uQO0QPLAeZD+OJXWd7hpmJS0+7
vnU78HpQunUguQDtBkpDkxf/x03MnOG0I8a7DQkSrkEWuYr0VS6ZGKVjkQ8YsZc/4upj2xAPC2Od
eBfNN2NVrZdJJek2G4SO+Bb83QWkx6sTie6rybMuo9rmm2pG0dhMAERy2OZ4h7eh92nZpe5GuQNu
A53YgVpLO/9HkVOlgbncNTRg1OhEuHymBmje8ym2Bo7ZTaX/qY6R07DWN07/Nr3oAE15nGgzyvth
8JOR6oI/6vG7eYlQ5bGJC/v1zwY2wt5++W+Zpe6RhGZ5Beyc83/15hXHPgAiYvgz5h+HaeNU3Wwh
eCBPEw2p/FiAPLQ/yeM8rTN5aVKczt6zk2WxXIaXIYwtYMOLO6uKQ5s66t6RoIwoN+7qGv8d82jx
wRWkvXZV7jhPn7SSSgMLrt1Lv3khwFtIX8LMue2TzT2UwHT+ewfU1T8M3TNv2zEed3jRdIUwsJnx
kOM1aF779cBXd2vFWLi9jVJqkHJtigAeHyXJSaT+N8OJ2aoKQ5+gjTsTgY337jzOhDaXtWY+13ww
N7qsOWC2Lcs/A6GrS2d5rgGqYrOJqmxyDz1vaaF7nWAjvOH/vQ7xtKhcCN3P6xm7UbX+jbE8YUA2
xcPewmBaFtcTbxtdgL5O36pRzKE5jBpqwf/+mfx/0frXvmN9H6yAIVy/3MtoLDRQl7NmpF6pVVgG
1H08yoLOZu7GtXXe3allTLWOgAOkg2Yvw7VdmoEIXmIzulSSUP+96uPGYXVTb3YjCNrEEX+XjMXD
y9jYGC5J4uqNt9m04A8dsgyPfdumBYS1kCTjg4CMF3uD7+K3fXpjzratVYOfVFkD3eZunA/nDAls
6bD4von4oIlmjvIeh386Bvs9CFs/gnZXLf+9fRP5Xe+WmOLOLN2/bkkhhB99Ui2U+0jfWOH8bOMb
81FbMwW6xOxMMlHe0uNtz5j4L9fJd0TL85Q00GCS+PaZhZl3XjGq6kaOzOLPxGPJmV9IY9tCQZYo
4lc4ZsP9xcfAnzqmCUarMKSd+6wlcWMzh2Sk5HHJpq3BEtJEhpBK+DLWOJHJKtKi9AsyegNS8RSo
MDjfluwMZXN8BrKNj0SjQqEdHL02J/T9X3V8c7QjXIbiiJrP4HFhe+qk2Ii+maNEMNcvzZwvIPA1
OpQkxA+hjwZXlIEOnWBCDXTBFtrw+hbdPKYxL6kF8TYhUinVdkoP+21lstE4PqI/GG8tXO2kdwzB
anEoDthFUoxXknLj6mhzSRK9v6WzZwziF2aVk7szNEqp6pspJDyt4yH6eOFbDYQz4ucF0vo248hC
e1Apgnx/4CU73KP+n27VjywcXLR4jTEZVBzUbEoawnCL+m0a1AdS6cROu28FqKtXaKpiREtEtLuo
fb0D+wpnCUAJzaudlNXLkL2Pc6iNJc7P/GzL+HeixK0g8ACgNu65Bt11fhuLTmJo5H4Bj52J9m+J
PGkKYp4YGrDTrHuGX6X1VEGgHX0R2k1m7RDP580HXJwjR3tWknBF11wq+J+17zaPNzQdTkXmjNL9
CtgAFrPUm2nWQaWche4i4aoEcwH0py+vpO98EbYkR7UGIg5OQw5fCoeSz5wo66qUOY3E+vqBDRHO
zxZw9+/0QytgwgMwm0lMTOErjvNc4ekka7BDrBCMcv6tmlY+bbSYyljIXRhZgyx4QWVSZZzI6zw2
mwXn8CqPiC8TfksIXG04IK5h8UjPyczVASkuRAqID8ANgwVsqmrWkAEhYNsEqFsBtchlna6gLtu4
Ogm4i6HX69rqviUcULAJl27Nu4jcTqGVcJ70bt46ndl/J+3ozOBzCyIJGLiwxr2M1HOgSS8TfxKB
mriqGEPP9PqfbyoUsUDR+4fL4dCVVXzzEO4y/SGaiMwM/MVP1J8xE8eTvOLpFoSlMUcG4jHvoqe5
bY0CHMOTiJu7JJ+/C62vBAJHXpVSt65137VmsIrT4VPX+oQTsZis4LIS+6dzVtPgQuGrYpazImlI
ziZLgq2FRfEj8uXWQDj/uQxblrp1mNrysZUaCXNMjNtpqMHq+jRQmSX2HlrXYm+WAUV93BMC0X6e
zsqm3tj3zMB/Ji9z6FzCrTgHtpSAZmFYTaJqJ8YKYTs+74lYteJCZfJ1ZEgrMK5LuCfxb/kaHnqJ
KgxgJi6an8wsyKkZ8ZsPBPajHQ8d8Kc7z4gX5UE7Lvdi4T4+HKhs3K7cLk/u660VasYNmCiJkC69
/kZ6u3lMJTvcpCwKhvfhjJ0SZlRnnmHj9P8IIIeHyo8/hRZx3rZ/wUONDbOjYFCgSPdgkTo45cjF
gCBrbC55fUiHuWGKN0RdxJT3zk/CiKPv5orkcbHEK54YPWEBO81Uq6y3wop3KJNzziEgdHxzetLO
1oiSqUrGC2u5McohBpnDO5In7xfHEdzwLuUW0cTdjgvwXWBhrpUP9JdmSqi8fXMgFh3wbaM44+Av
S1m9HXHHqULpcbyRRyp+yrGrCOAFuKHpBz970IBBuM8rBageCXIF6i/kgdTXfn2/tNThluVi9tiP
vDfkTeMp3XpzO8/M/KKUl5HYR5m3D2HOsEYcxuE4JyL+5W+e80UNzWNuK9rhr9eptJQ0OGyCejCI
e6Mhj/4op+H+YZu5AATJuVRgYzu6Os4inNrMBvMm4PySk+aXWYITqF8Ue+IrN8KYrrZr0ts3v2Ke
E0U1oC9T5Neprkt1UwRow2OtvWIb5SgtyRVIM4ZEyxa2JpU7d4WLm0UIuzlmfu3zq+hns1+44Vz7
+9w2euktdI1UytACJ710zOQY8EEKfBIm3ns0OEpTLVLooPUmGkZZCeq2qnR0penv2WMmYnS+qgme
mmyoh7o+lnCD8I8CYlLxqc+EwZRVs9a11bUk+39Ow1G7RefR9VwwHiBXYnCTjInNF2ccEQfrEO88
bhE9iKOKDl/rqsq9gjcoAMF109uwmBOlfOHqdzVKoLIDB9kD0HoduUZ2ZdaaNInM3x+KC5P1H4nT
i07UA/QAxw4VEYywukcfJo6XvuQkXdX95SgLPuyf9bzLzAn0xyNruGxc8pVTsE0YHJQdDHWtyPRL
qx/wYdwku025FWSjd3z2WEggZNbh5OPrfaIDzlBKy1lZGN46wRpIkATlFOyhEmo4DbDFoB2gKHk3
/UQQAHdUXyR3ibWZaHgnJUkvBB3gZfnFoRNhZfabn7cwOCO9Y2/z9iqyHSMkqaOk4Aj3tZNCw/4k
vB0zLa6UeYo8Uxh1qjWbVHkZz3mG5z5XpLBldZ0/BNFxxIQBy4vTXNQ9dmUjs93A8rt0KXjUzP8+
taGeS9YoVWENRTMyCllj5QYhQ1aKEkBueYn8m2NJdtOEIts4f96H49sxYUn/1331nzkda/+3y1dw
c8tJiBIGI21wHGMXwXNlvLIiER4dbujfxx9u/66ZcffS1omdVdC1KDjwOrX7ijMbHXPEEytKeasM
pMwoDKWrGJhIZtOd9ZggxY0eLM+Ed4CUEaaGz8jdhn+skjzeHWw05v/rAFSrapX3xYVDDm08H/tK
YPXVHWSgEKH7aGesAMUckvWOWoZASiRxMEDixFmoGRxay8OOSUNYYbaT7Nt6L0hq5IuODZqYs6HC
HYZbGLz27+ooolT/kuGN4UCHkPrulPeJoJaqdGiMePqqHU+gaO3dX7xH1AIUZGt/j8f7hfKReIeD
dostudmNIbfvHmjaEm7/mfTfEd9ITFta2B7XVSAAwtMM4Fdk8qJh9x1SxnGSUYvGbd1eJXlj9nDP
TZjEgC2Dj2VGGGYK2BvwCQVC1SDFhvJHJOeH4HZa1AUny4G1OLVoMxnH/cZkqTulEwcXMs2qN57N
nNGtT4e9m9rnewVvQLLPhnj5/K5YjiN8QWYzImtw2+29czaShU2e7eZmignDIWclC9BBTvOqFrHx
EAlk0jWrGM6el7Er/wTjoy8V878v5qxpksK3ppbzr+PGwJOnzJrqozIKO+e3fLHsyuxQmhehArP0
BJ5M/2F1Irx9ybEC8969rEDp/AB0vh0XZyzLat084Miv4GW6zMIo6hRO7TUvHecpqgnz2ED2Qe25
RPhwiC68MKbtbx8rCppyC0iJtjTrIyeeQ277zd5VsDH+uNGa3Q2Mbz0mbEuKt0L/aFjbcdK+Rf+M
3b9DYoSq3SJw+CYEblAc+C2tkauiuJ0JLIXvrErCDTHXSeeU4KD1a3ao1VtI3CGHIYnKMwj+FgzW
W49TqxEgvSvjcGArk9mZCqNjliNp5BYtAkF0r9dSGKRqNYtxUMadeLGZogZAGwZiBaEAMBx+RVkk
i0xyMzUR3F9VVBjRh9F58J8ptY5EiE3AdkbTBL6J/LDW/MQX+JEo0yQg1NgjQHVVuC80068KwKoG
cJTgUID4J0QI8Ktxlofwxu3RZJpgfOVsiCzg+aFyV8VYkFZkm1fkmqQxnum07zFOxumi2ctlD09x
eVX7/oRUV/C+3NMTciLmvEzrv4BSY0NPIIbMNYImk82iQyA6gStbVL937SJK/Duvs0ZYP2KWoObf
N7iPV97v0ekvKMPlvWFdo64f87wemAHtV0VRIhAP+J+h9kciKov8w/nJ87ECvUJH27NeXTOI+0JB
/A6JsW0t2TsGAvXh4kE4zNOQMCSbDS6zKJJk+YhE0APYT+/85fD4tNuEKKWg4wVXFrtJOXM2dlVY
iD/gsQro0V/x417KhBGV6X2/KsoQKbofjordWxsp+OYwaRRqlJeCIe5d4j+tYOfV7a7549xKbXLa
pJi7Ue8SR5QaNhr/F1NANhUPxVjbKROdFM9rUm9hPIoVTytfjFn8yqWNqfqIWwsHrBJGYjl9IrHj
yAiE12xd255dOuwhU9n8HvnEDHFI6s6zFPjbm7tl1eKn+678VZswJw58lT7vgNJINuEHKxML5IQB
luQn2RJPTg7R5Kfw8pdd6frhDLnEPeP+c/dQrVPGYN2+LJlMTJsWAwyQHkkxjBAuv5tFoJiEuzIL
Vt6J2G97JZehAJkSVuV55hsOFyKOnQTFNIEoTvE+PybYB1ZioFE0SbvPQaFv4R/S9vu3p7entU9C
QjeDnsNJX2ATS4PcjUApGTJk6nt6W05LdFcQeT7CE1++KhbpPA5gm8UChpohmNxLJXoEayFrfR2t
JwtFNinm5eQAM618ZuK8Vv0zfMR0TJOqCwJzjIAY0QYnPbN8R+zPGnGbAMT3ZF5+b7H/pBaWV32e
2yIcn1jCa5uv36K9rJdORNNFO/m/nIVRaLliDSuTjwLPSh088YbhfBEUgg6UIoJPeLNstn2uACrS
DXDt5aIn0TawjqpvtPRTdq5EUo/JBKXpiW9fuwd/6G8jlAepwddTbh0+P/Q6SEyNo/t+Aa2Rfw8X
IZ5wP3ELTzGPTvMH/D9szBDcisUf/Ufrypt0Cq4CFLWsIJcJL8FfjeO/Io//K+mWXU///i48hPHb
kJJux1/oR3pfK34xIkbxg+9SEg/Y/QzZTiXhptUrNW5mmahUOKEr5xuzjbg7W95Qch4p22AVr+71
nFsB+trZ7cWR8lRiGqaTuodIk2gwYIV3kyzdCsdMwsTPLST6Z5KaGz5z/RB2hsi4zuT1e2+eosvE
L6BJpqaAnEArWz8x+jP2b73BU8dsHglkq9ruspf8ia8I88EokNcwKg3pfPo9HZ2XdDScF4At2DEf
9QL+wAj/nn+lvPXS3aDJx6TrR9oqas6SpMtHglAJFArW02iKs6oeVXkCrZN8a5zfcPWPG4+EAQNy
9R1MIkFgI8tTHuAimCe03VDCtxBo6+qR363tdepOKQYGchOfwWhmawaJXtoU+39rb4UgsI0MOBq+
Em6oYtpeZZE1KN8NT5BHFBaN2z22lwdFNJTvy6w6D5K/AflWkmm6wXHk5zCBSzBqk7qqbMQcKe+p
6tx8H75JDNex+uAXT4B24gl9cUmSGe77BAKr6y6h+Kny9FVxWrxwCXpkz17r7taJq0lUhNNDsiBk
tpv4SRXMu+bSdqO+gUrFDXUFL9NeqsnzHgoBvIpLUC+UFiCtIEITR5yHXGHcyu/pW9j/fG4BGRQ=
`pragma protect end_protected
