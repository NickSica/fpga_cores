    .INIT_00(256'h01ba002da0701f0101b900205f42ff000188402db0701f00001200205f428000),
    .INIT_01(256'h02f935013002202a02f834015002202a0112010146c2800003ac16250002df02),
    .INIT_02(256'h036c10142002df0201d0000d01001f0000b0130b0142202a02fa360b2152202a),
    .INIT_03(256'h032c13143003201d01df30142001d004003ff00d008206c600bf391430028000),
    .INIT_04(256'h01d2013a61632544022c01190011d001032c3b01101325bc01d202030071d002),
    .INIT_05(256'h00b935123501d00000b8341024032091022c01226121d002032c3b14106206c3),
    .INIT_06(256'h019402060101d08200b43c09008324dd02f20f2d2091d01000ba362d30a32282),
    .INIT_07(256'h03ec97250002800001ba002d0082df0201b9002d20901f010188402d30a32225),
    .INIT_08(256'h00b20f14d002202a00ba3614c002202a00b93514b002202a00b83414a062202a),
    .INIT_09(256'h01480814f0e2202a01490e250002202a00330114f002202a00038014e002202a),
    .INIT_0A(256'h01490814b08206c900039014c080106002f80d14d082202a02f30c14e082202a),
    .INIT_0B(256'h0142063900020697014308110b92068f01420025000206d501490814a080109f),
    .INIT_0C(256'h0140063e638010c000b0131901122ffc001302390002066102f20e190e9206a7),
    .INIT_0D(256'h00430025000208d8014006190f62500001400639000208ba0140061100701101),
    .INIT_0E(256'h00b4382064203cff02500000c0003dfe0370002500003eff02f30f1100a03fff),
    .INIT_0F(256'h01ba002064c2003301b90020642207a2018840206b5250000012002064c208e8),
    .INIT_10(256'h02f93514c060110002f8340110020037011201250000110003ac48206b501010),
    .INIT_11(256'h022c3d14c0620898032c6a141002500001c2d014c06208d102fa361410001014),
    .INIT_12(256'h02f20f250002003700ba36141000110000b93514c060101400b8341410020033),
    .INIT_13(256'h01b900111302500001884011107208d10194023a64f0101400b4381d10a01100),
    .INIT_14(256'h00b935090060110000b834206b80101803ec9701a002003301ba00250002089e),
    .INIT_15(256'h02f30c20620208d1001300011040101800b20f390000110000ba362062e20037),
    .INIT_16(256'h014908001000101c01490804a002003300039036657208a802f80d1910125000),
    .INIT_17(256'h02f20e3665201100014200192010101c014308206b5200370142002064c01100),
    .INIT_18(256'h0140060112003fff014006226b5208d800b0130110d2500000130325000208d1),
    .INIT_19(256'h02f30f0113e05f00004300226b503cff0140060115f03dfe014006226b503eff),
    .INIT_1A(256'h00120001133208e800b403226b505c000250000113105d01037000226b505e00),
    .INIT_1B(256'h03ac75011310101001ba00226b52003301b90001130207a2018840226b525000),
    .INIT_1C(256'h02fa36011330101402f935226b50110002f8340113220062011201226b501100),
    .INIT_1D(256'h00ba36011352003300b935226b52089800b8340113425000022c6c226b5208d1),
    .INIT_1E(256'h0188400113701100019402226b52006200b403011360110002f20f226b501014),
    .INIT_1F(256'h00b834011392089e03ec97226b52500001ba0001138208d101b900226b501014),
    .INIT_20(256'h001300011422006200b20f226b50110000ba36011410101800b935226b520033),
    .INIT_21(256'h0149080114425000000390226b5208d102f80d011430101802f30c226b501100),
    .INIT_22(256'h0142000114601100014308226b50101c0142000114520033014908226b5208a8),
    .INIT_23(256'h01400601148208d100b013226b501100001304011470101c02f20e226b520062),
    .INIT_24(256'h0043000114a2f01e014006226b52f0320140060114901000014006226b525000),
    .INIT_25(256'h0012ff0114c09012025000226b5320c40370000114b0d00802f30f226b509011),
    .INIT_26(256'h02f20f0114e320a902f20e226b51d00402f20d0114d320a002f20c226b51d008),
    .INIT_27(256'h022ffc01150320bb022ffc226b51d0010250000114f320b2037000226b51d002),
    .INIT_28(256'h022ffc011520d040022ffc226b50900f022ffc011512f001022ffc226b501000),
    .INIT_29(256'h022ffc011540d080022ffc226b536112022ffc011530d020022ffc226b536112),
    .INIT_2A(256'h022ffc011560900f022ffc226b52f001022ffc0115501001022ffc226b53610c),
    .INIT_2B(256'h022ffc0115836112022ffc226b50d004022ffc0115736112022ffc226b50d008),
    .INIT_2C(256'h022ffc0115a2f001022ffc226b501002022ffc011593610c022ffc226b50d010),
    .INIT_2D(256'h022ffc250000d020022ffc2d10636112022ffc206bc0d040022ffc226b509010),
    .INIT_2E(256'h022ffc2500001003022ffc366b83610c022ffc0d0200d080022ffc0900d36112),
    .INIT_2F(256'h022ffc2500036112022ffc366bc0d008022ffc0d01009010022ffc0900d2f001),
    .INIT_30(256'h022ffc090003610c022ffc250000d010022ffc0306036112022ffc090000d004),
    .INIT_31(256'h022ffc030070d040022ffc0901336107022ffc250000d080022ffc0309f0900e),
    .INIT_32(256'h022ffc206c30d010022ffc03160360ff022ffc001000d020022ffc2500036103),
    .INIT_33(256'h022ffc20685320d7022ffc2068b0d004022ffc2d1000900e022ffc04100360fb),
    .INIT_34(256'h022ffc206610300f022ffc2063a2b04e022ffc206c02f033022ffc2066309016),
    .INIT_35(256'h022ffc206c00900d022ffc0319f220ea022ffc00100360e9022ffc250001d00e),
    .INIT_36(256'h022ffc206851d049022ffc206a509006022ffc2d100360e9022ffc041000d020),
    .INIT_37(256'h022ffc326ff360e9022ffc1d0011d053022ffc0b032220ea022ffc20663360de),
    .INIT_38(256'h022ffc2500001300022ffc206610b202022ffc2063a20661022ffc206c3206a5),
    .INIT_39(256'h022ffc01002360e4022ffc206631c320022ffc2068511301022ffc206a52071f),
    .INIT_3A(256'h022ffc0010020661022ffc2500020691022ffc206612200a022ffc2063a20716),
    .INIT_3B(256'h022ffc2d1001d002022ffc041000b002022ffc206c020047022ffc0319f2003e),
    .INIT_3C(256'h022ffc0b1321d003022ffc206eb0b002022ffc0100020050022ffc25000320f6),
    .INIT_3D(256'h022ffc2066301000022ffc206852085e022ffc206a520059022ffc2d103320f6),
    .INIT_3E(256'h022ffc010402b10e022ffc326ff2200a022ffc1d00120716022ffc0b032206d5),
    .INIT_3F(256'h022ffc010202b20e022ffc2500022110022ffc2066101080022ffc2063a20703),
    .INIT_40(256'h022ffc2b40f2b40e022ffc2500022110022ffc2066101040022ffc2063a20703),
    .INIT_41(256'h022ffc010402088a022ffc2b04f22110022ffc2b08f01020022ffc2b20f20703),
    .INIT_42(256'h022ffc0100822110022ffc2d01001010022ffc0102020703022ffc2d0102b80e),
    .INIT_43(256'h022ffc2b80f01008022ffc2d01020703022ffc010040b001022ffc2d0102088a),
    .INIT_44(256'h022ffc0101020047022ffc2d0102003e022ffc01080221ed022ffc2b10f2f01e),
    .INIT_45(256'h022ffc1d00020050022ffc206c33211c022ffc250001d002022ffc2d0100b002),
    .INIT_46(256'h022ffc2066320059022ffc206673211c022ffc2069d1d003022ffc3271d0b002),
    .INIT_47(256'h022ffc206a52f01e022ffc2271a01001022ffc2069120703022ffc250000b001),
    .INIT_48(256'h022ffc2063b0b001022ffc00c300b237022ffc2066319801022ffc2069b0982f),
    .INIT_49(256'h022ffc206a332137022ffc206ce1d001022ffc206da3212c022ffc206611d000),
    .INIT_4A(256'h022ffc2063b32155022ffc0bc3a1d003022ffc2066332145022ffc206911d002),
    .INIT_4B(256'h022ffc2fc13208e5022ffc00c30208ba022ffc2500001102022ffc20661010a0),
    .INIT_4C(256'h022ffc2066d2fe0e022ffc206632fd0d022ffc2068b2fc0c022ffc2069903f07),
    .INIT_4D(256'h022ffc2063b207a2022ffc0bc0622167022ffc20b8b208eb022ffc2066d2ff0f),
    .INIT_4E(256'h022ffc2063b01102022ffc0bc04010a0022ffc2063b207a2022ffc0bc0520858),
    .INIT_4F(256'h022ffc206832fc0c022ffc206a703f07022ffc20787208e5022ffc20661208ba),
    .INIT_50(256'h022ffc3a746208ee022ffc0d5042ff0f022ffc095022fe0e022ffc206632fd0d),
    .INIT_51(256'h022ffc09d1d207a2022ffc09c1c20858022ffc2275d207a2022ffc207992216a),
    .INIT_52(256'h022ffc14b0601102022ffc0bb13010a0022ffc09f1f207a2022ffc09e1e20858),
    .INIT_53(256'h022ffc13e002fc0c022ffc13d0003f07022ffc10cb0208e5022ffc14b06208ba),
    .INIT_54(256'h022ffc2fd35208f1022ffc2fe362ff0f022ffc2ff3b2fe0e022ffc13f002fd0d),
    .INIT_55(256'h022ffc0bc36207a2022ffc2063b20858022ffc0bc3b207a2022ffc2fc342216d),
    .INIT_56(256'h022ffc0bc34207a2022ffc2063b20858022ffc0bc35207a2022ffc2063b20858),
    .INIT_57(256'h022ffc20683208e5022ffc20685208ba022ffc2066101102022ffc2063b010a0),
    .INIT_58(256'h022ffc207992fe0e022ffc3a7652fd0d022ffc0d5042fc0c022ffc2066303f07),
    .INIT_59(256'h022ffc0be36207d0022ffc0bd3522170022ffc0bc34208f4022ffc2277b2ff0f),
    .INIT_5A(256'h022ffc205f82093f022ffc01b00207d7022ffc01a0422172022ffc0bf3b2093f),
    .INIT_5B(256'h022ffc09e0722172022ffc205f02093f022ffc09f07207e1022ffc205f022172),
    .INIT_5C(256'h022ffc09c071d000022ffc205f00b016022ffc09d072093f022ffc205f0207ed),
    .INIT_5D(256'h022ffc00ce01f000022ffc2063b0b018022ffc00cd01f000022ffc2063b0b017),
    .INIT_5E(256'h022ffc206611f000022ffc2063b0b01a022ffc00cf01f000022ffc2063b0b019),
    .INIT_5F(256'h022ffc2066d1f000022ffc206630b01c022ffc206971f000022ffc206850b01b),
    .INIT_60(256'h022ffc11c010b032022ffc14c0036199022ffc0d5041f000022ffc01c000b01d),
    .INIT_61(256'h022ffc206a711001022ffc250000b03a022ffc20661325bc022ffc2063b1d002),
    .INIT_62(256'h022ffc2b03c0b002022ffc2b80c20076022ffc206632006d022ffc206a52f03a),
    .INIT_63(256'h022ffc09c0c0b002022ffc2b02c2007f022ffc2063b32193022ffc09c0c1d002),
    .INIT_64(256'h022ffc2063b20703022ffc09c0c20088022ffc2b01c32193022ffc2063b1d003),
    .INIT_65(256'h022ffc2066132544022ffc2063b1d001022ffc09c0c0b032022ffc2b00c2085e),
    .INIT_66(256'h022ffc206af0b016022ffc206af321e8022ffc206af1d800022ffc250002200a),
    .INIT_67(256'h022ffc206af0b018022ffc206af2f035022ffc206af0b017022ffc206af2f034),
    .INIT_68(256'h022ffc2b21a0b01a022ffc2bec92f03b022ffc250000b019022ffc206af2f036),
    .INIT_69(256'h022ffc208b60b01c022ffc2092b2f03d022ffc2b08e0b01b022ffc2b1bb2f03c),
    .INIT_6A(256'h022ffc250000b001022ffc207bb2f03f022ffc01c000b01d022ffc250002f03e),
    .INIT_6B(256'h022ffc01c07321b8022ffc250001d001022ffc207bb321b4022ffc01c101d000),
    .INIT_6C(256'h022ffc207bb321c0022ffc01c0d1d003022ffc25000321bc022ffc207bb1d002),
    .INIT_6D(256'h022ffc25000221c3022ffc207bb2093f022ffc01c01207d0022ffc25000208eb),
    .INIT_6E(256'h022ffc01d00221c3022ffc250002093f022ffc207bb207d7022ffc01c04208ee),
    .INIT_6F(256'h022ffc01080221c3022ffc208c32093f022ffc01f00207e1022ffc01e00208f1),
    .INIT_70(256'h022ffc250000b016022ffc207ca2093f022ffc208ba207ed022ffc01100208f4),
    .INIT_71(256'h022ffc2b08e0b135022ffc2b63b0b017022ffc2b00a1c010022ffc2b3890b134),
    .INIT_72(256'h022ffc2b00a1e010022ffc2b2090b136022ffc250000b018022ffc2092b1e010),
    .INIT_73(256'h022ffc250000b01a022ffc2092b1e010022ffc2b08e0b13b022ffc2b37b0b019),
    .INIT_74(256'h022ffc2b5bb0b13d022ffc2b62a0b01b022ffc2b6491e010022ffc207b80b13c),
    .INIT_75(256'h022ffc207a21e010022ffc250000b13e022ffc2092b0b01c022ffc2b08e1e010),
    .INIT_76(256'h022ffc2b649361ff022ffc207b81e010022ffc207a20b13f022ffc208580b01d),
    .INIT_77(256'h022ffc2092b0b001022ffc2b08e321e8022ffc2b5bb1d800022ffc2b62a19801),
    .INIT_78(256'h022ffc207a2321b8022ffc208581d001022ffc207a2321b4022ffc250001d000),
    .INIT_79(256'h022ffc2b649321c0022ffc207b81d003022ffc207a2321bc022ffc208581d002),
    .INIT_7A(256'h022ffc2092b01004022ffc2b08e20aa3022ffc2b5bb2f013022ffc2b62a0b001),
    .INIT_7B(256'h022ffc207a20b032022ffc208582f013022ffc207a20b001022ffc250002f01f),
    .INIT_7C(256'h022ffc207a220727022ffc2085820661022ffc207a2321f3022ffc208581d002),
    .INIT_7D(256'h022ffc2b5bb1d002022ffc2b62a321fc022ffc2b6491d001022ffc207b80b032),
    .INIT_7E(256'h022ffc207b52200a022ffc25000206d5022ffc2092b01004022ffc2b08e321fc),
    .INIT_7F(256'h022ffc2b08e0b03a022ffc2bdfb2200a022ffc2b10a2d003022ffc2b64901004),
    .INITP_00(256'h498d2c94a085c6a1130fd15a90eb6b1df1a9a4a87532be54fd64ac731fb5b535),
    .INITP_01(256'h9b849782bed6f4439fb1028ea7ab9ae3a20a05b09605607d9a922d10333002be),
    .INITP_02(256'h72b823a88404285d70b0888138bade21b4b70b0057033686d7f2b9fdc8d9aeeb),
    .INITP_03(256'h30d897368900825cac893d57d8ee442cd736163f8ba74ef2d28eaab1072c1b82),
    .INITP_04(256'h51507a64ce6d7b5c3474e97b0b3233b2302a277d87050b1a95a16bf619a21e1f),
    .INITP_05(256'h53c7c2f4c045d2e7cddde1d85fc1404cd743d7c2cac25a5cced155d1ced64344),
    .INITP_06(256'h5562c2687564d265dded5a55f9d0ca69e370de7f43614c597cefcb46f1ce40ee),
    .INITP_07(256'h4754e1c1fadc72d4f67f71c9e94a4441dded4476c1c4f94d477afbf5c5e0c8cc),
    .INITP_08(256'hfa596043f5efff6fec4ed4f1d37075c64cfd5ae8ccfb5376f85e4546525466c1),
    .INITP_09(256'h706749f4dc585e555edfcf73fde2edfcc47f4e6bde54f5fd7bc454fad16de760),
    .INITP_0A(256'h76f4e552d545cf454e45d542707a4c50fd6e735948f9f9dbc6e4ec49784565e2),
    .INITP_0B(256'h68f8ece3e959615fffdc7e5be040494a45d1f75a4c65cb4567f549e1406f4078),
    .INITP_0C(256'hfc777bf4f87372526240ebfedbe57cc5e8795a79eec470f67c41e146f1fd5e4d),
    .INITP_0D(256'hfbf140f779dbd2415cc85d5e5fcac5c7d8d2d1c943544dc4c44a5bf65c49cd71),
    .INITP_0E(256'hcbd252e450cb434153ca404a5e7b55ddcbd1dcddf4454ed1d87ee7414af2cd76),
    .INITP_0F(256'h5247584c5b49c8dd46fdded44f4a43de4c4649cdc84fde7040c5cfde49d8c851),
