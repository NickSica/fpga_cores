`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
R1WqgqFekyFBf+R1EmSjRCQxUuOx6MT9aQyodTNNebOe0CK13nDxh2Wir1luIC2E+1RiIa720P7G
30ynEHVRjA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KNMY+1Jln0fE2Hw6EJV59uwRAjQ2BHIWVdMuSpeAltv11pWP/JZCrd4z/uZcVTngSRY8jZzhCZTQ
WJ4MxCfVaXUWBZm7mY0qLw6qcMnyzincQFakqwRdOx84IckfsGjNGJ3OEjUVkf7dW/J0o6KJvGRq
A/P9gVOYmGcnWb2CkLI=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
sL7gG3oizEXkzDHancu7/45cwKfdv4EnXAdeK54QMEX/eoc5P95Q2IxqcI+tnVljSH1drXWj0Eb6
Of0W/iXPKZ8OP77HA72GpMs5rDnQtlgP3rECZlxuTJ9RMJVfJzzO19m/vMWeqMysX1t8PW29rrsf
0Tqwcs84OG2uxBTuyDEWCBSCU7Yk0aBYU4VmF2rkELqh6jo2Q/udlKIUXrwoYSdX0O9uon++5ahv
mjzu8SGK6zkA4uqzG9ghLIe8qBE6KYXQuzvdlMdTVdy8eHbCbzVTNoB6j51Qlq+S5oMMSQvxBaRz
DIAN76FuevwCbX/XKHESsvee5Sen235LJDeW6Q==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NTwqMfOwske0aroynepwGO4Lz00SLylJkTISN8LAcq5uE8ZoeT6aFHS3yIuZsI6EEE3s5mQQ8Cob
RXh00Ler2BvOA4K7lNGJUpMzGqJI7MZao2GijCVpdWL1r0vSvaacAIY9nlusgQmU63NqWs7cQx1t
7NMmVlpgPTHr3KxO5lMNWR2EuXJ0I0zOxQbbrTneEEip68PBGwJFyFdSjQNe3iwSj7O0u1NlI0nF
01F/RGHelGngznubnZikT85LEu94GTbx+WNlMlaxWaxuIaRvhH8UG7MPhsxH6x7sS5ZS9GHBkFDK
gyo/ARDW7a6331M9HUgGOcgw3trs1/Klf0nskg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
F0eZzxJQxbI/Xk9S9oAxZw5Tpi91CrcqL3BrQB2lyqn9Vl25Garq+8JIOwcSUfEju0nEdI9Cvd5l
ooe0NMs4K3iY8tnE+FiNZhFGnmyV5djhXaAeRPiaySzeXAc0nSnoahW36RgdEHyPbHBrMfq1pT3d
S/0aa8cloJNV0EZcGFq/QrhQOhscPpDi8uk4IV75ihx4K3Y6D/SPBsIijokh2lVOyPsWt72NbpFl
R1J6iXczzSEND79HNenePfXgQ1Sr+h8Z2ujGHirxn/++xFCAHxWZmhGcFFwVO7AI15b3pfNiyQF1
2SACCg7/b/5q/JpHGBLoFY5e10UGMoGkaXNq2g==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eShHfvBzKaZ/Wp/QUxGlK7/6Td59dAgzaJsrKOgtjc73r+sFOocLpKUK8YR7XmM0pkfLOBkjrXYq
jGiy10qSwBo8l2eE17VZo8T9nQ0IB2FFGgVl0zNGiZaKSzE4a7K5so8c5gtUyyVlyHWXKqYAj6Ro
NzUEnqMqJPppbTPQbvI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
VtDvfrNdg+YlmytFZV1nO9Ch/hNzGllGY3c+wOLUGxBvYhloxzDDcAB/7/ljwrwghZilvxZm/DJg
2fzdltt6rugwiyCDZPTj9bYqZhAAM0bSdp5YpZP0gTz8EvbCxUo8+Op+ufZee7A2QX4lG973f4tu
FbV42AkOjECD3RCU/zC8zhB5kCMonmYQSEe1sGWBe2+Ga49sur53s1VC1GSUOY3PQLHNqtwSq2Ra
owo+cSlmwu7mHpq7nDvHG8vWLm58VKt4pglBRfC9BYdbhmSQeWT4IcMsVz3wzwUMY4HmFkj+0Htu
JAA3fKLFH4/svF3ilwX+klAmiEhOn+ftw2QOyw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HHgo2A7au8S1PE/PLf9TgssZhqFUk1LyRHoBPoQd7KZOhYH8iTwJV9W8hjvxzC2Na0peqSJ5zF18
7DRfKJ++XfNw8OtnyxfjOhMGRjIzpk9/xlZOxoCpZPFsl6WTW8CoN0RLlh22HuIAeiFQu4jBiY8s
f/eG3F7z8aDUIS222+2y8Lc0ifWDx1YbNoJritsavlDA9L9WOwq+EXi3pvUCyXszhqfkMn1JVCVR
qUhUx37i3M4UJEKXpk5rfAol3dwNa+jlOtqwiBj8/VnhZxY2i53S+bX3OP8N1Zx5wRoa1UkpaXLd
9XQOggc4VKKTgU9CJZPlRk8FrwN41qv2G8xfRQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 10144)
`pragma protect data_block
eeCl3Hcc/V4mGRBHBrnlVN/vDOpjBU3bqCKRovmRb5q9ytkDaE0KsUU7SxZ3tspyLPc7onekASiz
dTchwPN6hdkJ9p5b7elrEhdySzEs5IZ1IrJKEFAXY8IfcQXzm54HRp5m4i63Td6vz8SdEYPKmipf
487XCma3aikBLPTEMH0wxmY01BH8htv2keDI527o4lPR5mdgiNbZChgt+T6ySU65nV3T9DW0pprZ
cS33jM2hxXXSODQCgLJYBCK+pVMAAVHHQyPGQ3+G79Z6hlZhHokf92JewiHQFP6M2deEcIEs3BnU
zI4x3H2B/Ffk8C8W4gfRLrTyMTMfvloOuZ0X4yPD5ozPmPtnv6Z2036aTuqWwQnyE33/kJ+mRRya
UH0HvdHUHXeKR2gIMa8B2g4RLeeVgYWOdpKYFJf/agky9cmAo+7idna1w9J0ufV5kAA70ERgAVa1
e1tQBAgFOnJ4whHMEVU12I/j391FAPQuBf3xlOXX2r89/FtpqoT15Jf2QJ0cE7u5xAQzB2Z2UkbB
AZFCQp8Wh3I4sl2cJFKQ19zcVB/k6T7IRDi78URk3tfkcbwA9bbr4w8q7GJXXInG0rO7Fq1WhAau
PzR2XNPX+mrP3Vhu39lDLoAtYNZSuq863dtsTWOM/UiGby18YS+LR8volxTJx7e+1MkMpakK0pOj
pJif0SkA41w+BrBJTWPiB7PsQdpe2A8eArpDppArGpUnTpoKN0oCWkFKeuR1bZWAh/0EfwgUKZbO
mGYYSFEdAEkAwlXQoKn2LT2bbdpSwaPQmx/9iLOwETOMW2HOGKHzC4hG+juu3mqwdUc/mB11bRmq
k8AzHo01BinabZj04C++4Rz4pANsvbUV+9SUn6ihhGXLh2/+FS0Psu/iwbnlC2GxEytWzAfAv/cw
FCJnfBhwsz38dOr4I/Ij9kQwFHHb1RVIqPjAx7Tz6SGUrEX3pMTtXk6yBZvTGrEzFJFO0LySRadF
ABv2+c4u2WhfYhlPdhePCA53jkSbm71Vo7z2xXtSb2yVhWoQ+2ZwAVHmjtOQrub2BNTiaeIx50Op
oVwL4yL3iNqTpA22J8wBwbIkgfi72rDBJnk/lD5HXaPM+1l2a77/EsO5Rzef6s+44a1SqPsQBk7l
1y2JkRU+d/OKA4L7LA8cHaMeYEOY3o67A5KjdajE06sOCKbiwl2PpVx+PrRu/kaE9+kWixbyGEK0
dL2nFlkgBARF0Xdt9fsbetH4DCLh1QXq12gw2oyB3hkLzvH++ZEAo9hR8BsPKBuup3s9p8IE3x+g
i4enCB4IeJP14MD5JbZvfUG6BLiShFhrSENuU3AYwa9+Yi2k5WZzQgcFECclfqEfoieI6yFfy4Od
LqdqEw3QEF1Lye0s7/XRywwdtxbiL1ZnqPRXMLXbdw6ZTM/ZYUHHL01XvH/bbBB0b5XSkomgsK1k
SBIgZ4ypl7XmjsFcH4QFadyUtv8OzUF/ZAwCC2iLMKyKbUTXjQwDgW6eUMBftMZ1j6XsjcxrGbom
LTVHI08YSxQljv6F/O7szPAR9RT4Ex/kf1a/OB/TDj7Y/dq+sg65ao8QhnO85Pk0Q5fRvycpCZ46
pRXwCRvMdTejdNqp6dm/GLtxf0//dE4LPfyL93l7qwjP2B9kMQqE9WQvMWSAncKfWwG9ik+TzIev
dnf873NKS3v3Eei13mdxS98Km2dVWn4FC2XBEFhxzBYrwAup2eIQ8w7A0ucm8lW7ewwgk3k1sm1n
enSPM5OsjpzG0gMLWW5FQzkbR6G4elrc6JEH2VxxmwyO34fVWf0DhZF/h5+D5og1uzaUKX8GyhGe
3AGCkrf/Or6GXMgOIb3B/DkwRdEuMv9txzg5MVn7q65lgPKBiOB/Ss8CfzwxMYYYTXATl+3RhW8d
IkCTg65X2WjKwzKqdFw4gaSC8rMFRc4+TMZk3li0/II1OjtSBQgaK6LlbyxiFI+qSUk7umw5MUII
VuO3XxqNNFIpGx/I8mGCl1MJFP1m9bt0DjRJkHWdWO1kmTCyel3pEFEJ9v3lJYoIBYhn/5eQlFSd
MW9ilOh7pB82HlQrerP3Iu+lMZ7/I246dExYF01YyUMx3mjnEk488AtWUj34bmAb2iG/NMJR6qFd
jDe/wE/ZaTXwBxe/kyksnYI9oZ0e00SOt7VeMKRx9BbxoULVfcXIBDb7D30cKKqphrQq3QTRnoGs
bg21yAN91zr3132g5iwFT6gWZy/MA5+CfrtR83VirI3tgzOrt4aGTh1tEKIIMSZ8MeoOS/EmmeTW
khWXY+wiinF2EUVp1wpAQ7E2ildRwj7Y/Z/z6l1HEq+t2yIgVaxjJpMxTFMgbSVniytz8XFLaCQ3
+P0vlgiAV4CimeSuA5MQkr1ifFsv9IXY2JvtyNor03PA+J4Q2JdWaKiZk2k4uqbuLycIWqjiwRtI
beDtenWiJGXWLXFfKyw96B95q/OtVZv6TPvW4XJBsCjzAjvwvLsnUssBOEm3xJ2zztn0IJrCUsJz
jj7Sg0QukRPEwjSNkDUX+AlybrbCDnX6JGd/EKpNH6iWp4L//OEZKwSp1kYEy52KCqqgjzPpUs2V
0Jl0kKw5+B/BIXYKvcuzgGXxNMI8nRyRq3NsEKKOcIVkBeCTDQuwr4VaPs0iQ7PvZW59tBPHksBT
zYmvs+mZ+916nuz6n+fpWqEtmUOVKgP0Bpj2Zvi9HI2dRlTsHjZOBQnToEesTLo2z4vaFH/9DFwi
p+OlYWAa7DU9I9O2HUiQrTOCxWB/8LtkrAbv1W9r4x+oD0Yj0/XVgU6gMM12C727+t9IX96g4Ltb
6hmVo4bgwB1wdJnuifJeLvRKdzJamZGz1ELBnAaaSEfCHbF+8cZmlD48Hv2N2vQjHvRHHd7Y/zk1
wN5znyETnGvn2UHk3jUygoyAAZCTr7Krfav/TnzJdL3r2i/lnpIfRHYmcWb9SEK/gn5Sv1S7FujI
SKp3A+9XZo9Wogq2MImof2QEx8XDZVG+lD+8vIHC9XHC9uxTZGk0nLxl3+JUBrUkrmcocFjbo4r0
C7mVCNga61Hw3EIU7wO8GSm7V/dor2O6j0b3gEY21fT79+gtvlSQielfBXKBlfktQrWDzqnpd3sf
S7uT2uQHEF0D8ljrLJ1ic2K4ow0BzEUccI8hGV9XL6+/J5bV1QoxNjZTKhWvBPDJo3y5qOGYnO0L
3Rba9JBoA8q43kSRlbjvtYwKOj7xrY2Fv+cufACT0+vVBF1a13yTvG+oaFcfQXuVznPEJXCnnpgX
TbEUV5NVI02xBywQM/u68TSJcmshR3KNAghm2uUTZn66j0n07IW1JayR7y6ToEFICsRZCqcrkEYg
m8wqt6JT7Aj7Yw2GbIEobHc+ckAW6QuILOJb4U7Cd1GU+KsNhutQoaqm/XWVNOKjNf3Zui7sGWyX
BTl1wbFp8Xw2NRs0vRvPVSOnnrHobUUt96se4JaDcigywtqz8Xjw4nz0j60YPzkwTDPLeK6J3TTv
eDW49ke8XS4WL0D4JMFWcE1p0mBVY/fvz384aprrWx07tHK/gqB33NMI2NTycbEhJTjKynaFYQ6D
YdnRAqyEGooItrzhMXu9QyaYPwJbjlV+jcJm32WYCWai2IyZgL+wBVcSg++1h19M8C5mgLNNP6/0
Mm+D4sC961ZU0aNC557gsqemiGdnZdLfApmih1LLmfr44b2zhKZGbCv1Id3yVNA7vZFPpdK6DWUa
TS8FgxOyaeTL34lgZGuBfY+Ptd02+sq+QB2Om6t2K37vnslUMNUH4vKZ0hgRrZ5hD9sYnI3D9wmX
j3TjSZH3gX848AMpMH4De6BCINR6sT2Hr+y6I/xwt6j6/ZJhAYifSesBYGztki6IXpBDQHcCktCO
BcWXoYLoDpwy4FfN9FsG4wwWM4UP1ZSUmdRrUbCCxOEfCWDpnWXRWClZdeUE8Yk2F8Af4Lf0n89I
/m7IxVdqt50/9brGajU2NXgK7zmIyfCoHXVQIHBGd87P0VvajSU1VuWbI2VFlSOJuygKYp4ogXlg
EIeLwcUaB1QJxh1Mww9bGpwdO6opJ84oUwr577cX/w0Sj27k549Qdy/fXafqg2XRXFpMsC4h1Qhn
ZAjVdzVvchej6T+ezRW2q2N9KLhXrR6kC+mnAke8xxKfP70lhB/5cIdQBMR1OZLxcCMs+9dZl2qq
IWfjlJSAK7212nDdCWA0F5ylSn1iOY/NmT7A+hOiilXmUJACp3BFepfO5zDva3AKVm39vBbCO3ZP
C2VHsjM1Sa/a60pyluweu493dWxyJbWFrhLmJ9OL1C1IhHT3bYnoMYWtwTsdnROWKWjOfLvqSCKz
g39WIqfv22hMujy4O7U7CDihJMmqDOwZ+dQW0iPQODq7UbJM25kcrIFufdNt9HF0aUmF9YalPpnk
zNF0MhOCmujGclt8qFOvb+TdnGH2N6VqxDjyri6jgGU73XXcGu5B35iY+dK6Z9eGnGVcPxL7s2DS
dhAgFelDK9jHOaaZ24Mq3WccLnTAhMxYtjjg+qS3pFofk8Z/WZpYPx0aMkH1yyfMIlMglkElm0Sn
doaF3eus9N/ypCXtGVICfYoJ7COwtpDYzorTM9o424e2w6tEMjBdXcvahMgucj2Gw4p1hgmiUIUi
bGzJqTkG42laKQHIEHYBhg2K5RpQ3suM/PPchopStRFNWf7LlyiP/9l3jkH/rrL8Gi0gaQQMKTtx
Oaaj4Rs2q9VkJHUNaObu+GMe3V0Eou6QO3DZIz9JFhOCX+zrX0MjmBqU7ZKG9LHtNNDOolevPtfb
6Qa7uwf7GCj1BjZD2TOdQc4QlSf+oINzEVKaOrKyat4lHcA+S/gdMZ6ERNlcPH+YCWDkPDlAUyxi
5TdKboNjrj5Ohn1Se4O6kVV8degg120Icf8kYmKhN1V8yOH9OsyHUdGJrAz4iG6eKTfyhKkrudPp
DbOAyg6p8mag6ZC/Vz33j1ibVmWJtnRtFiMMdYJ5YYyxwvuLWuVy0yf+X9FPh7CQEi6EpnTA9Cbd
LuO78nHKMcQ56VBLJ2BPwMEMHWvkcQnH3hJWTu1VwtB7CqZCczCpJplJTsMhNIODibvPFvkw9WnL
28BUefuyXaCAdUoWDVQHkb3IIZeElkxbUPOFX7PDdledg0U6D6+Lh+MRATB48LBqD8ax4LdghjSG
5jqV6wcazdBKRrEkUaPlxET22K7KjdEoeocZ8owqJ3h6vgSNZhu3FBtJgAsF3lvU8P3/vzwxGVhc
mrHlfNj/Tv8vmY9nbTsK4uTtXXdane9rl8Sa3zq/I2BKIVU21Xcs24mSSGqAfkqvzw7SF7dM05eR
rq38138rFutnKLjnBjuAE6DVq0z3/8pTBMTm34gnGRbSLz+LvXTwFmSaD42KSaVrVWzqMor7aXUA
OI/jKJuO7luTSj0SEBBlrWKSJD+PgR4kPOg8BNl8PfwWuC4Xrxt+L6l4/eVnEcuylCdChqYH2EuA
xEzonqAKQeQnfAOyb0u1fBqq7a0epwMVyRH3aFMduHfgCDNsG8wky5jq8tOpREN7fiL8Pbc+Incd
JKXAq9UsUtntU1m+Qup0YGxm5w150cW4QCyxGR7E1WXuQSFHYxQxv3Hc49Rcu4DRfhdYUfOTOcPz
7pMTOKzCyt2GRYgDtk3d5oB/jmjt2o3eIesL0kWDHwF03F5unn1jC44DtQvr8SZrh6ugt0h0nwtW
jCWx8L59GLJFpQ5Nuaktas7DdG9WsINNbBAUQHb5V5dukIB2hIpcmvZQEi3SzzT4gqgaWrSjEqDB
aLUb/YQIxWzASi9btZ57U3x5Jt3qvJ0zSWwHeyARVWLIU/Huz8w744sWF034NOyXXOLM6+rUBkME
P6TZvNohICMsbrgL82g7LMchc6n/HwxAEGx1Fn+FCQ3y3JaR4xEe5p63Cvt4k39VPgsB1p6pPQcA
t22/Iy13ST8H3sjDvo/QrUwWLLsf2YJwWhvIbftBlhBTZQtQriD4/ZjB9U9y3/2NDS5p3IjPQxqS
eM1NkeJBVz3snXjI/XUKtpfp8cO9af76fGnYBfHFybZU0DyhDBAPQKFOivizSPmdivwrBZT0kNSc
PpYJZodep5/s3aZM+6JOTWw1Dcid3vZG6nRFkaorjWw4+v75dF1RMeRwZS0Ipk+8OU5R1NewFmKa
0Se3Hpe0IjjPyGKKHEUuQP1q+qoUSABgLVx2U5q6cmP+9QGISo1o3ycjFIY0FA55ixQqmfGKnCfV
VNwX5s5hp0FdKe6T6/MN0+fqRsRKRQhuA66RomDYh8bzRfCpqTknBge77vmsSDqOdI0JyN+NdC+i
d6/WXknjzl6+eq3tRBJjd5ZcEH4g7d/Cm1beQA8zlZfPDuoU+OVFukbVRzU0hXbs3DR5vONgkxbE
Pzn/0enRzqn6OWkMJSS2xubhhSQxvbJWIEbdJH30x7evKf684jKM9gObuHfTFEH8TaAFKT+gn4sz
5gykijRmbjlTDb1lBiNJ6G/kD7/e0kPGo+Rl24wp4JvGaXkwm/LZxMgdykkJ8KEWJAjmF76OxE7t
7De5mGbDWohvxpmqhDAcqGJECNgARZqwBSZx1K1Xzo9DsaJFTm4frAcgUIBrHakzzmeK7WhzblZ/
gkFhDfMuL7bScQEy50CMH2H7dxr4TQpauVQ8WYMxYfTtNt/G4nEJTJeiOKM0NO5f0hD8ys5aX+Wv
4YHVKXP41fYv+HsKeEgNzToVop4ZZZCw1l+PNsbxNUuih6ORcCIn9PeQ3cbVC0EFSbiY/5226dC+
KmbBzsWPBCG1tQMOU+wQryCHL+5SLXWor9+F6upmFwBUtoX9LuMZyL7kydlNnRpCrG3zmzfORbcI
Z17x08hZ/2w5mNxTbVxhojiOwoW7aGHx1yn+vR+Cp8PT9SayGcEfb1sKovfLRVqmQbdlp5eHf0Ul
jcVaHhk7nL1AUq30oktJKlwCYlWw2E6p5Phh+e4oQvwbqdFJkp48jO71CaFehh/+t+1IoHDUOeNG
gX6K7NK22EoUVndeeKjhJqEtCII7jTmk4xWAZOgdBx/MU/n51sTW6U0pUZeQCkrTqBIB8ePTikml
N8t94CP2V/lIXcZX0SOgjr5Nh7fkH7MDOKUBq8q4h9EiSZvJQhlN3mvPgjWttK5Ly0eq/6XAFJsj
JCNYykW5vn71ayGc6Mz+iht+Wc/jhKvmrZ9Z213/SjPLrWFZG1t8kHlRqTY2Q+MW0exx/8xvMzdN
qmfrsSac2D8XVzJHuu2pGN/2xuHWUWtbxcvczrCSa3E5t36vVoFjnVFZDYW8KXKaJx2XqoVllm7N
pN/aJHrMDGrEeP0iXl52AI0uhFcpcdv4EFK5CsLpzX1FBWGCGdCtwzGsmjFoVvby4LF5YDOZwgKg
Juk1dv1vVddONap2wNF/8KYvPMjunaU+aaW3NiHmJz6MrD7ZdMUoWzeZXkF9LVig0jhGLglNk+Yu
enlbJ2wCzsKOMvZCuujpD2XKHsO2gISmFXCOB7NVgJXeyOyNGzMFm/l1cLIKwj08DVBwtie2nwwi
Vxghd+iuh/f3yCqA0/+F487VhEJnj7+s92n6QW7vdoSrpxaLOkcZ+QqcrBWVBcuCtyCI54Jm5En0
Wv1tuSr6QrjNen9NOGlSAmCNyVRBjJCYw4x+ZcThE0siplj8yZXnnbG4nsC9K7WAIskT1aBKydi6
MYz9EMhALGRAxZrDkZ43VuuLCOwY9etmW8fXf6/2AmAX0EocMSuSkcfUd81Wu/p7kveEVSjBpdAM
seCiQRfdFHEtOGZtp9OlDRY91gMInZ0jzZ9tX6RXV1phhyXQo2NMBYZypb2FGf+nexUj2bzX6jAz
MdIrJzm+oCs8WJzr+pDHg7VcWTXiVcaSvheejsl4FXDtJ5jeS86JueVnYlFEo8taVg+53STbhDSf
R0i3gZFqbn3QPiUfs+OU5ebYOTY1ceteVZeGmNh1e/8YUQDZaAWBPukSRwcSmYYiTeYNspjwHyw/
0vj66rE4R36AvtZBMPZ+ZzZ3m4d+0WJQ65G1h+dAWSytJmeDHmMhPVNlgU/ZMsQ2vefWx4gEpLwC
JoAfmrYwuUmqqyOYWtL7p8yW1Y7etCfgvzw2IWwmtLCkS00biVz9i7IclIdDUGWjOEylweNKe8oZ
BVPA3MfFjawxdEten791pOBfqEcoVLTT/OutVTw9PnLFOd5tAfupFUn2vaWrxO/yqeMmgReGwWC0
RHqGdz2KdGPAgwaq2QYQUujozW2GUep43ogjm7pu5zPJF2g4K4Q16kj8MxSPlJMSv/mdFnDoYHKw
qrk+OoeZGvhybVvfankoc3sVe/9xsRIS5qUFI9iXNIW5boL05a/7C2/uSYfbYPvwClOyzi64woyc
ojd70zPyOqsBsiL6kDrqhzBsgrhvwAbY58ASh4rDL2xufWBHZws49MgLksJSfAriu9RDmSgB5rx+
H+ZyowJTff4MIwx6CbywdAqfH0/+f7xIM2+J6XbvYuSsrya1oxCCt9nLRtWN4YhgB4q+IncttUX1
5inakc9IIWquGONp5BgVWtj25QCCv5+ylqd+GzagTVUA03tqy3Sv56y7hZ95J0TfIC6Lf2KKykoG
XRet/Mjl7ecTdoO3fk/AwvVYc3+01qtlyYw51WxULhsuWMYLP3yro2E9Le9hBTXDpH4TUrwEcA/d
WifupmnEbNw21QfHFHiznZdIktJH0JqA17rL90SIFkutEhwTFsxZUquLtqI5P7Rh45JR+yiu7hJV
aqGin/Ds+GqC992Qi25fWfjmL4tIfPkAeSzrBVJ8wbHw/iaupI0kqsCACmI04cp9pJ2/i8bJxpBR
LvFe+KRBjgfHpAqwk2egVahjul5AgahmuFwKyNR+w1c3wFmegrJvoWy11S3447NSO12P1pGbzHSV
rb0ixN6LJ6yrIcSnXXEgT2Qjz36X85PAxIGAZ9FeLYphXbNWD5Tl5iN0unVuphCmwQPVr62Konfe
c9TvMzbz1igJOawWx1EVqbA1LZe44jQK0iP2K5IcNXcdSo3Nb82eL197AOdcdkhxmrnPxpcIoXyW
NUhDCR3Qh4ix9ibd8Tn40DfD6t9hnQo+TIY0QqLAUYsGOrcoyVNTGfK7EE9OV2tJQaQPRApu0wK7
+chLsFh+lohM9KypOIoFY3iGtwA5cqCc2IneuUHKXQzcCASRkQ55/PtsiMy3zFruGP18Jg2YI/pr
kWYoT9Wo4djJMnqBG2B1szOzWUFQog+I+xd5VxtzzEwEyGQEvZzAJf3hsMXar/92mamPRXok/cc8
SIRZe5vs92qUQZ9eoYqFc4wU04/T9BdN19IvHdtnhGrIpqHKeGqh2eu2VRY6l8DeCFnRcgtHFOlQ
zhEHLKS6ETPQaj6Qmh6F2rdVz1Ta4qosIUwiMOeU86W+rBnjsFJI0rdSR1hRZQ2Uuxi4GX4WKffV
611EIO5UUyH6pdR59xVgBoTpFSbaUSlikvutqAqX4ovHePYUE0SwyVoDELdtlXGkpK8gk3y7RkJf
sZcTit3gHZbvcI/qLfLWDVF4ti1bisPmFsMEeWSFTAMqRoy99A6cWlY9PxemYiXTHC3CcxLjZrFK
UICgy7PgyqVCAtJGTg6MSkaIRagSddE39vqsoJRTzkmtBuXbXlYCKuSdvVweNKZGfpZlwG/sHir1
QYhvlXUrGz/4OwgVuPzBcp8xq0SrP7+Ma06nTpmvVPRj2GhIA0FUXS02qku8AQbBO+Gf6BgMmIfE
6a7pBIsXrTlXC1+ppwgd2Lvh8RCPzaNq8+uO6SULbK/D6pjJkII7eKPX+cwAhsZETnGpMUu2P1Wt
Gw0L7f6rU7lJTP/f4Lsdi6ZUi7dn2IvVdSOu7esKhdo8bnIl3iatxN973p0oOtfzjSATOMHd0OWn
eXLEkgMfBkkpIBtpwsRqLT6F6xVYTu8gHFX19fNNevqcR08knpkiuvjnxI26IwQEfdzUIHlkIRyF
PNkWschviEikzY9lzFiNyv9CsxaIYgO8sYnmg5Zox4flkEWNtQ+6+XkgZfkycK4b2+7JI+AnbJr5
/PqC6FNKCs6ASCKbRDskTJD8ifwt+gTCXe4LKKB3wQwWUIVLczqRfxDRtg6Jjc3WEYIHdrwCcntg
A7EHCZieI8U4gXekfmz1X/Jv3WQmdsyT9nueSi4hYts4kVlU/31aPYPWAPhQ2OBLB6T0Ugwd/9wI
oRHJGJTCZ5EU50F6ioVoCLfqWvEX5LT6dDbgsAirckJvDb5VeN2d9qVWu0M0ZZI52hksO7LJEIri
ebBTeL4Y45Z/lX8DeurrnHTa3j+pQN+EgOyRVwyODytS3e6I/viAB5duiAAZqjXjKp9NDxcgi7eF
TmkvIfaWJuldUHitIDM3qjwsOqIMG6TA6o7cRo1R3FV+MwMk3KZb6tNvcWOrteKpMMpEYMObblHc
PnW5fpb2y52rme2DnNaw3dYkOS7mdRp69aEPMWld+YN+w3yuh7p0WzXzIxTPt2TLzh0UxRJcHlMB
+G1JAD/uBRYOUBSus1nuD8ArSvEXkza08CvWfmrZE5DLB6XyfUL3/D33B6S2Dfni9F7LOblZR4i6
kPFQGVBoIUpHaKeXf/BYKtE5yGB0TtR8Bq7JSBIEC/KhFuH87Q5kCauu/1TKozzI5nDcG6QwK+pb
RyOzriVfrNIJALE/eTXzbBrNNU7ua7uJuu6hTSBz5BJJ3H0Kr3wLw318jvjdObVFX1pVMdPCK2Zt
8F6sLH2p92KAXrBqgAp/m96fdJt8b8f7e2f9Dj4UDxCPcMF+CabvGeITPe4HEi9WjpciuopnvSx6
c46tCUIFp2GzNzfdBCJtz2uF9VHw9YUHSFdH8zT23Z86wXJs3GDcJuq9baI8wRfbNMbM211I1EH6
Fyta3YaX385lVt/bxu5pl1ULAbsDSqHdRd+wkVjJGUIDHTZqw7/Lp0Cjv6gt9Hl0UtIdwkzZMDWU
VHAvVGSEOVWGO5emHwQgbDFiZFp//BMy55v+IVE/EUGAg8wmXKSSoaNeaKmoZ+ubEUPRVO1Xopdk
bb2oKmkEA23velcNpIYGDg2gmY55ileLd9O/Bojj1AKVyhW4s3/4bqulZKjLcQRXKoDptV/U9JSD
mOw9XTvvqNF0Y/GumBmIqWn57WNMFNUX+ITFMbtMWxZ7EPE82DnpewRT+ggDGkgGa3iQg+KE4zxN
JYR556m79ywJl1v9sUOoH12ZcIS4HzCIDAYNu9trxIGMxyM1XhLmdEroJd9Zg1crMJMD5RvrX8OP
oXwzA3twMhXvkNU4X2LNWX7WNhpLYWMvip2wXTa0Y1gVKpHxisC6707U6AQuttLq+fTkqqBVmJ/7
L0uO4gzq/uEEAVfP/MPd3E6w0FSnFivD9pnsQ8PTvi1OAb42d5Znr+i67pGbSOyeUDE686Vu7wTB
dUBbwZFG7qoGX/gfMHGVyGzuN8B0KURf+3seI+skSUQkl3yzoAYW1deFNHcTZRn8qjYx5bD0dwrt
GGz0sOs92LumiOxW02axJKhq54EBH1/pkJJCSkMwhW7LiU9qGs+Rm1Ds4hxy9Ylw6GJ/5L6vxkBI
La6RM79Sn318gUW+xEcWroKxugL6wXpgJMcX6u86z1PSjwpFh98ErMetuxpF4UxemBboaZ2G1FHr
QPxKpCVFP/GL2117YiXcdd6X2SNMbowIxZo4Y+yCUZmcom0kUlON2egRmj6+btyLQ2URvnd3SH3t
N3PaeGvRxO7L98Y6XiZ0ABOVw0IS8oCQQO7W+9EKs3Jp6Kb2BH659pnxgRo9A05d5GbztLSSQofT
SkVraPxdeSxxlyuQ2M44+YQwgpwq5MbY8vZapkv9sPRt8M1X+3tV4kQpPWFdmgXgkhJoJLXMY/2Q
EQ8GJRGJSuylL2o2DzfsQZqbUgETbFCk20gTU3WByXXq3zH+UABOLnJTzGdez0MWCIgHYv5JUnTE
SSf7gyayFKwacern5SSH1ugWsobOPNc28z/qLolN8Qy9nLlW9OhGRUS26iNMFYw6LqH6TLwAx7Io
2ivUC4DMG01wYIOOuOZU3EC5uXhWOuMbKAG1rMLjVt7SWm7N9Hl3nG06sU89Ej/ocGKPJaVid1O/
sgFgnRuLsucBJPzwyzRjZlmLp7b+i8ohWjNzxi13xLI3lnqtA1IW/uRRblxICtpJkrQSOFUm/h9J
wmP+LDAT08jieY11v8z2fIYJ+s1lzGSNWRSj0MlC2jpphM0uuJa3TI85Hp2tUbuOzehvh7il6gjy
fV+c3+7wzna+WcgJYAQ9bOZzOty23lsmCqCgesycWn4KCOjg13lPWd5y+QLK1DPZ9N6lECFdFyTM
+X7l7tXa5su1tp5IsCIM3uAzd6hjCHdLuQCsOt4vRFGtQTmnGOkEQ5LZ5k/7DjxLcflWPOf29Vhw
b1RoKyIbucNagjJXk92eLqApClt67j1TTu05u0vhXEzSHgSaseByspZ5BcgYJCZLSM9RcWSOOGVL
8xatKzOOa/dmN7P3sg/MbZGEPcV9XTy0s/aiNzZBFR+4jGLt4zdTSZdSLR9E7izQmWrBIHuAsitZ
NAmgrRgabQ2C3GtUAPNRRuOjmftBI6t32gdMfi8XTd2YwzPcw2UfGLbj+B7y5RI/qmDQulfxNMnl
jvk88UyeUNH7mbOS8yOQFukZI1qdD9Da7dxKbKi/2Olr9higzmvpttX9eJOTGnjGDMvZb5Pc/RPj
CKjzHrjYsACQt88o/Yz8aOVBsY5oqlG06HLHelAXbBEumhlxpnUVR6UFLlVpYkFpgAolqsro2Nqi
nc7E2SSbgr3vQ0hq4GNbP6cWR3ie4FPAm2rS9lvDTRvi1Z02RBBctFjp3V4kNcWgNIC+HkyFn7dh
2YVnl3yvK1GPt0QLaHAbJTj25shRuVNmHV4vtUqVF/3X4yTOxMohjWWnyB9zVkiZdm04w4CjDmz1
fI7PRyQZJc2uU4uAEWDAp4yYAuz8UIdbSRBXX8urWpU8p9wI4D48j0plrTkzOcRK2xLaixbt/EAw
8nSzY2+r+cmCA3VBz2zwO6DWkIPbUqWBmeMbggjeMNytE/lgj1z9c2JSCqlqSlVjgUTAz8cUM9tC
NEe+761ZiYbQBg+0GpQ+qZwwSL+HTwDIQwEF1gFbV7TlnuWlzVsCzkOFnpXQDo7NE0lstAw6xYGY
RjTP/eKH82Pks152rQW2No6EumZZBs5ZCpFlNbtjPpBqJNLNfB6nfZw4swr5E4QZ4lIO9jb3FU7+
z6og9kjIFE20Ar+K45OAfvYaqWDY7N+SUd7zvurajnb019rb1UhTJYxGCz4hY/qKvX9fpdiuigm0
a/kfai6CRsgVGqX4FarzTSMg+cA+z90K9bUHO0cC0YAAvzS7AKIE+uN9cn1vLc7+oRmLfiS15o5m
YUeQqkxrEDDDC3LpZITLztB77ugqE4fyJZy0dTBUdo7KsJWznxPGJCUj16igZkTmQtNC28NIzBjU
HD8IENKm0zKUlC32aE/dU8sdzFOBR1iAheaM48AGej98hWMBL5Dhi7kbvNQ8gQ1mNxIl+p1MxA==
`pragma protect end_protected
