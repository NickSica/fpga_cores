`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
V82h/mp8FbHcv3//3zVZ5VW10Mue/LSt5dvjsUkiSGtG5WaH8H9Fv7j37k+xy+3/pQvfXcpqBF/k
iaz4/vETUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n4WSOWV3uUjyMD/l4IGcKD1bHONRRplCKgax9lu4YRYlORLHEpckVBvOD9geZHtnlLIjTLNUcuHS
rc4oO2K5x66eEf5+m+hNzaPYWCrVKWQI7/tyX0imMAsD4JQXzU2CP3ATsQoldRyYOQZmggmbIMiB
stLQ3uoRuVc4t0kXI7U=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zgo3FUzRcS1G0FRTCr4C/JBs44dp3dv5CUvkYU2vM2fDyGtu9ekJcjDXnFGi3Qx2X0BV1gEyWxsJ
xqQkFlu/f/1mutspkUjOMtKZNCgPGDHkGfwBEPN/xT22fOBwQJUR+Oj5KSeDWe2U4t5UJ4XXcGMb
ZV9syPFreDWYOTWkkl85cAKcf/WXC6oz+tOUowqV4nSLA1PaSrK4ohf8oaOGNVX+4Ji/w6ViTIJJ
OqmPJQ151npm7Kbt4RW80tp1OmABkNI+o6h4rwtTS1IHzM6bJ1Krrp0V+2aEmmqoZkuKINjX5Pw3
P4Vi6iUmJI0uMpdsCPr3MEC8HH4v95WCnjh0Qg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A45QQ9IEoKpoNXpmniz3AuFZmGAAZIhtA2hP4/pi+Iwurx8nPI4ZkKpYXPnn4DfH42bSsec35aiS
Ve+A8f1Q00bmFgtclspinRe4YgFesk40ftn1mzy6g6sLCNXhUm/IIjCSNk+ie6jVQS7STfOdio+z
cvSm8QQePoJjzlJz/jkNhsD110PhDAevJWb+C5fforY6kT0k7ZmJmE7btahod6wU3o7t2HM6+XGU
DDNZ5E+RLS+IiJYVCOwsdqQFDuRaWwS0k8Mk4UuDiVWtU0+QLFZ/8UGJhy2ZDSYlL/8TrrsWcD/1
Vku2N+fkWCj38RSMWEEe5TmUHSSzP7uBI6QwVQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b+wEsHDGMmVXUM545W/2toIjDItLsHFsIOyFDid8Fv6KhzBePVZlc9t2c1LfdAa6UEpdqcx5kgIr
+oVEglJG3R/fb6dRp2mvlu6+x0AYh7FK0My5t84q7uKZ6EPBxHnDds9FLGQdMDUFv8E10WtGrG31
lkto5q+L5WLAzYgiD3//MgdbP+aqLc/75XWIRhw/PfRn4OqyBU7xSBeoK9TDxBwOscUv0cQ+dauJ
dUQ0W2ZCXwF6cP5c47k76Ikfu69J0/IO+FTLKMkjAB7Wzsyqbpl6RMVdJ/iYscNROh1xxo2k+52w
4l9VnVKN7wTWZdW75B3V/MsNTrKb2I6dBdveDg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyn/owx08GdB/M0CwlYM5XwpK1DLRGgNdNGvCa53fvz5ftb1LM2R7yhWTTXlm8iqXlg1S70wvPmw
WVO2ZNZ0csmDdQcX4HNMiokrI2gpR08Dk8n3nzdOhqyFyh79/eVJzQItyKMQmJZNCvFfww0mtX5K
FbNe2x6ria5jEBEBp3U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J8WwILioFJtk4e6vNsFHYZhWTjvAMbsqHcnvhYKYzsY6fpaoYuWnjTNNNxS6JYZj7bKOFgPjdnBA
rKaGPLghV6UU9fx6UcBVLjNOj95AU3CZPEjWGC/GqjGRPxOkhGtDka91PZuOBRTBqJT8F+5qIgQR
vO7WJHaKezpaUm2zbeC7+ShM5p4Wm9L4dzJ1OuUGZNm39p9FbORAZNzAWa35wpfJ6PPOgATFMi7Z
sN0Hg00oxMFCKSg1bxvN3p4iC3rVT+wV6yuzOecq97B7Fu+tfvP+shqnUhodTpF0WYfGWHeK9ocM
Mg7nt62XJybi4Tm5rgYGMIIM0i67934etK5Aig==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AF8EDKLpUnsf5U27caIfzjHsL1dKCT4FvrlOxjBwD3ZJ9vsXwbWO+EJTOJOFymKnoSSFnuslr7C8
ZCAbkJJLJrLXJwfvC9hiPRksxuYzuxWrtwsjJd+5KWtue3gL5kHClD8Tbo/V+Dnr3gvKzMRNdFRz
i+4p8dC6/32xR0/NITJMYT1uOYu0oBFDHGLR02Wn4PqghcTR3gQMVeL0RsDhJibeNnf4Q0NsKqCF
7OscDpis6r9ZAFao+mdpLGI93rreTlZvJBUPh2RcpqOjL/8IUv0iM922KOCZ6j1LtvD0igXehvHa
5hOx0DDcMjOoejqJiwIqLij0FB13lDBsu+fjWw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 69584)
`pragma protect data_block
BMP9G5RAk03qFRu5UmzfhNOOXDwKJgxZfoTYKz/V88UZr3fa92qF7rXs7/eckNewUxlzrNjvo1zT
4g5opuY+vW3a88R8mQc1x7I6d4Naytx5g71mwuvh6KS0mH/P0lIxy1WMoPsjrEIkecYZzfPCQOv0
SL9V2E1j4mMz6Vv/fTMBhGTzEqS5xhwamjThXm4h9pjgnOMd4ZqvWGM5Q92hJLFf1Nmgb6S9adCU
/l93FEVvcFv78yxFQxmjn9ZR5FbJIh0eerO0au5K4S03fLil6DTkogjiJ5zmq83u3ynBOiFa16li
tyeg8HT5XOa1lU7vZZVOsNoiZgZTb2EHSnsIHXr9hsuIqB7hsHAVPFJIJHB+ARmqqQFyAVHK3wv0
uWoAzCPNJ994dtcyYXoj2MwR+g5Zr5wlJWD4ZkISun7wWyunvP4jS0JpKctABidb64ffiU24HKPC
caTeZl6SgfkT6oCSnR8Ifx7iuBgZkw0wCiDgGp9gGMd5zAfvvB73k6bA+TpLZjEyTw4y6q+rGwDp
gMs/EkhpBwE68prtkOIllsRJKdJ1LcI4+5LSzy3FBma4q3Su1T6K5uk3t16TyaJCEZra2hJejp2O
IoD2l/25hITleev4175fcKX6NmYsIGtlgc8lLNK7901uGSqFFNx4Gx3iOl6OmxxsxQGAeD43y4c+
hLKhw+XjxfYalQ10UKnAKllu0Kcs0n9eDizCXHcWZ7gFHv0QSR+tIcsIzYAyxDbAtKXpwcGsy1wp
82lau0yG6FoVLCglW85Ohp1F4mIcQsHnaoHJae2dpujV67iWoxg3wMlrn93nWfGlp0Tfc70S3fqM
g5CjMKY47J6ScAhwbFHqqPM6jepiqF8XIVj/Th6e2XJKrrko5JUkrMS3D7/q6y5s2R8OFyaK20P1
oqaNd/6PCK6UPKrVCLhxgJtPUdNk+vdP5IrcHqsO6+auIaBsSLi2LKq0OSo7gM/IFyZkXeL+KADx
xky9G+0z1Fb0gLn3yB3i5SCFD2rZTsBrW1kgkrwWsvgFKjGReDe2uQWZrV5YBOkFcs0NblfJJZWJ
J2XYwX11/8EnsLhPjjBwpuZ61XsVJUrKf+XeJWjKHy+V4+UhSXj7LMs0GuMFF6TfEKOkZuXxnr4O
+INsGhI7Rbp4b9mElrK4GEFjwmoMgVa1q1y71+Tvi2FfGJimbWy4A2ATEDWttPJwqKgOqZnvzYCy
Cq8U/AaCPlfqohJ1j5gRaRHUPwv/IVkJ7JeDVUP257lJj8z+OgYD/h0rwqM276hDgAofm+DR6JWG
6u2qhdOMInHq/Wvc+7fb5MDf1PsT72zZsw6Zg8nEAX4JtDT428kSurojntSPUiKSHN1M+IFVRS1p
Ykar4zAGfaeR9NfFCJQ+h31J/EfDj5+DqzVSDACP8fr3n+spopk8QWSsr/AXjM3ueifcXYTxK2nQ
YjcQ8jtX4cR/SsJSUMscEu+SzzTzJzNDJA2t6eH8mfiIcHDncZk5DNay3YWsolUMpJOtWpV/d102
vi/xCSJD3kFMLyjvrfdTeZB6NB971loJS+8U/Cwo9xOtE2ugD+aLhBWosdICtpwuLMCr//cJquM2
jS/ZXMyxjV8vPgkKxkFhBtBjWteHj2gn+rrOnEiek8MnK3sxbEpo3SkmyPpcH9H2RbtwGyiUJjnz
Gwou6pN94up7DDSNB2Z+Dq+qwhp3OI4LefAArN2spMpauLWDOWpjfoxAR8x3m3fkvkCwT7FiW7C4
fDI6TuDqYPHxFsSCWjzLqm2qHBfJKGd2Kz5BA8YHLMks3Ro/HE6DV7Gf7L0FEedjKR0rDtcCddVt
xdY79WEpxkqYvogJlGvXxBtVAQVSMcdywSVgswa66fDK7Pzh9wUVo3xrUbX0L+R9HlYaCVOPsDJo
vdtC4PCVzjkh8djG6n0niFtFR49QZSHdw4DtlWjd0CK7nVgJhDf+j4THFHCYAfYibCaK/qP6SFoV
o0sGjqKMpte3U0BpWsNfYWvNZI1ZNbeDIoyIaTtDf136K4O+zMXsKNTKSgRcdVQnPHvKmjVsFZSt
JkJjXorgiamNzuA//Ocai6l6m36USqoHHqDjHKp7bgapwnvzT3eQqzgnWPPrxotzjeZFd7kHd0IS
j6c8xMVvu4CBYhnkk6+Q1zpQOcb4yTM2ahOEXyRCjUNklj08QVDJA16+36IAS7xFHpwZWOkh64Uc
CKT+Gz0CIGt4RikCWWaEWBIw2jDO8KMulzOfzAjG6PukvvqtIjU7ZqhWm/D97Xif4342mZMG+On1
lPCSkT8RUymv8dkIPWfnSTnJaTxkC039ycsRltV/8L9k2wEREIVCd/hKaEgaK1y78i2cl7a3u81a
0Y5/kVMyvw2G+pPM7aMHpuZOH8s/kUWrKCzdjREcSnU4qHxKtMbm9TsGsX/6WGNUoYidViIrHzti
PjCIbBeeqWJzk4YMObNNLa4raX+aYq6NIWo2K6hWTW8+FlqGxc4Otxk/rKH9DhSOMHcmCnVgynXy
kOTQ/fEkM9fO9ju/7OJgn+HNMki7XE9fLBNDCjZNCALQOH7yibdA1F0MEWaKmDQKAT205jenjzci
3ix1tfa1O4cN10qoa1TDQa2niNfMR8MbD7YXGDBuLEedI7jO9UP2M84k49whY+BDoVzlrZFl1s1u
/qERh7AzU1ZrfU/bNMSHAqypEz2DmLANaEwbJe7foQq7I7Kh2A7Rv4vRKyWgX+Xg8TYPHQlsJMSY
eMi7FilXiI8gG5sLkNtXGRuQSpnpHVHpjveKdmE77P7LHmlbZSMN4kiu3DxMHRQTfDePyS1BbPks
W4kQyJbps2SAhm865moZJD9cej0UtQJLSjmHPi6KoxCKYMMksXKdCtrkzGG3vgbC2rqEw+/G7HkY
G4F3gMlRjZX0AxRDFelOM8LIZTOdqFzEk98bAFXE855JqZ4qaHRHBQzInEm6czZw3eR4go4BCtmD
hfBRDdx7NCT+qjA2m0jHUn3CSBnEayj/jX+pj6rKI1oe3W3oQ+1Cj6Ws+XsxonQXPpSEjXx+ochq
mq1AyLVdNtAKr9/NtpAp8ogR1uoFPAKtE8M++kt7EYl/dpRJzW+qbd4iliDCWIPl2mBm6dBquS9H
q7FwKkgX4P+nbg/BeE9sppEbxeZpiKlNU3a9Ft6Gq8CEdlLXFdrxDJSTMlohuyfQLyG2keYVQAeU
7/bAK0bikGLIh1B/RKIfOw3aFx+ypTfkzBW2s4LOfn7cWMINze6DilQZ7YUnMYa5q+QxGOmL0SzG
jJHvBEQX7OJ7DMpyaGAGzpZPY3JA5m9S4wfUdwUVg7YB3YM3b6WcRKgAot5cvPgl1tbWtiH3TzRC
PwuD7G+TxazEE2N9MtV4qvXRfbhbMUhDKT7KRgDOJakvU1Nldq20HNO2YBBAbOzbOhPyoAKaX9/H
JRuiWkokIi0ZJouAHWGPLBv3/xdo2R6ZFpD7NBnfoXECCpKVoqwRjrb86h1Vo+BY3UDyJT7QZ0bL
SF7xVNPLfj6RIvPbiORk5uGjz01hCMiXoPpW8IfwBe6bHAoJAnohFHjfwIMj9zOdvhqaZJTS1faK
PN99CBstVtHrQmy22pOXJLjw3oZbFP8jlytlful3kOcQrVD7vwDzMIaKJOjdslv5FS0ar/dWLzX5
FdyJg2gvg1MCX8NAXrIF/9LMf1++aoo13tLEscyzo23bBJ5Tm23w2rOBZTpmc609jQxLcbJGChI5
auBDhkILdPyXhJ/8uKEm25h5ziLbVugoiR8A1eXkn+xYpt9UVT9d3UKMwaTQh3OLm9aP6FkGuXei
KNgjkYga79u24yKmHG+c00C8u9EvVUAQcZGhGCgdLQRkgmb447XuCBLcXsBqv9Vrk4QAoBUx8JiG
mVenEaGl84+rX5p4mCnW1aZ0Mg5HoBaz9hK1Wh42C71gVYd2exhKaIha129XhFVheAQ1m4fJqjhn
E+OZd2CXlQwvN/SEStYubr/SqUmQLnifFJGC8S7Yw1puZ9ikHubV4pQzmPMvMWRg4+EZs/O0Nq3A
oZVAL5S/7KPYh2N8O7KmQDQW3oJuJyDieLVuM6IOHBPRWCi7TdFqT8UGAVycOXhNcBX6uuQknBqW
Kd8UKZQPhisQUmNhEvoGdpUdT57lhs8S0P2NfyrszpzlsQj0R/nhzNmnF2b0fhDuySBj8125VD/w
icJHY/F9WDwV4QIQA7pnnV7P0lNh4wCIuZwnZ8QswgXZpXT9FaFCaF4KfJIga5VrS7vxqEqdQ8SN
erVR4E59NcyYGtYrQOoSFAfdVThajPxjV8IDbdF+svECMm+zTuQQnTTOKOynSKe0h9LIOVG78nuv
yv8YUaBKWR8YZZqFhCD95oAUtbMC0bNknORnwmHeD/6uyrHO7B1fleK5mTNK8HaQoPP3ipGjXD+8
eQyQZG3Oo62Kx3vcFGODEahetz2DddWXV/OoOlH2jTMQUTOvvdFVViWzxFF+1V+VOl9AOhzbZZDd
mKIGSym6Vwf4uYnw9ieEnM0vedqMwJC6np4c7i5H9/5reU/O0TBK6ctS9ry4roBqMPL+krqXLwRG
EZhaDzKTLFDL8yf6eIEosfwUJg5cKFbViH66i0S7IiLHJq2kVtDcVq4R5qHUtoymYmAMEs38hx4N
9hpFQ2uphvaVGfchJCgWfUMiEsNpVj5FYRYhjCPJSWmD90NLzkPJ+uQCYWyt9ey+h36Xej64TJgV
FfAAhvciRB/C0GyNm0l1LTqSXDFRuuNiZ9+xERLSpyMWAeRS6hfKXGtJ0PEDj1Bks8wbFdmsqYmW
KSWMe+woEd/7UKvYA3ClU3tBDSadwsaR/POIOXPQL8xbmbraNMOlLVZmK3amRVdjHEs8U2vSesyb
4Bx709raPjAYDX8NPmW6a5njd7KRDoPIKBbeKkS9x/WUGP8TDrSBlvNGFTqlCDpIh/VJ4e4Mquct
pY3B+iA6XVq8zUhimSenfe/iqrBWlF7Bov+i2SmEDbMi3Uoy+lN/KpKG/CgY7hgBGdM4n2NcSXwv
7T1S7UQpuYwkEeFeDuFGkUiwOhvhEpGJompQCfwS9kOM+zwth1EaD1H4ytpZvOj7Ia8xUBFe5jLB
FM9VZy+xZ1NYY/qPr+5mr56wp80W/I9nf7kZPcru9EpbzB2rP09X36R/nRTmPptjsoHebqEZTZ8+
YOtkJtaCWUMshVGu/NAL5+J81I0oGnlusHj+eclXrGQajEUO/QpyAmGysa6i7C8vVKUcN6dY5qOW
MKSpePNv0Bt2xQ4PGhjzBjuryQIBGS6sQYv8OJOBu7dX4BPCf47wV2YLUNNuWDlYugqZG013dOJV
JAaJ7ezoYFBIwcP1KQNSnEvSv7PKDzpDidao2Gg4WVCLtghcVuiVCWgHLJqaiKnyUF7CIvV0ImuF
QkWQeNAoX/bLjqhlObDR6rurtTMZ5usLhozMZPDd/VseIoyCf/CI8Tme7BkX61eYO78vJmO/tsKC
J7YpbkMqHTlizyNJoElwnO99U1ktSpJx6bJJu20KVAHXmOLQu47phhPqY9oI4YScggq2WDGVS63q
O18fv2y1eWcrLEyDfGJGIR1juMx5lpiAyvLW0d4rhxO3O0ddI/BA0ttmkmAbc11qdkZnWLWI4HKw
1cS/v4ST/fDCvsPestuIacEzCEqT9njGBIAIVK6L6mNtdvN4qZ+EijHKwGN0thDFpYIxNouRraTD
JAM8fvwuf83lf7o9/ZdoAwFbC0QiA23cSpqv7M5ALwiYgQC6DmM/bpYphJbZ4FrYm+26cKmH9tcf
unaHBjnKNJ3lb1GYVwhJAtgjF6AC8Yf4ZxxjyLMzIwus9eY1qIlI3OTBSU3zaUcquZSRjjkNz7tO
7wGpuPaoQJ9GS5GLWtsaaplMi7siYByVvfRf/nyngX/7o6fXBA41Mn+3IsVcBs8zvdaP8l1B5/54
j+il6eT7uKB4UFLHSM+61Jt6IcU0qNiEb/AA+WKtFGr267RFuqODjC3TWgURUUubV2lk/16efTfe
hgXYazlpZXdJv4TvR2QM7sVnwliJz5RbIA45gMg8/LZPQ5XrrbDhZfGm39q1JfpdgKa6BNwvPQG9
3dLAwAXXwUXJhc5bwO9BUk+izJFYdPiD2CIHi8ABIdNMANksotfqpE8ti1brA3JoJ4r2WcwC4u2j
NOt8m/duSjdmFZB6yF1KDBOcqO6XzY1QS4ybkwM7spbkzCjO+ogFcP4HC3KyFYcDm/NDgaCMfwhV
nNksyl+ogdqDV5tXV96MaXJ8eldsNQsO7l+zHwWh627mB/JnZia+MSJZ0yJP/34FJPC+1gpeSK+m
1673qeROIc6s3S4kwBs6k+V+gpMGW/x8Hqmv26zFrfw1YNPclwfP4vN/3YS6Ir56ZtNIpo1BHI5H
SpOKgnfG/T2VSvTmplHTp9AplpbE43zeY0hr8s3ntosHPe04PPGk9uw5Dh8Q4yu00bVrt54w74On
JDE710mK8bDpXHWoqPUrm9nT341GD0DZXsa941LB+BIGdYcbcg+dLS3Sn5uZfoA4hP6po6rijGE8
zd76PilymtKBQfdn/3v3uZf8Ekzx91rU9eKMJFzBpC6VSHTkiw3ZR98Y0e3iz1XplelCxjkZLFG4
r7m1KvuDxzGRGBrOoopInZqhQrAcVbo/64X6ebnX/g4meiNmGwqaywUuHbbthoPZG6Ivzv3y0qed
fzfhkXvpC042cPEZOx8Awf6dm4DmYRdZy5cVmlp9u3ACfMFZ/rJxAmiGkszWYEMEv/aQxTx+CYor
0sIQ6j3NLKBGRPf8S8HuKLaNAjiokShC8duvcDxMKvLIrjBv7svg7Qp0kcGKDoStcWrRRuMm5mH4
G2Vc3qP7WWFxv7OcG4yobozJgC0OJ67x8yWh+11/+f1ohOmf1FkEsVI60p46oDe8Vb9p6ahouZPH
TBZ6KTpGNFt1MMNLc/S1GLjrblVmLLyeeO07UI6ckWbLkgK6X2yKC15i2CarJxhmiOJDo2dnyK6R
c9F5UwomlDIXPTT5dvAkjqOd53Bn7dbcUW8DQ3Wovkgx0O83sHENQy9EzIlFFaMz99/19nAxuiXC
QKBhKGVHNmlVqT0/1CYYEMcSVdDvHa0r/yVv6BK2UxDWR/hKROzQmT8bO4GoLyBJSpt4BUmMG2aS
+TyT8Sewvge9bZ2JaIFgY5xlzb2qB2X8kwIV+gdvL9UpXJhzl2JaFwSCeJnO5C0qfkcUSLUogyj+
7DAJ7rHl7NCB2Oa54+3h34DphHj0l46rWYTs/1r3r+1etUZSo3zWy+jQTxbdoFSakDSdrLN7RWCU
OH2+TkfPfLmBl4v8EqnZeHeyMOTKV++k2bkmLL5OaESN0T9+tn5OOmqSIhXW2gO0EjrhBYXYv6aN
4ZuoxAQY8b8WZoX/wNvCdWYQLB20UmamcPcSaceLqXplz04Zmd9sR/d6rVt+PP8FZAud04bpcr/w
59yXzIDI+6k9zLMzcP5f3j7z8nImVSIu8Jto96J4ym3OYO3S5Oaep002t1dkNjCy8MU1WLSW2F/y
a5gV1Uw29iTI/+809BmGUJJSHYkQd+MzvXlhH+3Og12OS2iBZELl/NlAuNJ7XzMDrQodVJsImDOI
tcubQbH+MmQKJu/VVjiqiNp9Cf5yU7Iw8Qx7wcQQ7085h+hBpvX45mKmmGxznuKuYMHNhkYEdImf
BdNmJe8KDSdlk2LhC0/NUkqUHIhjHm/ONrqbTtQaDjzW36h52V8KvY91PeKtAjmryYPZ0qmNqcIy
fpq2ROZ1QHcc3LYqJcQ/g4t864rj1BOhHHeqJeGV+D7DFVV3CR3y80fu0rd9u84B3vNWehjXp02O
5agnuyp9EXkHC0ufacL5GvkXqvwz+QU3jQ077/phqki969vfhetx8P2dQVZ8Fn50AZqPbdXSIxXe
C87h6YFEDcdwQy4kyYtRTDLyo2r1jtjfad52jHvxvsLTA6ACPd2s4Y3mjsoWA+GYxv8yF89alZ43
zvgFE+9lOkJYO0Y0lKnaFqHiK5iYDuLekr7Sg9gLdeCWX7deCpu+sZqs7wWTcCE+c8HUe92s1lGO
8w+MOcYETXnpyGuCxZWocfq1I4yFkOSaVXh9crM6Tf9uFFkOlWAC4/9D4uOjm1TtIFOVQbCp5BUh
QdMUbSJ9PNgqUcC3N9Vzp/rVizDsrq6yjtummp3Q9K5uJnfmZoTj6OF5K33P/7BP4jcGqKjmMagf
Xe6je0IFhrIaKm7RcDg7BSG+s+s+d2GzQgbfi44C3mfQn6mkhhOFD2x7JIGlX7orKcIOyNgJpLhv
oz9wfSdBtsBhV298ky1A8YZr0KE0Tcp6jFx8u9WXn4cZtkyMfzIvEyg7jAL7TtkoKGhntkd5aJie
tt1/S4C0rGT3fJlofdlYzLOYVI9yfdQL3CVjVIJxS1/zJjXwgs0jUNKNdqbE9oDXYVyGFYAyEvfE
gL274j8UQORc31vP8U3WMF69hUZzWmmvG4z3RjxvIAmRjAgrzKw6AIW+xz3+X6gGsePnoe8m89QF
VyPwXbstCNyCUgOB5AGpvT/roMg4PYhyoMsk9ybUCBeYYROFmlP/+fcKw1IGaqQLHExHbCdjHLeb
LhlUpCi75JEjQaLAJz3YyzWRfv2GeGmK5+Ahk/S9UQ4BgJsXcJcDWZ3uDixA/vSLoIWxiYXVKiX3
1sbTe/NCxTwxhmXDpceX4TVd1vIWgIuiR5WXIVBtcvHQzmsD13PjolaWvi9G/2sH8U370Ioh9i+8
YhYvKUa5y9efxRhz6c9x/NdbT5/Theng0mD73DTHwbvYDY3wQeth0sA45bT+7FZog+WYuUOeqU7d
4HGpb7WSs60xZexxjHjsg2zsNPwxt8imnJ3jUH0ISnZOgf1rkpY5GQY0NKAwjyfb/mvuFQj8/0kN
V0EZTHuB50MjK4xxSFbPQLBjDYK/UiEQxZxihaSebd3oswqjt2JrjME6JVCHpRThWVt8ObeU9ZFg
LTC8D+uKVR/p0kpZH8bli7SetqFAPog4dp7cC7Qst665xT9C2h/cY8D1odUUNUeZ+FNcnnmSGWyL
9linX3PZoksQhcZ8w4FHjykTIVbcZ6GSXEU/Kn7ckDjX8bFa5uMMiT6yTWg+M2Gp9GbeJLZw87jh
GD5vd9QlhO0s/fO9h9KO0QoFEE3CTsPdlkidZ4O8s83cRekRflYD64VwMkjQYt++4RFgURQ3MHKw
Qu482mATuJYKImCPMjnbJ8YIeBThwu/LU+GIKd+4XES6QV+hoBFNmFKRMGz6ek3GjKF1pMMCQt5t
HYXlo+KhQoPMTMJtYuQOLwnohzvrOzi1h479VQ9/IB8kBgfokEMUb0ZTV7a5feE4EXM3Autzaecs
lEmOSduZRKMDEzwYMgQfwNwAdtfPDmiRoX1WXpb+Gfn/moC+AN4HNZ6U5OZSmhCUazMZ4GYjO3hN
RhCkHDZGRnsbx/u7kRZdIKz2PjT1g599GQQQu1LHYUADkEg07fM8XqixcMcBXsW70Xu7Y5vLwqHH
kEqyGIChXSVPCVGn6hkIyIquHX/2PhWDYW6/7sMAYsXiyY/jIfUlIi3ZIcd5hEcFNsMXm62D+x6I
4v5erwdtlP+yEvKVwYYyvbOBs6aCFZodCkt1Ks834cqVEJHkxd/dtslJp22lHoUxyVlAiB8Tx4Bq
uFzV3+Nk2WlnNVMie4zx/w1O9HxxKUcw1OXhyiVyLI6OKyBA8GdTOFi/8xHEilIsx0jQ8VuprEkV
WC8cXBbxytk+4MB5WcPUNUOZ/sF1804MbhLcLD0PfSHk/5dxgSekBRUXQjapOKleyHNlVVxtHh4s
zDoijX/bfBBrt+cFDQSk2qypfB3sqP37uAzaJlCu9DmyAhK49FDfYfluyIykF0m8QpcQZ09JRha9
PqvWjaNN8WCXZX3h0R7UJjQy1fpEaEyasgrAF6TNx/PHXN/7CWOp0P+70DsRyuQOJbaknl+YYKD8
rBdE4I9PzSnPjzKEPmqvNkGiZVe2VhAvUMkyxURWh4awZ/g8EzLQFbq9Tg+6hnwbo4dW2jl226r1
X0k9SupwW4ilx3vZ97ttxTghiVGT+Hu9LjwogSBAefhM4jXMKWBvj8GYQ4F/iGu1w/RD2Uy97Xls
z0h8ooiWFbW7XGheAod5EvVw6P2pN5IMTa9TMxRzEdD6zDEfog1qc6eiNElpVdPQ6yPAEecjCO33
3DFH+B2/LjF+IG4/gOToKdlrTMvlClYcpcVktao3nnxyKU+/d/yqkSn21T1QZKjjKFKQNswqkgHr
mheUgyDb3u8nRx++y79Hp3iQVcoBKN+WozlqsPLf70H8bS39iOJXrSFhciuWhoGO4VTstdl9ezyG
p/ueN+uoOaKgSMJGEle779QeoD+tAgw8P/x3ZizDb8Os/nE2Vimuj+CO2yu1XDwIINco98a0D+/8
BIAuS2hPSLWS2PZKAVgzsUUw4tcrRHWwZMGWQ2sFPNyn6QZ70UvxNaPa5vo9MN3zarpjxnuQtF9J
Weqr6dozIX94Ze4mWcI2v1fFRLe7ahmA8rW9mHTRQWurDfNO1gYafIfJXSr38OFaTJMhR2rtzFhe
zjgIELMyD/TL7n3CEtF28c92RTOQTK5bhzWysoLNmrkhZewHBa7Ax8kTKYcEvRuR8wlGl5mQlos/
nIcCpmM5L2yQ1cos0Y2ZDiI8h3QKJNiHBu2dz392GASPxNOz5NPAk3WOogNlFdwrKGfXlin5Le4X
5ye4AdBil4gbiD/b6qt16/XDMZc+erPtTmals/3+0bdh7z9otdelc/tAdJCMhyFvSV8Ffb+pQ2Sy
RBYPqgRZxlmXrgyIihuRXWH+0XR09uXSnGe2oVQaW6j0kD9MQdiqyTiKl/fl24/Q7QEyDlPnp86l
BS5m8NKiC0u2hDKKeh+Dl51ksdHZXgzvauz/4qNh8CJHlDSEvM/oCn+5HJpnQz5eWspIY5rVcYAF
q0nM9l6F7SESd0eFvkh/rP02rR0jbeI/dAW9t1CvbahVJz1Rr7qWgx3PJFQqL52tPNP0zseqQfta
BwZhN2drtWTnMoAetOf2/MdRt17zyIhqiDoL7cOjtlw8D3jB6g2RALeMMyPv2qdq/d54nNxOLhuv
CRrbBcsUMQjRhxjehjqe882ghmcndNoxOuyGBM46SDMiCK03kmnQCyX0f5pb96yXlQtMqbB1q82c
ACtz7XQvy92FYIf8gp7t2ZM8uWpavkwfv87vtcdvFFfbqoBQ9sTw4N0jf6gzzdx2YPvCnGrXnM3F
cDn0n8wy5WRTSL8WcxVyecYmtL6EDwcreBsCLIcQEUkk51EKD21ai5OKqj4ueD6sbv0RQQ2XQ/DS
Un9xxdMjuTG+5sPBlObWAfIFAV9K15F9FWtqqtjnv69H95NQ8Wn9djUwdx6BQsV0F8nFqOEGTtGO
r3dCP/ucJkvhsl60QnFpTTo3Cd67aK6lKtJH5auuNXE3Gt1gU34/ajZ1nOPiDq5LgOQTc9tL1hgP
kYsG5lwI9OyzsUNTtryf50ESu/KP//Ja3rIcXJfELClNDLDRn0/6rzeGbLD2bXtQa1Qs8Rp5vblX
Ziuck5s0dvBm/WHvyzuBd3yFxmmrLNCK99thy17KhB1RC+k3ekGbsx7F2zCn9giZlxsJ2USP/6te
nTS1YMdwA5L34la5zU3zjjze2TB/eGbYIdQmOAAPl+ZJmblhlaooRRYvD6xkwmQ1jCqkQnfOV3dL
ZYw4ICWuTsbtob2KqRme7rUUT7A43eLUeib+Z2DNZI3S/0IV2NTRgYKivi+4+RD6nm8cB3McU97n
qOZoZ8nnOha1GmOm8eN6Tqfjp0bOx5/FA7EJjdXAQKoqGkFiB6hSW58EEb7G9XzYzKHsiwIswEZR
dMuPz9XQCVflneZ96d6im3Z/K61WsP0rf8Cyx+iFMr5eQuvu1/0kOJabVFAraoAVtk+xBgr9VZ/+
NE2assEIcu0JNb5RWmCuVU5TPaB2dKbRb1tl9WW1hmqjMRpKhAw+enE9iBZewgALk4DS7zUMtMn3
rGcpafueXajlDJheJzwoze+AxP+VuPEm10pv6kzwqMTTP7iho3uKQnmqMWW+onhw6z/EPK+pl4ns
zccXOj4dQrpwG8kRr3FW/BiPX3kemD3oxDxoTeaF42FTq2sK0012kzGq5LiG1VPoNypUEm2BvxMq
5KJfyJDdf/1NhZdlipOKoC64RfyjZddljcZzU56bVypgftnTZSdafSti9x77KNRXoY7RO2p0Ki3R
enXC6tXwnxIdZ8w7Eqxun8dbE0uU0RtTD/7e17gWcB1pWO4ODSSlKr2QWkKOq3Y/TLYBMIvxdTKk
u1HRoSDCUHGtroebo1HavJkkjHt0V8MNbYS/K7pG5+Rr0nB64z60rpMDGf8Vg5PFHILAl0nNfT21
7DCfSo/RIOpvKG1sIi4ZHiUhn1PXE3hGEgD40LpN0n5B1Y/PGWrzxlnWNW03U81T85jk4sHloayU
2rCdT7O8JIJwswvhzxOozhRaTxEfRIgWXg1kY8FVFRbRZYDx2v+1N5FUCHW2ieYrTgDP8IZeqAii
7hEpH5qG2CRTptuisX5t0EKHjhsvwq1nmNS6fCbit/uUVQubmgT8rHQtPhMtKVHgO5i2VYB0bgbX
1Fw+JKKMKzl1erbKFNIo7V+3z/q3Rd9EROE0/75iaG5XfNFT9M7y0h3ULo6dF8eb66kmJMEUrQNF
dxhZOABQ6QRWAWDf9R3KXqnBiSFJkOiX5xjDw28NDZNAhC3j4QQ1EIUSGznrl4JdMJL+S35Dl5lc
vyfoIMieoiyEfc4cdlUOWJI9wK/q35fl9B1zEAcALPwfkbankmGU6YM6dnMhDQTn5fuMNukNyMIg
WFKNVo8M8eQNsTUsg7AXpTx3JDYcu7DurVqUAjD+9vI3UMnMYEhMfx2Pal+Y5GZfZCa79xYHW13e
PJksq4yOMvVFh4W2tjBzhUe8qCBXTw+l853q+AGqMPQdPNWwpgA1WwBtYkLSJJPq6Zws7pwp8Fvz
U8kmHDpG5/MfAxA50J1KYWUMYI3/2JfnObev78UWXQVcbAVLza++CaN8x1JshqSqb2bWJzzW3Ebu
I3vGmamyNedIgewCCwrFirml48kiiUtaJB0VeMq8uENxABUVJFk4czqH6VlZE0A2i2ElUFgAFNEd
prdD6csVvyB3Ktb1iiyrcUUUdp/r0wpJez9EuPWFafHqxij1p7837ZLkpTEuHyCywbk5TRqDif2b
4a0UaSZBFlGN5kp8dnAU+jk7/4WXe/9Q8WCfCEWnunU11AYtYP95LzgWzQGqGXLjzvFzeN4AJ/Pm
AOZyMNN9Kcspyt8/n9k3s84AEIADv6j8FXfEYLEBqc1DF5oxQUnU2pj6iuJXWjnwG8tH7TD6/gbB
nbBOuU9zsZhfz6DujnwPuuv2d8/Ar01blT8Xc8KqIiftz3mLWpauagX6abtCkp/xaN/ZLif6q1nD
QnO8DpekBFJLUGmf8wRT6J/zZPoMmVPHB8jWezDnoXCM6K85CTA185huBADDvY7TKTZH1xtWuKxa
FWH3c9IGFRyQ8Dm8Q8QswCB+945WnR8XXDEdf8VRwM3lRYYoLO204n0kxtewcI6t1y3jHB8/UVZt
1q+27na+K2mk4wkNxTIE/VzCpOc4IG95Pt/hNRzjrX2eAjz9HBAhRn1gcCU0FzJu2yDrrSTi0c9Q
8sMyVjBKSKE7HMMj3CEQJxI+/FQu1akg2ilzVjytRlpQFaRkVhmJe7IBrKXsrwEb60hQxktgbc9a
9njJs9xYzw7LhGaaWiky0KAIsd/0zmZBTK0wIkux438ehUjiBtLaWg8Bnb4VaTmTNhiPmB5455gH
RQUy6Uj3TM/kbFgje7699/cEqzCo7Ijs1pJ9mMXaDcSyIYXtfT1Xv2kDFJ6E7sPpIxQssx1vjsIS
jgVs0YQ+q9EmUWXA8HRr+klpjfD61p7h1DJr0fXHblow/IypIs2cbZu9G2D7ArpWx0zIebXhkdRQ
SoRrbDlkM3XzCkRWfnCvGP1onwf7wzSToXgceVDBRbo8q7pGCJV9qxNEhYgKNo1yCvVrckSNALMI
r7Ujdm1xB/EOp/7BZAvOISNODhAaKmCCMaRRDfC864l+ojXndmFurt+Nh0ZzvMXJtb1xPeBjQ4Td
2obXP0nPX2xaxF6oJGYXNspgH/pSRf47ebqwJNasvAcePioweLC+uwxc2q1iFxuKaDLHilGYLl+S
+Dm/7upsWNwyOugBuHQFaE8KKRxueT8X4UiaTm8I8QYPtCw5O1UIdJsCtUi3vHzorPISDfJQ8fvf
1fhcNFUp1xg9DeD2HVMKFVzSISnUuoXVYgUZP57Wie72dIJw6cmVX33axQ1RrBZO5GfgpfSq9F8H
7KczUoVJerRFCmS+ruIGp5Qkg1NAHuB+jLXj/mp2fiWJ1CNpooq0Ai7XKToIoW4vn0MtebOeKamX
tBHQamg/7ztvXQq1hPTNgHOaionWj5hM7sGk78LEKVYDrAUh5JYonYrJpCFLfBZ/iuHEJ6nUaNCV
YJjF8oAfqRwZjuqH2B/o5Yy/8jfE7sN2RaO4+b7hPyXYBmKOrVcHaA8DL3x/NiNRJDUMY/m7SbPG
Z0HPKod97WeIl2ya72Skk4btLKKUWaaSIo6f/0EmnO0NWAo9zzstz9FvWzb2Ge1eh57qgYcGf8s4
KCWGHnuHyKUGEPtO1qcK8v+MluF4hovg5heNkiDcqF2vD4AoUCSgeQU9jnTuY65SuS/ZVpEOOL5G
/h1875QsDz6gNURehP2byUxNIxFPj2voItOhgGQn9M0UrI7VKsd50iYCmmDgyEHMzd9QqNp8hyyi
/QD7k8/GC9reukNC33yGnteCPRnhg13/pcTfhstrbR0NV2HholkfGEZPh8D4hfLalZQkAx4RL//w
CJiEwvqBDQ1zlJNlBwLtdt9uxHzZhiW5YDO69Yd/xOat0wa6CzjB4HhR5QHeBn1wziQ93HRnn7E/
AQZC6ywIiVqXKS/uxbWdnBYrTx7WLu/Ryi7w0HMWljNzyxmrg3GqvLEvG84thBr5qEivCUj1+AE5
LFZLiwjjbSga48seAru4ICtNLGgBuTAszg9nf3SmHL1Siv50jSGo3WOvFVSyoGKRSlGne84kDc1z
eVwm9hoK+Y2qWN53mvRnTIaA8VeUMjDfmp5XWQjAT7zWJkEGDWOdhBk/ZR6Wony5+na7EoyhmzUp
TDlRCZck0yBHsWny1IZgYgSi98KR/KCGgmQz0Ua5Hbh6XsmVDJu9dKiyLvADhTXCojgjLG1OLlIZ
X4NjU884ruyvBnPr0lUMBWPKwqAI0GumI3YXw1RNmbAelIPnmIZeERFHgyLErreSbnWdVqioaO5N
prfcDECSWrX3vLL5CrAwZGFqTCliG6HznuALO1Q5GGXfjsc7ahbt7JpVZAFUMokkXl2lCxDoFRx3
AQ1PV8lqcgb0I1bFaFJRJeLetACJWaLI+KorX+DoHnBLKcE4WRAeU9HH4iGdbAkZoxEBFWo2H1lK
UD8cnlEWpZToK1OJMBEeJS9qc9pVyKH86J+4vsD7pWoo+0SYCo3/iGaDTmrvqH5PfzOgFBU1BZFF
PKzzQtoRIM63jYHi0OYo377FmFkFd8V+Ok53xsuB9iOMYq7iftEQlCJoA5cxSA7UrVCRJoQt3kR8
sHUaIG1pbhQ6B7g2kKF42K045Dkrqu40JZCgVgYRmEbdegJ8+V7kF+JRKZD6sE1+JT742URnqxi/
GgSlCHXch8ROSzb7XEg87FaqnEvzvYBGvD5EUJ7sf5Vk61a/htUrmnpJ4ap50q6O7IZRjZvBBqIp
/QgT+8xZQgiXYNLnOwPxUWJO5iuTZ0Ad4BLu0RTdxgZhwx582l9bQsQQfN6YGVy4uyrgX+9338Ei
vOP2Wp+bTaJ8g7gGkD1YsZeRNUZB13XJciJ61DuA1gkvpLJWpJcQzdRi48nc6bNqS9doeS/AGO/D
p0ciBQ0Zkx910GRp1nL0qe5A8lHXgaQYI7psVtawz7PUl7932RdV5In+XAM8/iBU6tZIA4NkkET9
/Jc4T08qHGNbvW/sB76Q+uxtdBWwpC2EqFcZej9QlaHT6KNnWuN09Am9hg1GBRWYK8QCpeh4LmTb
Ag4PEdiQaSrzRsG1d20m/EiwIv5At7YEeujeZN9ojoMhNytDm5rAE4z86cqEQE2/PYKrS/wgek3x
DeIujsIVqNgw1VXIPzb1CaM1QSeJfe7Kl98+A0VvctCio0WC7esx7+q/5i9x95smRIh7g2HdhPKd
lq1TYMKTHsW3+pY5GiBUbOIk5GivWOAQN0wzx4gxuSNfaW7B7QzRRcv4DwfjVDZqCKcb36TvWZPF
xmOf9plxynSDT/LjkeaBFYw7flvHtwC+XNIrgRK/o9I1sb3o7wDQYgj55QDhfYRAT/rJCY6tDPWJ
GazQg2CFG+f3FnfajuaxO8nHiAYwieC66ur/dNK6Tu9DSm0gljLNvV7IYJ6HciJhfWxfdrgI9SPQ
dpkJdfydhq8BBGx4LNFoAIw7vx2ms7wHqDpqsBaF20i1jDOUUof4G621CCfU3cK1W1IyK/Gs6xIT
UhANydNOU7jjO3tP+fnl3GLxiMWD3v1RGbgQ4bxgTu0Sk0WUgxWq1Np3mqjA3O5vto01uHhc9W3B
5Y+amsswKSw8ukZlAsLyFCso2XF8xJEUruujPT7onnES67j/kRVyu2REcvd+/biJycEw7pnJV0G0
HJ/Cdyzaac7PzbHv1CPg/C1vWkqF2mBpfSZk5y/Vb4ndKM+nOuLOyD8PVgvypWaNLVNwRg07aq84
GeQe48qljN4aS724zg4UjwaxU/Vk2eIj0ypKMCNy93UCQ2dnHkar6l1moCPx0RLNPc9wbliAl6H8
NfK+2VcxLqGkeBdPkL4+bn4FErvy7ZUYdVST3QVLV15wx7uRYRnyn8QfmGPIusoLPMzOFuh9DeuV
v/UE7LXJV9LPO6g4yjMtU2h7ehcSy9IqGvGbEcFYDvG1uH5wbkDMY4Ru0NVXRSJ8Y1aTMOgGV2o3
lXihIe9BqRjw58hpmDhGxkJ3LWSe36gApydn+0mvIIJG7a4eGg/G7x64mDV0csZnlNv3yCl9BFHz
ESz36G1fteIxc2xMV8kxhHNJB0dkdxgZy8GUtZlgocal3ezAZG2cuJ95BCgabtW1wK/ov+Syqtdu
NWshJ/57gG3l9BjTn53pTcoWmxXjbvBJ84iB2btxO01LSRXZUK07pG7kWEp/0OESp7t5faa7+YQB
enBN1XX+6gFMmBLs9oaOBS+BIKQVWh4LiOlpQ4jBkDyknF5w1ZSAJObMhuyUrs1BB/8QgBBLSsL+
Ask4Y/dg+z/jG4jjksGTIiLfu+bDbB1Hb2rfxD3Nybqppxp2OvvL69T/iE6qZFd1G4t1TJWa1S0F
QEZxAlHcdLAcf5FM8H7mZuvOFKaHevd5lo877OMeS2A29NFhu1VBr1ZvU86f2W5BLBnL2Z+Mlmrb
nhNOOT9FIsVN12a/dbC5J2dKAD7qQDZCDgGBiEPxPlTtp/Ilt08J07/9kZU9DKIF4Kr2PK/2TPT6
NIDYHpzNh+HzHiEagZ0MANw/pMXT1tDQfG+wRKlOASRKJTqdBcXMe1ixiE256CcLGnOTCR156UnF
8YtmDDYErDFdu/TIkUuV/lJDAjjWfTk3s0KksOg3LfPZ/dVoiP+kmghoKm6z2c0StWBb+VO9FlHm
pXpr2HfOyfWiIdBpV2SiK160RPDtAEb1StpaXpOQ5hKZhJ3QFy4CYStGevFqwzpZovI8Pd/NJXLT
i0FSjn0ZeVBVFmrHbV6jpCScNbDGGW7Kqy1mKDfpaDykCB8z+1hmgssaYDUnxIHh5nh6bxdJvDsW
LBTw76MnDVf3QNGyDc9w/F2gMhW9j19fW/MXKfVY/EMUobx6HCZFW0nqxdbHMWc9oJM/RYPS/oc+
cBIZkO/vwWNUKYGNZSEB3qrZhFHfCh85T195RefU3iS9g0QrzIxdfoyu7DzlPC9ZqTRLCBUdFzgt
FsfwYGg/LNhU6tf0dbNnJeW2odnaGILXgIFdAOP9LV9wypwym3fpJaPSQNhESyrsOE2Bv+hsYU74
5HQj0YoMgkEjgV99SZQblwn2kH7qKjUSA7acuEXWcE0vsNoCO0oXfP4+y3YoK2Y9IJ9ffrD96dpK
bAq4QUMiRKv8+NKqcTSBWK7PEuyWoDRsdTljAkAAHoN+NgzPE3DEGQQgSQ4DYGaO2B2sFOh9a/FB
C92NxBHYDRr5CNTqdONp6/5K5aDPsK8dCCJgpRKp5cfdBsELHHKMmOOSfOEMxHx+MZMsobQgcFNT
oCvZXUizpe8drGc9AwTKorPYlslPhiaIrYWwDOmOslHsJJhCPe94J6FVmwuOtdULoKDqqkpNeGFO
vN77t3yKOp34PV/2r1TguzfafwVEgp0Jns8u+EUvS6LrC86wm5LPU8beoyldTz92izD/i3ovmBzW
YYmtbyHJ3oB3doW2jVLvdQfl6rlER7NlcZDNyB9qilMVDi8XZ+3QFTmU7F/5iGYw48uaA2jMbZm4
gtmtqkorvKRRrR3dshuroWGAzURa4q8Uy9e3L25rhasBjWSLZSKU1B17x45khNTEFrLtNWnECm6S
PW+BSthbhAyCYsgtqxmZlG4PgIWjB+HZtYbTn+/KpGu4/njvT8LN4h9L86/QU9FHcZz4K/8luOPa
4rHbU8z9FhQ61f6BRpvjXTmpfJi0JXMZBSCvf2Y/56j1gp6z3YUPNFzf7yG4h0ICZqsXlxBizYJS
HO9gjGQs3T6h+Pxr+0m4VzJLohc9vGsQaM1EMJtgl37MdH6khbGNhX8ob6bNTDSl7Y+3LYcFxN/V
/IyDHrMzRuz8Wfy7sldI8E7+CAjxv3ZA6aKwHTJYoytJ+emT6JZtw8T3NdYraahO5OzGdxisKbe2
imKq/UpbcKKiZ4X7eD5x1zZIzUHd9zHywxKaTZm96HDcWDG4B8Sr0Wy9/hrBPKrDVFclNWHWz/xG
6q6xIhPqUEcqkvgiopBj9bu9xNIeQHaJMbWarImbEipbiIbXrdgT7c3bKIku5o6jQ0osECB8osWe
JK/zt4uFvoY6+79lUQ4IOodCa++XPUPo0U7xLumarValfRDt42KgFnULRmAQ0sYGrMWlpBzG1bMh
QRxYdiMnEzfaGozAqViMTFWIiGaKYHu9EeWefNwxqOhDI2kdf5KZcnXhr2j/EZ7/RqbxLlawifH5
AjBqPXegQ7mjar/0OnQHpTmkgc00phFdA5sdmzyyAdKbqgbbzyfdQUwMs9H8PTYfz7oc1LgXnjL+
ZteuG6FpFEX/04jFGWqAgUdlnzCmmHwXQmRNasEtllUzWhzmlT1ijT1lxXkpjt3elwj7Lx5e6+KQ
y1cNyOTURSyOj4bV4oo//TRWJZI0BuOv+cCkIesZdpii/M+yBupk696MI1XlosOXTnFX+Eypp7fs
FjttGlfEm6VEC58pIKgNy7UvCZIyhbaXaB7gqSvQLIXL/RKBrpbLKUACtWc/FHf5tKD2FQCGuhpS
j05eHijmzL7QKBNOD4i55R8PqFdmXw9jcDorAyMx+Ft1ZZl3ZyvJi+dKGFsXuV4Ma1380agaiTk3
7KnE/jSNlBTQNtELMxotbI5yOQXcVOYss8rDUKmLasHpnq/N1E0fKsC8u0m170l9pt1Kh/kUgi7Z
9XB/16TAq4FMteeeR9nwdiCo/UYaN8m+0aLfqqpJiaBYGekbuscmIizec39am+E7zQwSmkyemPcF
muDw1ODTpITT8life3xRvRq+HGNowF9ok4dB1xObz4oaZlc6gnzut7laPsHDZp3ej73JkWNQKh3I
4f1JsVdQFzN9sBToFC2wm4IncXk5ueYelSaP3IhMJ6bcEZ/1+TrnPxicm3Zqalnzbdj1D5BoCBJT
/e994shpPB++HdnM6UsmAMEjIzek2XjeRM1Uk63b+UNlNeV3JbrKXr9yRf2YVXgyku8vlfswbByx
DitvF04u4VeeGbc1hgXdIlnRwiSgSOQrmRbf6QFozZF+jC33w6/8Aa5Zv1qZkvOStnDn8503hzfR
JmwKyaTX7JsO64tbneKLjILK/HyhGdMzPfZVKbyF7T1dke01rTn0Bd4lwNMQHkA09T77HlHLtzOc
Znk3remA79pNh5PmrDCrH7nC/SsN+5hcthosvgwVaDOF2dxb8AHX4QwztPNhBoZzehghUZgA7DYZ
iQeoBB2AtplEFUvpIghFwmpsDCZrR/iETxxjoF6tIglJRGV0Ki6xb+8pQwyjjrzUjy6gFO/ls/oV
fGQNRmU9VteSxgE//uHfHGZ631hfI39vOYybZXzqGRI9YeRqRY276sb2lD7WztT1wyduf6Z2M2r3
WE4VhcNLkUpgZmlovN3Q6Mst6y520LgUYtPCSiiIY96EwxvdluXM1VCFHSKc/HMRiqT6lg8XB+6n
a7B7e1Voc8+goRxn5HMcx8IyMuKrxTz0pwUVYlaQsuax0ECOzfXiiXjytxo4Hnm5ETPup4Q7aZTo
SsbFBsxA5z0vFEhu+8N8XAt//C1fkS0UnRs8xlD+TlsS99Ll+fBIkcaH/P5VXdTQWBycbs9+qV4h
BaOj9/4GmwWMGQSJDmRWLFMF0/6xUxqtX+YmWhLJDoZ39h9if4Qvw9/MmRGEceTz00pjJ6/8twsQ
3mCZrsJ0pmq8eaX4qJNbrwkvifHdrtVwrY1vlHcn8mOdIc4B14Y6h78yAgZuZhuYeWFdw4SfElGC
Ll4QvWO29IeRaxnf58wxXAcf0E9s44ET6Xwljd+0yV+pPhvf3IG5HOk/whyGwNMA8Wgk1yAd6GD4
vOGN2oThpCufk+/X+HpsTDDOKDZHl/4WeZrADaHgjqb4RnCVdDJCAT7DP6kn3a6SspGe63ntdvaP
jb8wyKuemGFOKbJmKt5V1EvnuD3KSxd3C7MXhoeb4iQVKSbQb+DVJeIQ9X83fV1sa775Q5nM0Nha
rUyFPuUGLLlj5NCliwju+PV+9ue1M+S6lKZRaZlzhmGa4CHmChOWPssFDoQ3zhzNEQNBnCMl7BgK
xqbHnGZgIgU6WdEOEVIxX5czQF+FyvdJkjxJ7AXVPi/s0G/AgkWbCtw4gcwUfwsRPxVTWQDKxKs2
dfDrlNOYMbeabIX29DxlgKoUKG5o59xunvuE5lsk7zdYVQa0jxSh13lnPCRiLvaIMpwuJnaSQHrA
QDX1s0HO7TwTSlpRmOZBzCInxJJhI30j9/XyVD38CUKkdeK4xw/nef7QuyExwzLkGhUZtGRdTK3c
THhICfpC4LaEU1ZeA/Ur7cgqCidMnTlDO5N49mvI9GsYQj4wXuokiUG5Ft4FC1X7b175PbH5rkDK
DS1OlxNADqDrA2qqEsGzzZNTAWy6TxTKFioj/Lmh/q9eGOeF+QdBPzL7Eifjui0cPAZL3gY7bTec
yRAg+5ECqdG64aQpx6rH2KyzMjmXpGIEQBWB94OG9Wse8gkcqaNBsVslqR6cQBvqOr7/3KcsVorQ
Ng9LnrooE+Yj2Bn385rPrAida8tG5RV/J3b7oL6zT2b0d8SvLh9vib4CktN5GPOvWtdfelElJ/vO
IXwnfX4qCdRHU0NM36d4+Pm5qehUaMGkJ87qQOhEM7brMwNZMaEn95FUJ2YMzsJUR3547b68nFC8
vMbspRRcLp9DWD7HprNSY22vZTMECqFYfJWXbnN45PUUHD+g0QeVXbDrvoUExzBqPNeZFxi0vTBy
jOIvgIk+Uji9Ol2vNfVRpdJG2hgPeVxY8Lg/xYdTp7XwYXg7nLg0ytoKv7adU1jk3ZZL0P08rZg1
o/vIT0Utw5QsnbvqGStJMYKrTuvncpajOLrB4B5K0Mc2mA/r+sDHQxPHPdu2QyI60gp6MjWHnk1E
VYEhb6Gjok06DQDb1dbY0tnerarLaiLVqyD0283i0Dfk28P/jNo5z4WwMz2O0XtS8radDEmTe9f2
LYCWJ+Mn2fXhG9JZbKlXRPaBhCN8WtNzD5KA8TSmM5wjg3rCnEVGiQ7XPuGI0Q+M0dUpxCeU05b0
GGkVAPEjzvLalRcTe00DdO/McpOaCX1+gJKMdQ0khhpwC0QGReBp30bu+h7YF5FpSKtSKEcgslZw
9eevglcksVklaHkp1JvmMKQB3zpjWDFPaiiQEMGupwvXOO8Rs0pL6T2Wr0ADITGCbH4wiSQuqjYP
NE24qRyjZ6MWGae0zjcnxQoVaeTIWBriKsmfa+OrymHwaBU0HCe4fKJZlhZetPCruIEbgVPhT8ER
7e1hPLVlxx/EHCJ2Xd5nOox3bf2h1HmFGZoeWoEm1kCSS54L0kenRntmGJPwwjB7N+Ywk63HfvVC
LgM+0wTjcC5RMGSeEL/rRRxYsES59zNVSX0YTzj8J9CdvCZP3V9gzkrn1SCnD7qJtbi1B2jUlgNj
JXUb849pBdmSqQpL3Pqa7eHwPKOLoku5ExhGm8Yxli9l4SssUsqy9GBoTLsYONwq77V+icw2ZqB4
8IU7RIvbdnSLQ4mOqycotyW8y9uGtjn5eyyGBG8hjKB438anWNvr4DvTQY+PBXXih3c9N9YDsZkY
OyuN++MXUA3k8AmYCDqJHAJIUbbjvZNvXvCqQ8F64reuMpJr15Et0GZl7MbAsY/yTH07dfFIfIbH
HbTPPdJA5Bf+WZIC7Qv7mBWcKfzVqv0wgEx2RX7YijSdndUhDyywG7yj0XiAQ2Ss9XKJf7JsRkd6
6jP5pzJzdQXPy7BR44wEDiRcraWV9iaUPEX+fuGK6KGB2XYDVPzdxc0F1NMAfg5ShzA5JAAO0oqN
BuAgo7+uS/C1m1ZFhqq3+3gdDFzxXbfDDlFnjF45scAynYl92eHYbtmaJsnaa/QkupgxYfnK+iCD
WyMmsoLB6q/YEnzEn9u92KDPlZ9idehjRGW8QWRYFgS5XKxL5X/4RcW0SE9YTsEUMAvEPxIJHU8c
cdBhR0cJE6+Fmj+2rL9TMIbXZYj1MiGkzG2sP7Ecx4sqMgrzAt1HkV9kB8O7wnyK5TUShfUYR//3
zCaD3JAOlQLt4/cYJpPJ+Tg/TcFBbkaIGfVnH/FcV+PMTNWITXJ8vohMVxkHvr+6M2mSIAzn9EHG
d6qVAoy1FcVunbZdDMWejUojlSYWlCX2dJ56FJbaW1/VIf9sqS1krcbGOa3TzNutYQCXiZeZb632
vHwLHRXl5ZuqNMxyo8GFPVfccg9K3A4LfFOXiLmd0XtTQPdJeTIMwc0MPh6gzwcYC55BM295YFkg
VUMfVx7Rzi+Ow/QRawxMNcwfOqnCheCcXQ/Q1V+P/YjmHkRdD9AMbdjb33cBFOKGd/KYYy4YsOES
mBlStuP+yw3FO2hMe1/LeKxL2Q5/bnPgNCl1k4KYcVOx8UO3Q9pPjDtGNUgQHrKKokdj4ibnNYtk
gZJZo/I27+XItghRUpGgUxLAVx7SYWtUvLdyuOECxdgVUTGUpnUyMogqEZ6JojHOW7pFYHIKGpiM
9zDKzwvnvfEDProO654AVeoQ4lKCupfuKnCD45qSO1Jt3m81yYTAt5AV6Xpzojtq0L+SACXtakMC
c4AX3Y9FJ+tdvGfkcAMcXzLokBD0JN81y2NB+WVpNS9b3+Mk3q6ZauZnWV8c5waDylyasWQru3vk
AFVBOwHM62DP2h0Lu/vq7z8Y3wvwN5jNeBFuO/nV+q9kzOQ4NvmSQrY7oRe9wQ8vSt1G+mZK7ILP
q+A19ppRysI3Hduf5KQse9ptLpD0EQKG2bBQt7PUzJZ7CHUAfoAzp4poGkkjmqXtS/pWEiqjIKGo
58wDTokRxJtiOlJQnOpGVzqFmC1n15jgMNCQtJjWIgZfeP+H2W6jiAzrf9Xfaw2F8Ohqa/3hDnfM
IRUsJSLQACvEhW5nFR5x50WfFZXrB+uGnXp6xNalKeB+2uJ6W7O6ykL8B9/WPxnrHSpGXI0Ay/KS
YaHgUD7GT8EuS/8AYDgzTPOTkpglNsRSLnJwUsfSII0K1vsfBKRcO7UL4aKLES8dHIjB+vpOqhrC
ZvzWat1lkxo981FpGnB6nRJN31rSGkOvFpKdKLXbaj+zxcqqNx1T1p2okRZc//XHTvH1pMIeE/cB
oSU+wto7lvhuwyTpb2dGDaEIc3hbt/pfCSuHgC/IdHXyrCBYGI3YUNUZfb7zN8XR/MJUFxJsh+gG
0qXUxXuPPNt8RJ/F19a/DDLs96m1wnFPnROhJW/962Yp6h0Apdp1m5azaEq7gclKd9PqWIJia/IH
7Is6WnVEFxWI0ICV3H7o91EOp0nloB27xqRleim0bBMei76yQWjOz8Yuv99e+3etjiA0gH7jorrt
lmXnXSde84GsT1qqX+l6XD9bxSg5rPdVVvDLs3iKKoVSuBZQz/QCiQu9IItbsrlRwXbpSpkOodlr
MGi/Oievqji/WxjxZCqtICQOVamL/PBnXM34Yqu4mqWmH1dbbJcw+RLy3l4gWLXA2ZR1pwtWWQ/M
UBGSNfBhA5kuUDaS5vdOIDKHVa+GGEwQrJtDYs5LFf63FBUUUmJijqUwpJKU/VerhAbTD+X0VDiQ
zlUcT7Sz3j6uqIotxk7TH0pczlXMdlCOql7VR1qWEEL3wVWoTEjRvjJLe2CccVbSK9aDTUxn9TZF
JcZsgE4C0AaQi3VyBNifyTGc1G/nKjncJyOUPMT6n7zg+zZWqHhgWlISg7wR8iEtKVfbdNIC2sUM
t6OvsAG/66pnmaTaQ1wL+wI+Ao89Oq8af/KLX1HfDEN08GJ3u8za0mdgp8Dl5dkatIXANypByt4x
v5KQw42YMgkL+i2qM9ENZ7/hYXrE9DQ9rqKkTWJzPZKbjiqrCg/hsPSSVthdfc/7UY2p+bQmmbj/
Q3M1M4wplxg4GJkZu0em0CwDEhojdxKaD9LnM2Pk3EGsTuJ2cLRtq8Pw/JUb+7GbXZvwtH5kYhcV
CTPNIvRwscjp3swU1yZhlcS77zNZluunB7vI9wSdkqy0wcKb56YOAGbxGS7sQyU0SS1MH+Gh1gfn
8YJy19qmz1SNTgZKG4fb4aef/BwaBlDXWvUWqoKscQmUK2N3feGZ280kZ+E2infFZnynWVcgEc1z
8sMt4s5Tic7GV+iGsP+/8TVyv3C8K5WnbMvthw97t50IfNIFYeJ2Dzqc2RaWJJITFkAU9IUVPxLn
MT58S+uJAJ9fkbX6fgBeKVbma/pLryLt95VxynJl31izvjdDptshdJx83ikuqElB3g9rWZcegVTv
bQHgB7nRMggb57OEnOwjw3yhC6pTuZzl/ItxYKIaBcNocM9QM1+OYPwn+68fVPk70A2/0RX7dMZb
jWZ9Qyg/AQByillDsEzsE2HmB0u3KuwwnrPVYJ3ZNrpnZmM2L52wPDsStoQR/Xdssov6q7wm8Q0r
ETK+YBC1EnjIrS4gTE8CKaylabLVxe3XtX5urf82xx2NaBQ+ypaaKwk4h9C3wA43VDKfPrsUIu7H
e13dzZYsZOdQMUpoa/qFjCv072L/QObnHOCKW0ltKUhsHUdyoESZbfzHfTXur4i1mAO5XFV0KScV
Qhhh1BFMWtFzGGnZfsOgeMvTldfceVM0WOTxKbInzPrzJKTEy65l7LlnytvIo1jED2IAqMAwfppD
YLuPOUBqpJDJXsXL9NWIowZXeuUGKx+fMtDqYiInnlOG6InVH4sh1YQ7za6kITfjT95wAOHQ1jFU
w+/b+RCvBxuoP/zT3LR32snBMnUPuvXAtbxWv0mtw1c6YFA5rBVBDlyc1uIv0kJxMqUN2dPp2CxY
YVlDP1nABA/iEBDd4Ra2lX2jeU5PullZMBZ1V7zFOKZsgF1kPomcOQrU3D1Jef0QovnhefR43qgD
OME0BbSbU4N15VxMfnae4C0R5PMX8dYxQUp1MHj/C56v42zUhBT6U+jf2FLOpcbQIBr0Ppe+gcx7
ek4misBy0+HWCGnLuD1Mt8dMNFVjWfudEmtcEe82yI/s4bDiGKuDs2vGTRQBM0jm2xeUk+wpKsfx
7XmhXGcK/dKb2DfZhSCA9vb9kCjoe4pOOvrq2YBuICgTbp4ZEAcoSJLN147WQZ/F3WZzDYdOXlxt
Ays7bP/uNl3yLIRJpew8SJHxGvKkpWqLJnzvYyq/3/2vNhYM2ztpNXkjguNGspdz4s/d02IxC53n
/Pf9e2/iinyX03cqMFtXBS6R8t9wjM5MW6CeOl2qpU10jyjlLjhcsFGBvwXEi72DGABhqZD/ja+7
Oz8ce2FlFwtw1/eOPqHzdgb3RqH6LWwqERHZu+Mh3Xfk/7+1VouBCeMOKPCBq0D3i8It3rIPJn2m
AXEInPB5Yn2q99M+Ym1YrmHM8nAPiuEcD/0Fen4pnvTjeI+M/Tv2aRZA31nKfbaevYHCrlNKB86r
Y4yJSC2Whg1uGQ3Iu+fAV92d3q56Pgt01rbnPLRLlrgDnjsNUT/CpZ8iBvw+0WL77w3S9xVudmLM
t9nWDoJIMdBgJ+8qkYV8gHqUrdusvP3rEGH+XPtWgvIRy5I42PYkIuqkGcFgMFnUABE9bJU6AzDG
qUUcyD2Vrmi8k5k8+ujYc0m+i66omr9jL07PXjmYTBWa+1EygJcoqGYXHXS+CxYLirW6bXV2RPn+
NwTnnjYVyqUPJQfmmC4zvidBzMoNR693yJLmrEGs4sMhd7bB6qOUduFYyqdakvlyZBRZ7xyDlKbD
gT3FVsn0OG3yeB7cyURqsbjIJT3LAvGodETyg3Ol0LMK2smMrgXhegv9y+Vkpe0Htl0QGZRu7YuD
EvKK2ciZd4r6SIpOz3MZmNLMIMhfX7YnSwjv3RYZ+SHn4tcoyHgzeBuzajg6Pdxwql11YMr1Nt8u
hgflkMiWqbPE3MqGBZItJbnzXrTOOPor0tZg4m236Fhc8gkbSTrAs1JBaBDmvHkVoEzoCqQNR556
TLbOJp1lv+NcATz6mErBvhKOE4kTbphYHViRoP20PmR759QP+3lZocrWrjvFaZkxRoJLxGx7RTrJ
j93/txS0GAvnP8SeyH7tTIIAziuD2/YdlrDNe/WKiv6lq0gnJwqwQhzc9rsEVs/V47fl1jTGndXr
X2UvJB9ktR/oda9i/XrdZRc3o6yNgrOaQrAHdNqNKgYj0aSbXgqkdl0OOPThGrdhK0BGfhzGqX7P
A7jcQ/IidWMLDbytsVWBvPVy7tYCfA28aoTYLpUbz0GBuKdVwdFQh/twqdVClOQjqIjn7InXv6rm
sUOZ6NxiatiA0ngkHjU4yVg+mOMfRZVgFQpwjjKD1efVOUQliH8kPpRg5z9vV2zZ6mEcM3TRjz8a
y8cLnW0mowAATR6nq8QwVtSPFWFZZlks+BIgKIWuHnDlPSv4T12tc6zcfQrReo6JJzn5dIhkS7HP
JnRn6Jp0I5T3BbR8lnWGQbhxzoKvctOPzdBgWhleUDbU3IuW2Sbf6Gq3YXmRZIQ0LVnejrHIy9FZ
1M3E8DNVbdViLZlRro+cwjyKJHi/FQW6qnJ5BNzm9YHg2C7/YmlZojZ0pnRN1b2qdSDaO7+L6gY/
7tMWtH+1jVK4kdxkiqSdbwgnJUrrFlZgicRneouLEfOAvczvdIAVG4WZvn8PjA7NMtCur/BlrPSi
KaicBCF+zZF26fP6uADdgy7GTuRlPDWZZOlgXkpidIeGLaPKnwcuvO7oKWZY2FVHGG6LyO2k7v1A
sciXm0Oe4gRxK0iTdyGzIptUIQsvH6RaNtSKAFDyVH7Yhu1wF8Zh52gu32EJG4wvv6/A/mPF7SzT
+8/oBlm6pvOPHkMvOUG4NN0GbU1hMRQnbL+l37QQB+99EoRSAxIf8LGZ6s3weAajsxD/KQFA1aiL
58TatJXliQvos4FaF6bIjSlyVvKGi/SKRztkzdbTHLkUF5ycoW0iqEabHYZDudy8O5Q9c+EzYZav
5Go4ZAaAW/tTYwI4kbb4CxWK/7zVX7/OP5A86wt5Azp7oczonHVRGKB8BnGt4ayB3/k9AX4RhNA7
mdebow6Y36rcgeskGWRPVR9rGahMoJBYn0Q2bab/WV79nCNYxI/JUED4n/snPLjdfmejn35GdEHu
4XxGe7Rjd2CfzdFgOY96VB8+h9a4xke/xYrbEsVVLQ7FnFIE+NjXEOo70pwklzU0dQhSUW51UFI2
rASxbGtZ4PIXts26erEqd0bqdG6lKmjxApcwIN/E1l3zP6j77g+3pRNt/lytU9m7m8v+/KRJh+/a
YRRTOge+aveyVU4J3nmxiOYPyNnfxF5VFdUe0c3U7MbysYuK/oc9KBqYq/Ea4iaoQbBIPRFnPIUL
hAetvZ4maBIWruJ0UrfZ74x+O7Q7By8uT5tiiVwEYVlQK4gkf19GFlaxEwTmGZpAgfQi4JUTPXCC
ZJenmPIDF6JUip1mqV2z2N0ipB9WjNbAse8dirWqVYV87sJmuzks0Q2XKx9ODiKUFNqbnpNhXni4
LF2tH+0XNxpih4jujR3/H4Tt1Ha3ki7d1HSV2wgvvdB/OV9aJKTSNese2dpULg5RuPPAXTmZxjrz
fMpu9UGW4JeuIlYtgVMbQ9irA/t118+ixCTqaSoZAIx3OMLD9YfAciOzxtW4MExUkFX+y4sEwhh/
aTH5/tbRMQ0k0Qg4PI8ObQoiPsFKR/uLcSLmnraT5c+U3UT3wcVH1YNjfXoygwMwyJdrwno4bRmg
SssrWyZOSioIRA9xvgdq60PDFYj9CmZg9Fej/liaB+cl5PaddmRxAaDIhCVv/VU4FjIYsOtIn74A
0QGYfDGUy0v0Zer0SQiLgdw07dFJobNyZhS08tcPyQbUCAVOz3DLl3xdOFVI96gZ8va+oLhs0+Er
RgsLbkh0KHSYbteboCsX7n0RvP+zeBFIsaf+cUX4ih+3UJQGaaBiLgn6vemqKXQwV6qAFuUiZgKz
1nuv2ExvryL5Xj5nfKC1eP0VW+lDwTCqxJRu99KGRJp6uHlja8qWS1qS8e2+u+q+ZRDYUqvD4by5
gmTtwCOehf9jLrx2qMQjf7E25eg8MIhxXqSbEKB027TihESWLSGLSwabYBAIQ2r++HRsUoXq1dHJ
hA/csavTTdYInpgGgcoyoGiW2O9+ocMIWGHZmMbSLODuL+XRQ+XpdGmfbJO/yh49/rhm6CN91L2h
+q6yEjaKrKoUsH4Hxbx/sM932tPOc/bmoP8T2w9GsYNs2jKrFllCwfqR/eWHyPDk8i0hApDO0Mfa
KfSpVxRJNtn2oz8ABdfCXvL6kKGlFqoJd0D0YoJpItSFtV+kgsplq6T7crry60zQW+orh9rbigOw
S76ylQuCLi3K6E/xp8062Ji0/9q0x3a5cHm2XRU9xJ00KajCYdsgM+1zfQKf5ubXlWuz2EhJNYUx
fzafcy+vDHXH0PJTjCs+UOj46oMWNLC+Uwxn8OkALYqAREmJC41gK6+OWP7P+rRU+BjSP4v5ZnhP
epzR7JJw4vXReB8e+dlekkyhdhlKH+QCzORi+XP6iXYzPPPse0jgLMQ+1CBSBPyhgxCkkuM3tIGi
aamg0w2x3qNamd7KAKLKiQt3ZRiGn8S0XRsdcGWL3v+DFef/D7tkFZBbxXY36uz+Tqzjwx4ia2wF
mcwkYiF/WePV7qk39vTmWoYN29Eqb9uxVj7gg3Xhxve72xhGF3ERY3QScaEaT1pcaieb5L6i+3nP
Mt7BMTRDfE6Pa+AGDnu27CuatZKF4QFx41WumopxwMlOYOVBZM0Lud/5KURPsJ9LEJ1L79oXFxTW
G2k0jtAdkniR5R7gUIYgHvKW0SwLuXe6mjG4PUNcZGhufJUyDm88Oz834TEAQArbqWZjVtUTMYFz
JPc7LA9+fhg7qWY4h7/hack4EeN7enEt5do8lcHNKbown+riSeS1kDTq3BjC6AULMwIHsYiArJ62
iO9GDeeJqMx1pACjusN+xbPfWEFGNT1Woybyw2tIO7CF5yr4Bsoh1dLmIxpLxMSUrLLnHZKzB2cu
zsufSk0xiBegLUUvVfhyjaDALzxGGOI2jCTesDBmspnr+vidvc32kKKcfj/srbPpnfmEtVeLB5ej
R5zMGwWNqUGDXc01moUxZDG4m5y3hhDrF/tKdBmW/33Y3TepnbxLTMjhS2lHglzzuwjOerGmS9yb
VPPQpXMTucVV3IQrxixH4pzyG6NlVaRHOvOZAiXTivRAolNBQ8sYJvjBE0tQXy2dw4uKSS23qlMy
sIzTidCPPz327tkUGyyxyhef03H5O6huP+tuH9KGlXMrPbLEp8Hrdh5HfMxLqRX4YqOBTVHmd8My
hOti/hDq+UBTpUWOfcU5+mMvLCw9eYAvIp1xenhQRG/oc4g1jKu8x5bc3kkTokZX+c0cDFi+8X8m
hTCvzY9VWlOQF5SLLWrlLnGw2btpj9SQqGZN/gW7FUXtO7ux/7Gh4bjii4XtgDAibPyFjPjC/E3h
eY40mvxof826FsAGTnRoVI8StoX6iu+ntA7ck27LZfggLEzi51ZJdg7xd1TcITUYpyBZqwQuYilR
1gh2gW2BgRhspHvBJ1rDufT/iRGR7yq2YBBThk2zAfVh7O+idZM0pSKzFhRIzanKID1ICDsdKfuR
mi2+k8qV1bI9sOfa1y3GgD1nJY48G97/4Vi/OeS2ADWhEXBuy9avUghkdCnuonFmu+I5GvtXea5X
2lUTBwUZTbcTXk8LpDL3h+OA1oIh0rkf6ha/eDNMnDyLAvkayKTzWS0spSEstdPskW6XziGCGV9H
12x7j+uLanGdHNPmqOZEp/8SHonQpy10AuYTf+pLqqmZ0ZusU6N7F1Dw2/HZhF1Jb+ZR8DPjlzws
R1SluVHwAf8r/pIXSGVdouInK2xCP3+dmQu1mGL9o14KHcntG8Do/S1x7ZNOmPuabIUOlr2Iq6vE
WPlJ0yzxcODvU7YMDcgI6lXuQ6JO6kDDMztw+cS2geDWs2kNZJCsTtUIUdnuZPF8ioL2nrqdHybQ
s0f67pakTii6biXVG0zlv1u0EIlRdQ4n04CgBhObTbY7ph4tM4BgKBwCxkrTp1h+jhrAYKSeoI1P
fz8tFEmbgfW9LELN0PXAR5XPcQyNPSgIAhoYYg4+HVoQKJBockUmP6bC1fiLxeG9k7tQAvyFtxNC
85wKZr4JFa18+Jg0Tjl69jHjOWbLq/7wDdnSAiIZTipmA4PzvYeJHxxX1PEe8YjYYc+05rhuqosT
zPZmrm4i3OJ6f2RuowNZ5zgiGCm3lF09FX12vUD2mG0RzroGCBH4hH17MzPOO1nm0BQN45Zy1FY+
CemjRzXSlTFhTtg2fSM9M96ioOGX+t1FWcG4zdY2AWzZQzvvEtJYB1KEXiKlbuff6HxxqET/JOxd
I8OgnqlXtnvYaW4163X+AGx8LG65OYvyTV5Q5D3CQa7M1EpMVCiN7ozsqvYDBMnKyHntMMCrrrC3
4uRbPUAS9hQGVmhG0kSokxVVgKaB8pokUcO/fgA7U6P1La+2uNdWrcp48nkNiDl8bI1mYf+S62+S
Uwf4d4v4i3X4mQeAz9PcjrVblB3nuASG2HMYsqyEbjPENakBDKWHltIoxuc5vOsTLBbRIRo48YGJ
cxWGHkzu/EM5p7DOUEPO8hBoSUtI8txeXzkMD2/4juKjvKQX80RWp1DzG+X/VNmQ4lfvfp+s+C+h
/H9gVMPPuvgfdTPbjOS5HytFE08i1SAxG9B/EMoFUtCK0o/LgThYoosr6ZMIlhpMLVEtipB/ZYjm
fGpEe0wHAjtdUf0QZvIA1bhhA9M79fpuOaizAYC0JPvFx+WsSEOU/R3ACPD5mrTAET/C1kNy0y7a
S/Z/IWCNlNFkURvFdnFpRsQb11yCK9bgWzvy4VpXB51r1BFxMFYv7mtb3JoYBbnwuGCLJu4Kxxtt
yf3QrKDW+PncOMATcSMZZSZX0GXXIckGm1b20L4o9ym+4SrzVraabdsjlEMqlgxE9n/Rw579KsQN
Y+viUVBxdZt5/1ff5XVuR98KNS43kYSAI9SkhFWMXb1tAjnR/MKwJ4VIBfH1/u3/u3AC2lhlr5bj
zF1Uf+fBninA3Gte/2Rt1etMU8NgGo5Whbz53JnWGmlUcUSNuvitOJDFuDUa3SXzcvzAAAL2B6+4
/CzII551bzdZ2D4ObQ8noX1n4KK788F5U9mwp7UwxgFo8avZSeumBZZ0VQhvI+xhfqGEWdC/aFF8
OxXe7/kGwcPg+Spdg2gL9gC0+VpQOAx/z30fzxPpVMBkwuUU3LS38jNOHx9zvdD48t5mw44LhQPS
082TSwtlL58qTqaQrEk3mP3K2+ylwfdRZHVRUzt4Idn0riRnBIQreU57LNJRt8rIU64gEgeJxvWa
lvnGl5TeEf3hIEQWFASOMjS7UKIjGFnrrnGJ4sq+ZFViDwx56/mTpyLYJ300zpevi3YF0hcz/9Qv
s+M6FgLVIKZ7oA4/mm/+BPC1H7pvAx0kux1LSqOsTcRcef0OYj6c7bUROcI9wyoZulCEivzQy9pL
QZwmFDr5tgSezXLaoCHCeFeWteBUBNXVfBQkaapKfYBz1LYMPZG4sWlYx7lERwtzWmQacqVg4e+l
MJ2CoGvnNnDyuyVC9k9kD2df+GXsOhngR/W+Dsgzn+UNrYqZlkmz+CbTFpv1qkIQu8vwAxbxnw3S
0SC6qz+tX6J0w8XY1eO2yZ12bVWFv1w/+HbTRNYvZM44IDMXxFJcYIGj+BCrNN+0t32C94lPtxZX
tQ+nvEchu+7FfkLosfEUjBS7B2u+uQge6A79mc3Blt0yKk1U0MFfIu78XtmeP+yvZcHTBKX/wg1m
G4//qXdv4grWuJjS7Md/WvbzApn+rntNq1ME7mG1ABtxUIsYJ0bBo78f5eNUCdKDVcAFdun1M0UT
P+6NeTC4XA6p5nT+AMO3qzosBeuygdEyUiYROf5k6OLcOQtCT9tic3wodACLWaOfeboubdG8bSGs
Hat5Ijc4WNdJpb53ACjtkQuP/ocL5w4rkKzPAQ2NG3I9CKpIEeDD9uGIvX8A76tAWLOpXeF24mCC
+iHvPxUr5TiTjeFw7loUQ9+EnBkV91022pxpqeF95Msig9uNRrBfET3LynbgbbBGiFcUOI/OX670
4ZYQ9FiriKLUO0aT9NCXYgU0eaARFYAoY0ScK3sMV5zktCwVj6dyaC4e/sWavQY5rQBH3s2pWs5v
oHP1xrHF0qxyruTKBQPv7lN4h0LDU+2WSZDWGGFwk4PRfho6JipqLk0vKztmXVx5mmULb/omFITZ
gUPQCnyyzTGDIcJvIFWdYd5IoNq+dIl1e/M5IQZ6oedb/2C0bPFYE8nP79zMdydimo76WAq20lPP
wScXA0gT8DvHZUk2Vw7le9Vscdmsr+XS0puWg/x8muJEV0KqfI9aeoQ9jeuQWPOBhujbZolYDUGb
knZ5u0gb7EldWmm0InOVtLzXiedMRkGiS/TPbhH5AktYn4Xa3+Q2Qij4/PaCYfuwIM2uomh6VsjD
I+3Mmdvl8zTwPx5XoYUK4T/69mBwoKWW5kyZ7ke06HMPqHXWAV2OVP2VcrsB8Xh34DwiSJs2AYno
YSoj4e18yxZTIVLGgpkh8RaQAkwY6CrWy7Q6GWeljCKqi8xo3M1lldzR8kdJWs7TgVW/MUQAoFkl
cNKk3tmIvZI5TSYFUceGe48uwUvORm0csb0DVKkXfxYimgGgTPkoGA0wbs4GsyCIEafcQvIV90nK
mOLZeX9UVQTeuRqSFqVtE/JgcfvVtwb7vjbb9ucnjHyStNDEV7uvyEeTgxK2mbUFpXumkhZB6avI
4lHI7/vl+HeH25ZJ/Nw7GE9fBbg/2zATmieDmGwwIi7bbmRIfG6jmCVqTuDEiiXH8eVJCtiTZ/Ml
mUa3jUNTDn7q/wYHA8xtgG93KN3s/qY4syVP8Cw9MfyUk4IpOFKRaa8IO4wFu+NbD3JVmbta2D+j
TUVWrWp6ZUiAksAOzwrjhpOGvDo2jeqbroIi2oujIhIrh6K43xeB+LiVDUU6hswjS3OdBaI7TQRW
KPhFC8+dc8QaHeM1fT2AX1NMgFTM8Y2p2Mghkr4Wt85SGXtk1AV9XKpXvPKfKGBVzsZQeVfmGwKt
p9boTgguqgXj+9F58YoKKieCMkrtvcmiRQJv7UJ5p6mtVKhZulpLeZ9QAfyfulcfUb/HfcGQHL5n
HV6ooFHM/nSRicONUAScNxTkrUOY97dtyrBb1rzPwskqNbEk6XMuW/1yNdmnX0W7xH+pimKF5MhW
VjFrVyVs6Nh5kF+zSLWBnFvIDYCv3ZZNZO5l7h0oup1Il631Idq+s1rgF2Z89zG5PbBG73zJO7B4
SKsOAybyb81q/MkVFQHlFzAdVLyUn93x1dazEZ1sfUsSVbm9d18M+gpMoD+rVkfZ2Hn2rS8hfLbT
ifKrHbAiXwTLRMjfU4vkqvkhejzJ52fY2Itvz1eN2d07YXpN3FFp9eyprSxkLVHgVM9Fa/dAlUWI
rZhtQ5Ub+RSZ9MDUnE7Sw6MpY/coylvAW++mDvGIOq60RpgdiRYNBNCYP5njvNSXsx+bsgRsh5VV
JDobrCsYp+AojAAVYjAicmW6oWKbFLsfFdMRwGkjrVhdlxFYWH4RDofjNoSxgVqVEVen/LKKKd7K
0I0Zd04dBUdb2FHSQAdUun9MBKBjNA4q3t1ljUMyQ2iT88e+LAQruzJxiH7rRzc+XtybOk43QtF/
lS4SOzbg80dr5HoYCbtVW3RN1bxL0Hq9Bw3xoBT/8ZAANB0vKVmSU80BpYhrpF6cNGDOwsNgl2+p
SKM+oYYZAbUyxGHu1TYWusBtV7KAtU5W5Nnq8Ou2drBf1UR7gd9NoL1K66GUcPzqiIdbUAdnn7c2
4Ah73glvtbRAQwWPg1x1yqr2ZlM2HqbSqDHbogpbQ7Jmsm02M/HqT8LFV6I/0gb9WTD4CR7fzrD0
gQM6JBRlrAj0YmTK2DNTrQfxc2OBo0JkHe9uK9Wi3DJV9F5gYrpS/gU7NWqCD3bLN+VtAvEUPItv
Pzdhq2Hmn8huLKIEvgvOZY8So87J7RPF8DM9a9U8O0CN0iiYIHBHGkt9gZS+Q9lV+QE7XpVkSr58
SeZh2eKZr2nP64XvCPPL3sA1vYnnsHLIR6LxG3rSJ2FD4hDRYRy6SwNpr9mezUqHOCHDG72IcjMA
6gyG6pbvdqHDRUJgOR4P96bsciRZ+azCJSsn65aH7cFfkS31UmW1sh07+M0mOXmpPj3RSuMQdJVv
FM99Y4P6Qakz30o0B8nJw5Hd/eLrZBMlSkkL8ZD5XkTCRKCRkU1XnsOEck3C8ug/HVce+glTKtPV
yGG/dURV4DSKhoaN/yRbeEzPhiqvkO4GJkw/tu9z/9HcVS0k8TcchnhL1P+N4eFsDbGwEz51e4Zx
BkwOTclvYDVyJyGqo832lHyJBoV+ALmgkdaC1f5zHE9nSzYEh4j1gY+JrB08TS0u1f5CFyXwE4nt
0fq76UKDwD2JzooqEkCOwdKCFu/o7xhq7/yMDWVi837Yzl/b+IRAkfTfw9QOPT2QxzzloUUUdZw4
qjeHFuNJYIhbq3TBirwtKA/RmapK2BvqaEVbj0htfmcFnqC/kH6fMYfRar4tJq8Jq2nMHWJXS/yN
MpqAJh/nIwq/PnovES75MxH31JqDSf1viUU/z3ERo+GLt1Vk3ew8AbX5wtk026wE1mNR39lkhgMC
4PToMuO8XyARRpg9LcGlw3UuTzhxJewR4oG0hohhl3STBaN5iChLY3jpRTQfbszbYfDI1TBaaLIT
lZrKcRUX4VZzb2iFcX+s2Dv8lT/Rc1mgloQLcD/ewlRpgPU9HAmDmyNu8Hg6T/67PE0A+mHn2mPq
ykdyL2A1ELRAYLuNFmagXg0xUY2iY6vEk/ohyBehfTR6uwmbbiEl7scKPs/iIbYCZNEtnJnGcAYK
vS/0tL9EO/7+sTloIGMvjD6hxm/CuLYOgJ7uSX5QYsLeVHN4ek1P+QeBxzy/SlKhyfgia84l/tYQ
90EDEZ4z9n3WyvVLOqrAtI6BxnGiHjrssiox2U4MzPQEIwmWb0uio9acVXdp+tN/Aqw36DR0MsYD
GrOnNHDikzdgobJPYueIrXgIu7sjCQFsD9qofg8i9ploV0bxYg7WamGukF1HScp+XmfUvA75tEqH
/NhZMv6SOc6odwd+MQCKWGtYMJx8N81NsT6m7s7SRv72J+uquRnEjo4uOHsh9nOE3+Dif3TYijXK
E8GkFbSNEWzSmQjH1FnJ/LoETGwnNsKg1b4AKzh3hF1WyWmAJNhwaSH9rpTsS9M8J12B4FFNEsoP
oXhGVEcMQBdz/iLlZSxzLMu8IM0qAtDNXawm23YxTVZmgm2SXBA7FOx/JgrvErnsmkoYC3EUIwwk
IKno1TuQDtUc5EsDeLAPhC/z9Jrwn5I0bPbTt0wd0wZ93J93WPdVoAH00QCpYhqkuo1FY6FL1VR/
hW8UTH3T/AAIB+90mh+P0uT3tAmMv0So1W46uXdKO9Z5y8gt+4gk8l+Tq2xpb5Z8LSx503TAmC5F
jr7ugRABW8tqAOV/UQNz3aiYKMWVPhzwVXYSVeLbj+B7eJQeShXt0b2PSJWLzBFB/FqagUV4lANS
rkla3AmpfdVklZDjRRaWz/qLicy/NGcQMTq2BAjDo0acr7J+R31q2wH5NF4EBL0vwxlb7ff1e9dB
imPoLXfI99xFkSIKkJ8NDDwvErrFoKvloS1wlzOK0lcxddu9BBf4tXdt+TXFCyzBS/i6HHcd36yW
Tx+zt1tRYeaArInxVuU5HjIZiq4hiwEnCeOWWz9mfCvlkRo/7BI0lyxs3ZAd8wRmkbPuKbxy5D6L
U9lDdfE4tKP1dfp/EtFuFjX5QEPAd1u/hzbhQUIdaKULFdVn4NDbUbvhF/dcWG5twnz+tedDArvo
qLmdz86SiHllpDJ7VVpJgR0taGUAcicRoMrmZp8OoxHm9H3UD1V69jiR4z4rhurcsTqc6DN6Lj0X
tu0gX13tmScujDN+Pa/MV3Mcr0ObNxsCBGCeFy41qn1DTZVBEGJMt6/Hz8xhukw8s3NF1mYK5GQ2
+vlKZ9PS2MZnynn+FoJA5dsQIqb1ICy2j4k42bqTU5uxEt2mgr/HnQ2QrpgUi+Feh9zUZj+W9uYg
llvpxcItd37LveE6bIT6J3c7ACuKE+N9nCGCdKt4Jvac7ju8XJMF3yhLoGj/6YkpJmtQe0FsjNlS
neqyIWkQ4zX4G3eVhTpBlGN4t9/7y4g7mEh4HsqZ60B+pKKjt4iU1BJpCg5IX8KjLMpFhm772GC5
9w2beB4NVTIKzBY4ylOa88J3AeXTmd+w5Oi707z4laKMdLbCHzYUl3nExGuliN/lTVdtHNGudxIk
nmws+bGjmWk7+4ZLH2wuB5gAtlnScvStGhCLfM407ejIXymADB+8aBIUb+FJPIa0AFaQv74nRliE
OQqSWWMAhxSCT0ohgBkb/LtTsw2PugSbcqjHMSwZsYMoEZXMBK5BDxUOWm0OzChFlnq0cqUsa3fX
s7UXnBhfG3mTHxLZiq7U8iHYPIXLQQ4t2gKRBx5BHjNZzARYCKI/KVVUmnwrlzqxSBRTPP63ttFS
PuSkQSOvFQRdets/l2HBJVnlCBLgkSrtSbgGfcfqKrwpZqfmRXAmRSmGi4APKDSYzsKAEYYrP6D5
dK97TcXRjH8HJzWBR8s6kDryWJLwLF2+iZ6wTsqUT0nH0+88POZkf4AuVUfUKQuk+ZyGm+cY3eMv
+VQ+JRUcrepanjUj0LO9899Mq8u0FPWbxGuMII924772XazhD+zki/Hw+w92TtiG5RDadd0iAlgm
q2lfwl9goy8wuTvXT9pfANU4sqNnjy8Cprj7K+vEiefZKJku638amlM8fI7U9UhKMsEA04BuNbWv
HKO99hYRMHXuJHx2mtbhGFShpW5F9jr0uVCryQ9wOLBtrOKM3ReAmH/qJruZZThIgvqr+amAn4I7
ZiUIz1BrU7OOFW8NuEr8MRB4uCWhIBgwrAH0XvgqX7pods0x3bD1K2YcHLgAC7+1rU+pKm36n6vI
Y/MAcO2KWI3lPHMNRg1fE4QZU0BHJp3aXggBLVTImNl99r+XsD7W6SlvTCkujF7gV/q/it31Gne0
5ukF8bZBvBJG1q2gS3HccaYzMiopUnSzafbSqAMBPzIl7T4LgPv6Tp/jLRVHOZ5n/DXp71blhFcd
N2gP3uWujL61alB8Sb8UVktVM0CctLzZqysLLsSVESPFiD3SXaOaHNTPgoM8VLOZkWCz8I1vdqyU
ivtjvakoGDI4yK1t9IGBCrH0KGMO6mL8C1xE/P3YjW2/LmEjrBgqTMo14Mwrnfs1p9UtenLORCO4
LHm64xEm738FdCL3rP2MmUF3395/DKXTpdXQ+/2aYs35qO2NncxttMt+o4LhwCenJYGCNWhSnOrW
XbRbU+xWKAgdwRCIIueEOaIJAB5nHCoaCwvwO55My8+o5VJOAJ9CmfLYWM3bOPrXS02NyoYXGD1J
X44mYVNyf8JIjCzNSHV19mrF84y3yhtVncIb8NPoplX30PwVkFw91NCqJylLJc8lBNt+6lgY9a+n
cT+3bZHzrU4R7gTHz1js8JD1DqSYLBJop4qjlC6ZxMviNHhTD/bqGTYEOWCf/Fofk7VuoQ00sF+5
ypsdsr0FIZr667kU8vjltULVU9JnJgzPwsXfiX26HengtdCcmHqBNaL86QnGycrlmRbQkSx2ci+U
2sc+p5O4V0kAfJ0eg5zve1JO3yWQ5FYMSD4froWEc5YiKauYKZ+b0b05/xz2kV81ci/j+eETjfg3
Dncetz/aiDXXaNS7oLatqluxN9LmpYyMcVdzT9gMvOeiBb9qwt1+fx/6E1sT9BRqwzPnC9KbKUjQ
fOBOaucm4eVRbZyhdYjQtpAJ42W/GwKTPL7zgI+5Kdk9fnzvfM4FU/qmkGKLPvlfFa1zvE6qYD0V
775ocHjwS/sM+JV0fuaPEiH86zCuSbCPMoA2eybC8AhrEe/F9+Z/VLXd+v5MbXYb7x+8c8Wf+Llg
qNku+hvDo+PdbvnX+gCmsESIgu8srGtlQpwS6IO1NatKJHVNeoXuzLCMQosw/fgD9qzRzGbWUnJh
hJKXUBFJpuxcG/3GvzyAmtd1SARA9E+Lx9xgZc9SeN0eHo4fTeaFhRVDl+LOsNaraMbVjHCGZyZ8
XVwkfw8iFG+VM1Vc9cmcMOMIlydK0uF0l7NjMQTdRutxrX2ycJkujEk9MT1sW+QBdUV4cykH5bg6
8lVddeuO6M3LWPVy+BIZnQlZilWyHSmJ8k7GUa2fzWiyVlTO+fzWBdsX3fi6TBV7WiwcGeYk7ane
iDpiVMW5t0wiSp6fOMXWTs9p4zVxe2uXeBXPVsp9Zsbdezd4gkK7Zu3AXXczpm6Xzt5hgeOYm9jH
y0W3QbXmwuP/yrVRpw7gMFB7DN1keV2TLsVP7zgsFwRTKz097mOlvDFpirt3UPB061NPWZXSLvHb
uPfZFzxKjXxmFzpaDUmJFxVjwOXoybAj2IJ70HPHZogx1SMfuZIr6DrSINpdVwjInJdsrX2b5K0S
bRAQJER/FHwUq9JL28/5fGEVBZTBRGSfKUDxRCrOMLPvkzuoRPSuc1UBGUv6B4CObVhU4sx0sDor
XTozvDc5pB0TmmGPluFvowZvCvA6sz6WTX7qG+nmbe95UdKS/EVcm0mzBYUkz8eKY8rD5FDVehUR
ykrCeR53x1ar6ACdm/qiLsirVOGDOTfYtzfFBtNLHMc0sz8Mrxb/QcY1SeDwP8XtS7WnWnIe4wVg
HwkKWzMFRfFd2bCtFj7Q6+bBlSEIAJcOThzFlfuAqhz9o3NoDuS9NDOikIuF93zl6MdCdORB6v1e
fPDRFFVma9Rk4/0f1MuyA1InkXBterv9utrUdtvqE//eq0u8b/D6zGCoQ3rw4ZHpQ/QeiQbPabEk
ODaNCJMMZoRCNz1gHHjU5A6F5kD/hSI2J4L/pTLLm5JAZwS0OKlAAYHYxtKavps6isQ2ZxW8TIoi
F1wv6CqUyWmgkL8f4SafBmOdCMPwt3v1Ew/Ug0w9pHJpKmc8RkMsrRat4mq9BvXVPc/7WAmseZg1
9O8qVHNYptrEOlidPFocFKn9gh3ZcqEEm7jzapgTQHdXtNjY2bBeIvfWyUb2xGucnA0yklsUk976
/qHEidizvg+AnqCdOkRINNp1db3qm7/Q3DIXgVakfeWALOpQIkxjd3AesulF7eU55Xqflw3Dpbz/
S7pQE2F5KPCQrdK3hRAOX6y8Kz7dImeSgUrQgwr1MJ4mFbiItKEed/RZE+R1G8duGHVFX9PPCHhY
38pox3BbhvGuNgO48PTXXV1sgIkidxqLSFmtHZUGPUSSJY2TPJWkSsvMK8Dwlc+QGQDFnp+ElwND
OMt2l9ybC2ynCm3xJgb9zS6Reit3BKAWRpdaWTQ4mVYGMEeZLxvdjBrnvxh1wdbDGC2L+mw2vWfd
HcNAqg4OShBpS2ZbqwTPv356EZJ6lMi6pNbAUDwmNz0yFSUui3ch1KcaEJwOagtxSwEuqMBurOA3
pjYe45wK8Q209tjDTC/MQrsnSap4EYEvo+LG9pGnLLOQIxbnIeapK6X/1hdGwcuurCJmVhkDJuLg
pPCTu9MedERccKHmyjaJbKMmMqa6jelWcCi+rFwQdxqe58Uth/Gs1PiqFp39RlacsBcg7MpR1k7J
Nlr1ZUU7TUlG83xBzGDlzUf/qtZq6/+cl84yhbI2q236QAe5FWi00jTQNSuJ6UhIRLH/r9AqEMEv
VYzqrE5jP7Uv2dFz0lrUZqmaLvtOoRs53T26fDzZncxIuzObnmrxHAcJXFE7+lP6BvHhkOnARVox
OKC7v9P1NUMEcxhlPqtgxcxEs+jvmcTdfdyka0YWVedoOKZqgHYbgR8WvBWNRrPIIFYKvv6QakmO
TqM94N/IK6wA5DGu3Ca51en9Z0MuD1loxfSBJ3HOIuVdtigaE5SaDOeig4VAJkVdIvCkal6cqCSs
EDd6NmkFjNJvugjRRALNCuZHzv5L98wjYtHtahW10+bWGDle2STR1jwnxgYIYBDDAw1HHomhNG39
4Y9VICP7eGWGgPgS29q6HuuMP+5dDOjgYWw+8Uqx6bP4ui2MmLG/7w3TzJcJICabmKm0rS6cbYh4
Hhf9a8lrrpXXtrxVmQ3IDbQNpOuFBhbMlZCiDOURgT+58b59ac8zA9CzhYXmNetR7qg9waSkhV0r
eeCI1LoVwELetc7TvE7epsCsgbgy7IE4yQMj7zM1p0MqX1OkRsHZYdnec9EnagdmUzli6SeCitKY
BhbOXWzyjee3Rl+L/bZjWBHcImMFeb83a7umacKy1pCIm83sCVdvVGB3kkNNWQtYxTI3WwkiPCdw
TTRQ0f9SKgvwgvt7SogCwENjPTQdGCX457skCeEXncKMxI5eX7brRlOKya19VX1nC9nr0Y9Gy5LT
+YDMlH8BVJsQkZCPdgKdvty3aNvejLIhxuQwYjoCn68vTRxiiY39RlWwZTSuLqteiVMG4B6v55aF
yp71yB2Ifr1Xv2ryABfxgIN+kw/qMCmj7cLZIghMjC0aP/4Waobodf8pay1CfaGH7bKjcTiw9FRX
PkrjW55iJGPOCDoZwLBN0JaiY62Kr9gcmtkIEJSsiTEdsV7voF5vQMwfitvTBxwKVYPEwuV7j0YD
JXBDp1r0lZzZiCCSChimLhLcdrsDR9npe70xQZmkHBByQ3K/Vz6AZrUJPUfTC8QOOgMRsSplUUaq
kUZEQ/peBfNeW0cLTQVhggWm34K8ZcVJBBlMTgN5LGVPemNwIsoEz2rNSogYE3xJBmS/tFqqc9cz
kXXtWi7tXHjbVDyrZQQI7E41MGWn78c1zHgQu5PiSQaUl938QoMsszq2rSOdfvZyMcNJKGBaKF1p
GKXezHVrd4P79ZOhVKKrnAiZJ0J3RZ6sOmz1k+c0QJN3V2Yqx2LgI4oLnAH4Dp1KKX5a0+bCp6u8
lBDwO4IknE32o5JO7jEg5NqCeGSewlXbySA7dUm6tNafyn3ju6RgjKN8/0D3E5hvcpjWXTn2JbLT
T79w4VQxiMzgT/KkFTXCA37QIz/TOVse3UK18NBLi2wj5Y2JMFRHwl4NbpdwPshZQhsljbKSfE4F
FFmoH3Xvfp5v7o4aIVl99Bgkyds3VOkFHlw1dpaEpNqxI5ZWfkmYEUxc/wfwiw8ipJ4kbRre0tm0
SF7mhi0BnqeL4AUQy9Fn7UNPeULgQZYUB9RRBc7faoc/5tkd2GsEUlly7fs3Jp7fmWyGCaYVIdBl
aR9+gca0ZAcdQIb2roOrB7I6FAqi2Q2WtrRpE5VB7TEU2SFunyRYs7ALCEdVaB2NDCVjXxdg3G7k
WreN7nc7uS+n21sZbsEHC1HUNaeUxf2usaEGb7EJQaMXbvL2+jBR/tSBmhQMUHiKIXNRQ3FXaz8L
89wur9tStFxj2ilA97lUGqksnuGXJdDLHB23RYIVS53OHZNPMfbZEL6+HbSCWQx3/srIwkH7brXO
yb4W7asdOA4TOKCswFeK67QzwN4PBVmdQsU44bHDjzfSwBDZVKAlbD9E/tDNSHi4FL0fXLwaPusj
4NKhf7b4YwrN5BM/uOp9RnSg1bYEUc0m5dGouQ9uOdns7GH0l0lCA9c//1S56cFdrL9Vo3KMJnqc
baW9hZ+j8s7vH0PpRUPN1gPr+KLIm1WPxJ4nrcAYhcx2d4biwiiWipLgb/ZjS4AfLwp6HTm5gzuJ
zYxnH7dEdM4Ri/X+8Ao6F0dkcjV/qHMhJ7Wh0n2lZPzv/ozsailUNMX98yQnxa4QN0To0kLGtYz3
2piuhaT9gDnW2OUdljLRiTfvUs0l4RBBHL0dV12HB4S2Yh3NrkB5T6O8U/RdOUFs4KPkaaCI8kBl
o7b1mYzcxEz/H0mSypKYsKOD627KEVyfbQOOANjoMU2+iKy2y1YX2UUKZBSpMDJ3dkCZZX11Akif
Gw/iNBdmqWDoMab8twYGLGcl4ZevnrU4FwdBK8MBYa2dWYy1J9cgA7um43fwZkcfnxdZz58Pblys
mHku2QFLwkQc5SeSM6FMuPxfqXxY7eqMtcWOCWQeApZUPluM/8aDbq4HIJ003xNlm+HGkt032tkD
77q1/z2lN7fTdTu7PuVnxeRrNE2Z1vwb42DsKeeu9mcR+h9/ZT537e4FF46W9hAtTzJ3Q3CEkS4A
CA/hWv0AMoix7KA8oumKbjOkTysBSPev3rBg6w/wRx/Zb6NOg2mxNAhoeiaZZ0vzoKkKedWksp+v
YjXD3K2M43UAZLkaR3zaT7EN+aRtCeg3m6NsG//Lz0VYxR8N0DP1rEjnaQBEjj34hxGSOvgzBZ5r
vDGXDGourORYRP7KBjmHlXtvII4L3tF8CHeZ4M02P5tKxorzQGwlRDJknWh+tJROHdU/0cZrJS0T
GA3+H+NPNpstQ4hYy22selyN62Fdw0IodrnOFnWskBym4lgcBY7TMO1uit/RGnsccM7cS0LIuK42
VKQEjz4mWMTgMzBZSuHQyfjY4PfLwk56cID+0MdMpfzIO2kebBFi0eVKpUjAwWOM2Hfno8ev9V1S
3/GNZwy1/CQgYeDqvu1XX1eUqrOD0ZYzNJvqjNPOzEYVILt4FnRLT/HUs7M3SJ2mJfvOBRQDZU4z
KnBbyiDdTsNHYK+MrlsZssTsfmxVnhUmNqGVpzzmHhB8/3/ZRhttR45PwjcMxa+q++QJmDsaa7Bm
A2qEg9eH8bXl9IoXqL/xTDLVmqJQR8fjgGB83i0OpPOFSgLTUEnErqySd/DYysXErG0cYEa0nn4K
Qa1F1MsUg3dX6Bh2IcU6++FSU42y+ctFVpjgo5+rHooMn2EE7WBXFyI264/aaMRGox2ejYQH2e1M
dKK8EbZmyUDsX1bCtA1QP5fDDWMyvJ5FXx7iamZGleddpZpov4QIAMT1UWKZlg6UpQmBcvBwUmLt
xkwsRDzyS/TA0yqHC6e4KgS0NkHmIhLx7Tlo2jI2gACsMdZnM+Tp8UAIdI5j6UFGfiVR7743eW4J
9SyfnoXWGfuEK7DZ3Lq0znvvuY3uvgpVn+oXM67NEfjWlWMFK6Id6BOUnZG2XWfufuGEIa0t8IXk
+31+jir5WKPBSHb/wsob1tJYMCks55xw0ZCr2e8GluOnaIt65BnDcfeEhhWM9dUJ9FWJCXAK9xfN
i7nyMLd4upQJ3zl0TdVTWZEt212Em7kfXVd+ErGQZqEWiTYee2C0eh3lm7+xHWMfV/xEdWBKWrLj
lJopN8MLiVuhpu8q1WanuN29ySfp33ySCVL547RbZc/QlBjyEpCv8f3rK2Cxz2GsPyHvqFe5Mb6A
dDvJTT3NxiaCgjDGBeGSMCDE2k8kwXoNXe6AquCUtuNg5rUgCbt5anVg8yaj5XpaZEZp9yJoBmtM
XAjrD9fqPeYSRJ9ier8779KOCQvNOanjTYth5zONQGZF517FHqifeYLSouhHLiLjjGEDUnT/Wgy8
0o8Bl9bMyg7QUVqo4D2/yCtdKcGzcx0uwDU9WqY/PoR03gdG8ueVWdOs3GsJpgyyyG9Xz7p4WYYr
sBp2P8PRj4dYjuoE0JTH3IRMf6wdhZGYu65GBhiGtW68a1VgYBk7fdHD3aPLzqjV0DQvLdkkEFW8
f/ZEKhES69W2/PsjEhLelNIfCUfBGWDOLrFvGnURbKQGz61sjMg8/jg7AbZDKrH5Jtlr6wizQNPM
W2MlrDkREOzETGJnukhoX21XIjDWXMWsy+yroB/DcUuj700Mi+7+0FZx9PEPaOCASIxn7j72Hpxg
TMfttAY1EmgLsSsWs8KAfcmJHycX0BrpB+PB2HcU/TX7yBRUUQOmfG+wboQ02qX2TWH2cyH0x6jr
xnqAoqvfiULhGhuCH8DKcLIzS1eBv+9LzJgBpT6CRrFduZwaam85HVPQet4cxAwGBJsH17QoO6t1
1YsmlORNODWnziVZeDe8uBWowL7nInJcz8U1l5SiBapsVSSsamZiLKcTM2/mNdlhs2ZB/Pj/45HY
LyQDDTcxmVy07RSXduDoJbiXZBB/utS3OGutFtPYO+6gzTUjM6VMuJ4I4o7EbNrx+EqYuSd6lA7E
KnrMULNUVbWtF/XGBkWPP9RSF7Yr0dQHcgikUNWt3W0XdGdx1O11IfUUT/xYp6hOiXDBJ+4PBl11
FtgDOasQ61v4iVtR9ustt6xiSSH5cO2PXSqsxwz0oWQss+Rppl8JT8KAu3bcLVNNOmVpiZY5wnxN
DMuisgHHwuOSbnZxKThNqR0KNywff1gbRuQRO2jyASGe+ToSM7z6rMxoUVHPz7S55CWXTn8sCY41
Oy/89+3lpbMNgJ2LkE07zvn/hpuHtHxG8VE6PIZkOJ1+XvyLOtc80auLqHbdhiHiMVV9bbHLlK7U
o4QMEhAKASrNnyyAbcmkejWg3TowY2TSjcVyfOUdQyvRTYfcF7K9Tv5kRhX+/oBvkzX4wk13kAXX
eS6tqRThrb+Rx07mIk8zmq7Pn5WbUad+AyndDR8uy+im9Y0S1wcEivrgsn+sK2BhRJyo9XxxvGCN
phDCQMRjWFQiS9sHmgDyORRy/4F4J9ByzurCaURezaZiwRnJ7bQtniBNML6tAbXohFEs8+fFw0ot
XlqBEUbMW5WMVMxCKl2o8vO93LAXDHpXtcXPprOmmtPN5t0uO35brxs7VxRFlBTe6RIS4y4WBWLd
93aKZFwfgq2VVBHu54NVlMU8veKH+Y0goJNuDWUC90Wyet1jY8O383do8RiisJgVSbVNi7viaCDl
+gRNHzqdEDYjbUXQqFg3RKjIRfX6x3nN73W+qg0HcvhjBT1TQv7N4WDtw5qe16TNqRUVRHpLsVOJ
FA8Z5nGat5deuOTd7I6DaLkZNh50FWL5tg44DRqICvDrOMz8taMjAUmrTCMl+b0vkmbVxvSrmnz5
/5oMhYpB0joAsyH7Rp7NNoHptdtrnAoWa8TrKH2QfTQ76lUo2YAAsCeOZPOTBcCQ21QcrCC2aDKG
uNxcNY+yvJZ1ORovCf8U07BL7l2GE/99CD+WttgFJOxvnAON7JajxYfx9mU6oRV0IbZpcmyZ0NuC
W6NwFGQpgbSfu0Z4onjlud8gp8ggZsxrTli0Z8W741JARKutFTLVMwVwB7dPqXk55hT+6sip+dep
z0EEyJRD8s/XkX+nLFq8F46Kqt7qkm55DrqTfV5oV5BUYPZ+C5MqsnGgJ9EKgMdF/qCIU3l5qf9N
0HjgOibAF/cXI0tBqKIrniYtDCwMwDnMuOvNeadd751VDFOZ2/xts7tl8zqs5M9Fkih7iui9c6ai
tlrY32YjViDNagyFqMgZ5dSZImQhVYQXiqp5V39Lh0+wGfbhTyHWNValoaXiptxL2WP5AXKV8pPP
ImIrHfO7/hLSpvb6X1ZU1hRVYd2nZGWzatGAqb2hc/DFI4nTFFCyVJv14nWqN8H1GVx3hH5vJH4k
QB2Vhyhl72YwBh5YuGdNiekIY/DF+wqhowlWzpl1gf8h6eFxp3Db24BYPrDVuBvuzjlBRa2rBnz1
vugTe/71ykVsOvnPQLPwF4q02wlQMtTpUFkLcxLcoOQSV11JNgro4cphkPVF8vyB1Vk5luZJ6qZ/
3rzXNUkoprhwBrPOyVVTuVDVRfixvu/tWgfW1zNDKq2rem9leQKJ5SdMnqq0Nukyx4cx30IYJKIk
VZ5J9yFSLkaxe2xFKuq826FIYW9DnC07RhQH3cfaIji/ne3xNRrYuuWQYxn8cNOLsFdNk/cZMNvP
j5H5ns+DVCcoM604gJXdnSk3/GXIjPDr7g9ZTE4qE6WaHLGXfMM6Z9yF+6ndBHZOfT3ogGgQyIXS
6ooSnACw4Axz4FmlWuCU6aB21Kx+Lobpk6NhmoMNTmT7s6vflrS/gf2Pn8102WnBqA5bj/75sJUK
/vKQfcJYgFI89nrC8PBcR/P4Xpkv5PYZo1E3OyIwQuOwK5COJhZOnCEeCT+tcpg4laJOTvf/BIT6
5cqsf6Y1WgSyxKTeBibYIB9LrzyI8HvMT1QrNd1GahYa2UYWudbPGt/UAU/dyG7o7JmK+H/8Z7cV
wH/C03Bt5ZDLUUBsZPpqBV/ekn5qXYew1+EnSqsexYTqHv7NXAzf+YezmLnYzq3GL3FkZH+zpitE
PVwKkdxtfr4mS4angOfbYBUG1gXSZnNnG8URC7CfRM1TzwfV8rKJ7YpC1TpcGCagVg1EJoNpg38v
odtCKdJqW1Tf0efx2Seyq8b8ANjOPZy3tCSMGsF74v+d67+11OMjHQmjmPfo4fYT84ljSj8cYHH2
HMkTk21dK656874IWfL+f8ZVj5jdW1Pk88+bvwLWC/T99zm3qRJz/WDmXFk33AG3I2Rte9IsJf64
1iLYVB+K0Yfto/JXMWHA9qI8YsNDhSpZ17b38hBLSW8cHjV3SlV9hSWeWkPmucVaET5JY1sbbq8g
JtgH/2OwjQvFNFo/vsdEsVDHASo/ShsIRoNrxKKu6IMk5EHGeOpyvH5JMFFsq2Lhf1ZxG93bEQSM
DPpnJL1QYSKA4YMuKU6GCecOIsu2AzEIFLSCb8/1Zy69n7zppczDvPiTzGY3aKOj30uiki4ZndQZ
mKbG7M3elo+EOeoHnqlKwpIZ2BgH7SMZaTv7uXDpIzU3iK5S9ETfxnMIe/u1EMaOhxam9RrJ9iHz
nRxyU4aVxsx0C3ttcv7cqpgMRAhQeWTIU4A/TPQSVIU1iAVptJBy3zbawTvNjCrNYENIm/xjIvWc
uQUQ6f/X6o6c756UswiYgWFJJnhUNhwfPu6KRMddvP3X0/bBxKkiDVdsi/7pM36J/IWo1/XiV6CX
HTZ8hFtq8GqBO57z/tEuX99uJkx4zEinvMqGKLQ/WcJsLHPoEbbkfZGfWBpXXSUJUQr2slJdqIKy
myhBOhccCZ0GM6s6TN+JX5a2I22Bp8WcCJ9biJxnIf2rnfQ3WUUAUrLqAEy/rCHLbU9Ia7m83j3W
J2xiNRhP3HZYMC2nWcz2iKajOJAtR1ogPIaiYSYsDf00wiYHJy0YdajjHSvzXda0IA7cgee0GRKG
9FafNABXhDsuTIZ9tTuqCPui+qOTn110N88RzPrDxM7ZKKF9JQrimsmWB1M1SAuwBVnJiL2pQvwa
T92cpD7k7xuDAM70NNNb5SrfAN9Fqron82t912OFk1bbcQ1nCCbgalS0iPiWqT9lPsKpMUeZb81C
mQEMl8JIuTrUWRbtdJLZwnGBttCfRFZryHqS9eRuaP55D3dlauhoKTQ35B8z5+qfUmqlCp9O66PH
v7b7Np0y0f+9HHPC9pFCx4/TGDVSNiG+Fn75k5DY38p8npQGc7+ukHZzoboryBac6Yi9N806gIlO
ptGkMVldqYmRgvtkGGZw3m+30APlzE/Ra9XMcsfPePKmZFbyCZeapqF7vB7a+NG3wsLxskuA5OK2
x3WZrfSnkXMT6zjZWy+j7qPPzZ6zVaYbeZuRZ/zGcmJ220NSAQ2Hg+U+HKnDc6zpVzaHdY1vfE4J
NtoxZX0PoXRErhUIaNEFq62k9ym4zGR7CEhnWSS18nkipuW4KYxP9bKMhjdcEnvKtJ0XY2Ke7Zgl
hR4hAIhBelgjTSF0vMgovYkQ1t+sCWDu2xi5nl/eZtWvHpPsFOqU+qOmDLK6+QvLWWbpW9Qlpc3W
GVHfklu+cFGzZ1mXZxUy2hsWeEh5TpnIMeb5KQDaPhfKlWycfL7jUBSP8Y8D4kYB8wn49t9SPdSF
nx6ZvTXKlxDWcsIUltjN9tVzAlkGyIid2uCGp7eEBY9L7mXSZIRs3L/ktmag2cD53JlS0gysAZ6D
ZV57v5eNAbYrVEOR9vpqf8UIwjSCDwdBu7RRcn5s1KBAdHxnQIjVKyuPa8eSCQFVr6ztuFAE7jhh
PaxOVSaoGJr3J+YNTLktUxlTotZEfR/64xZbCYPit0Iv9/3OfypmkcK43ea0WEESIoJWv4hxuIu/
zPFRiiV5TN3G26ZPTC+uDMb1wegmTjDOq0vu1xipaUmP1ccmDq0cx4RnGak0T9+uBhurhbOVQv6I
Pt8psiefXUPz4vGbVkU1O40I6NB1Ai3pnfMw0nv7s04Y2zHRiHoHVt2l/3kN0sRvXsQuCoy7OV9q
sQeUlnmcH7Q3/F0IxCUacUKI/w2J7ZQqG51sVl9zNrEya5D3YS9ByXfkAFvY5q2zroVAkCU+v0Zp
DJlTHou3SNLJbFuj04apAqqXjAJq6KWLzzLOuTElae/BmchUsmQPwjyvUSS9WIeY731Ke4Y1T8nP
be/tEgXkIN97aJGshzTBjG1GiE1zDOO8TR7dECsEkRMpjkNofombJ8En5BU86PtWrDqasyghyCm6
b9TW2CrN88PUoSLmK2ujSqwdJZsC687igrLYQzbZQAsJu1OWuE9Z28IOEpMoEMqzehZLU0DwnzSx
tCXjpmU19xknXEmhXYvwf80iCu2SytSdOhcpYG9IWGfqmkx5dlmNOpQYbtuaNL6HLX9/kSpS1/5Q
GL3u6as6j7sJDdKGWiJhVXaqySQw5/p+2UkUSeXuwf30DPPtCeOXFv61QPZmuPi6GRh/Zgk2iMqO
9lCN9hNSznDwobTUG78r0/Kx3XV9+aJCca8DiYuAgdKQVqBZwMBOQeXAPLsq0oJh/x/BPoT08GSp
ETuZezQfnnBFrxr+dEzggue6kpOS9+luzzKjGD6x0xkVLz9G/xe4DpKy7BCZEj8YIs4rPC1VmkIA
BVxtJ2xHigdR/PvQR0BdmVMvdG25hJnhFE0xwyw+guW6s2cESGQKD3RA/eOOdSIltFqiHrHIn+xp
qDi/wD9tg9srU7eUUvSkMagGQAnNd1LD9HisrKPQiRB9HYnWOOBYQJj0Sl82QcLZY4wcggh3If3Q
OI4iJGS1qcXx+E0LgPsHOYefxbRGm6rVL7V3Fhm06M9w5B41KyHxAhQug3fO6hU1RaewyqIegqI+
wEXb7l2OGpx/jg8A40+CAAAkwtlHTY1sYe0qXCKbkUw7EgQfldxGmRHAFIQu2YL71CTh9qIvRWgj
gDCerHbbHXL5osBqBdgXdTXXjmKboel8Otmz2sclHu0TeKsE0PLImZI637jrPmpvE8xSZbVj+VAW
ncic6pSTswttET67BrbV76BoGNgpTyIJlEqpGDzo8MbfBaJtM36B8rYrLXgX1Q8sCpuQEqDTwDIa
6fuvitRicGMmRse8Tyy+aAav5ckrDo+dM6f3Z4pOf4GzJCrgqi53DyZUSLKa8Q8KO4OTwKYmYxOu
qF62j3ZMcOrIZoaXyzXsgat9D3++zOmqFZYDx46bfUH+KXLVY4hLzgqoK3Odx1FVzEyHcMwz0dID
LUw8vj4nAFr9OjGL33bDjgA7g+VKzpvQfVytgoY75PUFBv+8u5Md13a1wU5hejjPOedzI85gDc3D
INSIeiPzTGkjyZSR+hu3qlYvKYcAOd9xKngERGLPHiq7Mh7AGIk5GMzqsBKk05H29w9O1hl3ObKs
zXVJXem2FpOf0l9onw10F68qqvTNAEYVqemyF+TfMZOzlXnBGZkVj+UaVcgytr5XPUGRvoyAlih2
YS2xLH5pnnwHvKIihQ+ujUPX7xGJXDOEbFctphw2mUd1SeCtiYZu1qYCnsLM4ecp2MpxPfv/b6F4
KVhl4deQ3fyU1KTpncpRNiZM/UlwgeZ5h6aQx/Uf7qo9+CFtshACMl1Y4eUCe3l9yslZrA4IdlPm
XtBZ+Gi2feWVp2iP5QVD1DgassPUZjYe4UkScSbmOkrCNcAqnjw5F5SgTlLHEiaKtf9GwdRnJpgY
B/jZSu+qaYZ8Wr6NnS98kwhKczvrgA0CaObMcTP32GuoIA/GoCFaCCJzcQz4kbathYLEDhDMhav8
01l1iJ1bsa1WoseUFBWE0x3PoMTNxZjK67ztQJdkN1cwY/s3RXkgn6NVn3MM/Gc5zrRIht9BdJqx
KrhaiVszgrmC4A0dmUO1SmcQVjjSAXSPmziB67khXLpWor7dQ6X36AcWqRICxxliFSLBD0U6EinF
S+uZ8AjCL0yrPrugq/a/8zUHCdh1phAbEgckMVttZRng8guFdtG3UU/+T2Auw5mdtwrN6E8akDD4
5LY1nhdFDuBSbkz6L/JOWBxx/VnU6d/GCLraB1JEsv7Myyyw0ZIw4ctlRzTZHrBUg1ugf9PoBoAw
6Xyc7HvCg3Qq+GIyrRSiMXcLNFqS3TfGeNOBs/zONaBROOavHYUtMPooF8N3M4BWpjB4NGG56dmy
zhG9M13pOXzftsTJddpRcaozIcybeS4HlLdzozfBLmVIF05xVyf41Le1bKB299uhHoMzHwus7MHw
sN1/VYXMiXuJe8tYJvqq3YkZV3ZwFl+QjjJo3eIo6pKmbr06xgnH9penfYqNpBGqEzn5SwtkhOEu
0Mw+Sn5aq5klAy62UnqOfXo6rfJuqJ9nCalgjDSe9JpSvnw8PjLCHsxlJq0auKr+Pv4N24VF6u5o
O4fizga4o4DHz908MwmIkS5IeNd1EtgB8qmp/vdpbNf/AZT6K47LJazoaNelejdgzQ79PStUZELy
zopVIHzbwFf7Nww1A0n6wAPXp2fIxkzcyb/LZ5z8u1g8Wa1PyGp39W/UqGKsjtsdQ47je+ClFg/5
7syhQMURIQ2VjeUJ/hLTeK/gnTqTtppZc9jiv9Ny9eyNjkaw8tM+zBNO0KTFBNiWmcr7z0TxskHf
V1CE+cYJimTyBEhHTXvHhJHFt6LBdq1+Qi0VFNXJw3J2FMVBMtylHVpCqlwUWX0daJU3EP82k2ic
Yi/rgLKReHNj1Lpeq9nXGJypXqy0INSL4+zRqnKMX5psGPieUtKzeeuaI2vi1gzGQJ0AShD54PVX
awrD4eYZ/FZuYzSfzBuKPxr26tu+aOIdaMoqbukYwq10q9HmojJd+CUmiV4ymVE1TYevhozrm0WD
4L2hORxhLnapOJQsZJKbe+JcxBpBybUmtLT/mY7KAEeSYBarKWTxyXPXh8pkftcfZPeHnbbEEwsd
krIzU+JRAW8EwnxsuhPradXYu+KrwH0zIigJbSWn0FFGarDye8I6LkOBNFGouw0NOy3p3v5S9PCf
GZYv80vpLnt1yYBfYEpcHqpujFDcWIMdchTEtt2+LQIexWXK+XmshqJVvjv55tp6+IYFgSoEv2Dr
H7+fPrGM5CJy9d79NbQOElSFup+jGXW33dzJZVrQe08NnaKeg5BQWwq3YXR5dCC7lhMefjlnM6Vg
2aXN3h0WbZwUWxQTlskzhwOjMVzS9PxKOep4uD0YujCzsRwYbgXQEY2PWYJm/OgisOQIXzKWL/NP
JoV7hX+iAehbL82kTJlquPX50ZKJ6Jn/agh8a5QjfV0etn4m+VcmkeBSizq4FvF2Bm56JnUVaZbL
qcJVtpkDJucviVn5SxYGbtAQFV+wuwfV+oGKn11NnJPhD7yN+bRrJWNq176p32CKWKBdYfEn2kXL
rpfipATk6Zorbnsu0y9z0rfSM61BvSRVPNVMKW8Yb77e4Lk8ZeRY2tMhJOtguDtVtNL8GXes0Q7R
AkcYC99nbQC87APhJaDke7FDcNCtURm6w0u9SV20+U18hQBYxxSt6VfrG7Pxam3qTRUslD6iXlJR
TavAiWr0HIo+B5XD83xhVst9AahNjzIUDIWLGjmD6C60HGWQPxHzSdh0WVd4lvIN84o9F3DdhuHd
aaLvmxgwthvTNJWjeI9YfL949jFYumy8OIhsAoac5xgVP9ECPirc1L3WBlWQthfTJRqbFqws5dwj
RcxdfXhlRaNdn67sQDimv4IswJzJVrjB7EnGYgqYFWxXNi9X3T1K6WpXqTnDMiYxa/r2ibebffiH
9dgIIT++BaIj4L6Ib7a3QB2kr3nb5JDv2mHHPSFR3UVfeZqke2tBO6VVlFjDkxHc7Lv6PN2fXoDc
VuWoManJUVYsga/SbSqopR0Jb/LZjoWcKnW9l9H/xXAtzYDCYiw0THzktHzSojEKAnDAM2MG0S4t
RYUfGgU/w7B8FVidbKkoyECOBZwvysFW/uStSPPjJWrlTgb//w1TR9+HNSb+Z64uLvYCBJZCfst8
JjuWXoVdaVuQO5+0Fae05vCH/kXjX0hohVm7VfRpSoHlcVVb4QrEhlnaa8696dWMT8qimWa+IWB9
dGts/CimWxXRmDTCIc6bpoOaOxzjKfZjl14C58udns9qYeMCD5d3k735+HHGDjs1A6IYEsN65sip
3gkJ5EnVqvhhQ732khUrvHa7Uc19avkjIto+QUIjE469Z3E56RWbA607k4R8uyRJemZzRjQbXdTR
8YuhZtZGqs6cmUFtZAApZSXzpyAw1WJOfWto5/zhMoloMn7TLfi0UeDl8lYvN58rfPB7cmvcAUFh
pFuJ1Ua69WIw2v0Jw9shFNwC1kanAIMZvmFHYk/evNfK245mfefks8Me6R9QFyzRIdrv/NDZ2FDu
i8sDAqYxc0gga5FQO00Su2Y8B4JJ0/2R7QMgGyfZSIRemq9ATMJ5hzZMRaxoeFLHtE5stpWSvktq
24RgO+aTpoNjjYRHwYNRL3gTI8dWGgk7Maf/ebhDvz0Qtxxx4qk7WQf27l23Eq49XNeKgikYnmh9
oiH705coPO/qXXatBYt7zXMy+JR7TeHnwiVaklf7Gc02sdEARcXw0XLWN6hDTYS0fpk8X41GuOiN
vg0iqsuc8ZJwgDaFZkVZRB+XimExbWKQ+Vh2MyiX3dYcPBQY9lvEwQiCZ34eZiHVn0ioSKZn/MlI
5fCgn1tOEMQnW0QnIbk4Ei67RT4wTKG/LM9y9lgXOm1qEwX321PtmcsewbLl5i1Fr0IszntpBxoy
mdtnlJjvBbCK9NziBxMfWXfzsXaM2OqbqfDZQnOWSKF6u7t0h/H7DZQHaNAlvE4Hvl4bLQqQ4aXP
NCFpxhpfIyI9Y74rtJv/NLLybXwivNXno/2i7pCof+dPibn9s78Uxqg7JoP9fQeRs6KP6b+cBiSd
yFvcj0WU/aN9OiCfAzgCIprRGnb4Vw1NU7hodA63pjcQolxMRw6O2dT1+zihq+A0mGPdqXMAye7Q
0ArKTMVmJwmcCbVMGqBfwud3UXx9jDHqbccaqBCishWpNfwiLLFkMGipPRk89XGcxhYMk/GL6V6E
mThgAd8kJaqOHrUGJZNw9iIDHR/ejh9YuB394eLiO2yN9CRtTlIghYaojMXK855q7IBI4lOMiinm
33rRdvdRRNKUzB02+WkKgIq3GfVRpDcBUdlI8y+T/Hy4YFz9o2i5gR1w+XsoyN8CJRkt6yoNX0Mf
re6YfiuhI+vvKQF5mxAvAHXR3taPVKMU+xVxYmorh1g5ax1ljn19Rz9CbEpugsRu3XD5kFiGYWKl
76g3SnYD+jGq6L/QTsY5ZmooGkYTVc2MkyzlabiYGFb/OaQryfL/RWKj7bSfJfCf3N73sTbOFGOc
E0OwLR/onO/cejnqCtWan2p4uK0v+pg2QATGCHlGWZshfG9lS0K7igTC99h1/gQf4pvc0VPgW3R8
gU33//5o440Yigv5zP53g7gsoxJsCUx0f4xmXKunfrYVBoruv/9Ug69/EwFOdwxK3N2evQ3eWsMp
eQmKAnK/Tn4k0TBN/ACngkOMZSJPRKtF8YQn0lAZuWXaTdTcipvPXWKyzB658kRQYEmIDaw/bYMv
Zt3K/A9BDSKJkI4e4AGlGEDrs4bT8/x4xJXKUOlgcnheDsk11o6qF33k7Fkf+yXlvlreFWKhar32
rzhrBr34jkrwmCC2vEB48mHxLaRLI7MzsuSNE7gZC9ZH/nYeVLGCoC2Sf+2wSbdNbvsUXnUCdhYv
NOC9CHS6pWMMEiUyHbITLTS/DAtecsfMnKLbPuJkrUF4H4BD1rOFx9jyaTduJOd75Wg0QOSWbd+6
WZ2/8Sj6tfUMXiIriBPLZHus4WQd/yBhYmkEMGGLAY0trInroP9Qdhm+DcOWHLfOx089rbX5tn7F
lvTM/5EGpycv/lkrfRXhk9jcws4gadMyf78Czda3/puu5lLC84Et07YLYkjTzQQtexGiYJ46FklE
jTc/ix8tGYxMRQ1uTjejCbe7DzTMoECu9An7HApl3LoemfilD4j8icZVyTTe+yjJXpQp914+xvtv
LTMRNChPrzef9W18nfZlp3uTzQuufc2LZ9ulySB9Aiy9ZZhpJWuZa+VQHT7zxhjAufdUetx7UCfW
/gnuNluBceGnl7wDE4HTFvO71kag3iTLTnQ2XLGnhggHnLA4nU63GyLODZ7KRO6K3bCWkRA7TgIn
hjLmsFb2EO1ThUBqvmIl/Vcyq9TgiCxa5o1komxn19PbrktWJFq7RY9gHO0kg9iVa8i4yMcfNIG+
eZSXzFHlPEeFQulj2Ti5r4ed8QEyteehLLedmvzjCQdBp2QqiFT+Hr5VhKHnunbyJqoNuCKCg9Oo
wa2OuwfrGPvsQo0iHQ7mTf63OOYcKSF0Ut8LjxHwEsLfBIiKMhtN9P91qRr8s/PQkC5gXek4epns
l46hK9aZW/WE4c3TlIMnN0TtzfQRNIZ6JUJtdOM6KPXNLVeRHl0a2+6omQxZPWSEE1/pYYHYtjYF
E7uY3Hh+AQ8zlhmoezBV2S9X4TVKomfH6FfCnp+CQ7P+PlboVQ9DHyKOrJ4qvlYObj+uzGzARUwz
HrCzkl387HIinFndfMAbrh1Ebb10b7E05oupNWaRce295+4XLat2VUa8EyuMA8/qgWYsLFKByZXm
yI/QnGcyH25DYCem1FSmynXR9yEvqJnYWlgpDLOB7/HsViUHqveVFc0VaUMcxr2dFEUZhdBLQLcR
wOu7kphQJROnyT8xzWl1BgXCrABjSI0MFuM7O3MtU+kpuwZMejx2Ph4K3yhX8sUkNohkm6T101Wj
qtZBku55DPr7UyVwaI7HjQAsXk8uZWaKKGrBDQ6Mp9rZR3Im/+NGsxodePndpgaMipJr0Rz8qedH
IuCZ5rMc6XPJv0XfIaCMaXK2oPQ8ON8HWS6y0aI/eEj1QbmDAKsN6eHiAP8aZ9JM9QyKWIyc/uqv
gQtzegoD9MnA+j+g0/rImSZ0Nbic5DACoq+GbLTdMqn3ZdOuGE0Y6CJnBjZVlc2S7snc7eCx297K
ns/0oD43pStPTk/ST837YLLkrVDgTRnxuNVE+u7lmw3Ig5Zd0W9YSNo9B8Ob21RATYo4FPfIo+kv
XEVWXm845eBv7w5vAdhZhfs1hh+IG4vEbSRLQey0YaYOhPr0UMdqXxyb6ZBufhCgkhTGfRHiYb80
sDP54FIrM94xIvOTS/zNI5EfT1NS/9kAdByUI+3JJ2fpN8NrGC2ccgOpVGAX/2lZluubcxHddhtU
cOR445fEnzkyZJIRdqCbMi+KwfhN1FAHKUudvPhOtGQhnrEggkhwL/GXTrn0nuEykbHV4XOsU6r/
o6teKF7hyTHhxc8yB6iiNR/674kIjG3R7ZBIo05h7AKZ8caOzprdjfr0rA8NOJNt6TfuDO7t6Jur
glOTAot4i1Obeg28JUArgrQdQwcLrlXE1/1kpAMnEgPxU6+QZRLWU4tsELvFrgwdsoHS7TFIGYS8
sjGO8L7tnzK5ssITNNWgE1YWj6oVA0qgJv3dfKoTUtmxX2NhEY+HP2zWbXqQ/ZBxyczklatP9K4v
BjLZ+Xd9LJ3EvgXOlFfmjhgNmZ+xusjbR/IJJ2rgiXUVvpms52XGK49B/UYxZqg/oCIg+fTijgNG
y1Gpnc0P7HeFo4vsorFTD8rV0ZSZz9IKHTK+SzZ3tYroxFvrqQecbVBJ8qnDLk8C4OkFGBS9PTb4
gwdxM27GfkhsbAQes8SYRhHN6xjXTiHnQzbYugDAlIcJMW/MFb0OjRQeaHDf6foeKhT0i1YaE/dM
Wb3vHnFaUlRf9fp2LO6kAR7Y7//AyIWu4H2zpi0bLe5gVJQ8w8Uzfg9F1nKDr+YfvO5H1X7dDcHN
Jdh5MiH5abI2KW/i6V7BnwxlBD4zCVNofhEo/Z9nTPI+1Mi2WdtNwYqBpmfblyhoBq9lFoU4Dgjg
sTQMdo+XNCk++jOZw1dFRewIjARjxHhQQn0BLQlBjSxIJmiG5RGcHLhMu+sSydSN7mIRFxnfOr/s
fU4UmZF6PJU20Whv/q2qjnTPYIWQMuawtSJk9ji07bW9s51f2wknKOG3TcbWxLYzyq1bEfre4BtJ
rZ0/yM/OrC0TSA9y4aYPx0CRXLBl6f+aS9WhYi9frOx3bcn+Jd/pg8XobuAQPWHz8jevbnnR0+3I
kB8v9w0EsXNgegw6lCMdqFgQfbj5iGkVhiuPY0YSf8nppeAv1TlxxpXaW/oU8nBB7Wh1JMaX/uAx
xG8Jes9pfZPe6D8+3dsilWVzRB+XDydTo3JDbdtMs5ziOQTgM33rY3hUPM4Idr4wIHVA4Idfqjl9
dA/iBHg8lfAH67FtQpqBkA9lhDuNyAOSXVNdQ3IoiVl5KUJWVHfhQNPnQcwUYIzdtIiw2Obgol2S
KpFvHbbeApqnY/bPy6RaBTHgzgip+jQQ0Tw99EgZ7/O2SdsdAx7kUE8PEzOizuQ8RHEKTqo9kTIW
0hzY84YqULS7sy4aZhPaeDV126wqEMRGq9wvXJWsDXJQGH+pRQ51LtLuV4oKcPpcJVLxa2anLs7z
qo1IbFmWUfvHS1w3exkkfSSn9J4mWSTmZiEppF5PGXBvher6GXiynLbya4IGHAYKmWGmFavrc7Ng
ncHhoyDEMHgiHIGaklUQS2ikxr0M5VhwxnYsKDA7ZrnkedRBufAKjCK9F46AYcEZ7zh2dnAjpe3b
B+CVUyVaDFC9mJfGMkyOM8zW9P8xzuElsXITK/kt+sPJ9YIowwjD0kBa3KznQYDioOupj+QtawaF
5sY86txaUa/Xa5RVuZNjvVwYJ6p5D49FssAV0SeMHUBLO5fXfKaQMqUnJNbi6cc2IBOuT20PW1IG
Nvb42qbaGtO37q9cwZXLD8UhKtDKB4sDrk4DkP5LizuauzVfmHLXpi+UIue7xuTmSgFOBumGe0MW
mnapVYCpCKCqvhk93KcZxs/J0zVTETaHBK4T8bMU0OrsxcgwcDtna3+rM5PUC3hTO8wXU0l4beCb
padOjfAh2tyjToqjNPZVCeO9SiGVtAGeSMYXzueUIgiwiXb2K8jYPT5ccwYpDQBklQnDNVkjKL7X
5rW8xyYUjmH37JSb2eTx4/letN+t6JmaBDmWLFzBCUx2Fg8+W47/8uSePNpB5vHcUOk8n07CnbvF
K4WhLukDPDNMZAsAgrzYjhiRp72O/RuSGxjcft/pthEHHS/6sm9HS2BO7l20Wc4upPeVB2xhOaQi
TLahTikPR5czWWpuHixn0+SsMcTHD6KZE7c556JMW7sgSO9dkA+BJSTtEwUpYYmLo/viX0o4/cW+
pZK9uI7k/ixXgPjKg3uvl4Ged3Pq256tzqilLmYhl9bBjhwWMG69Vrd5JPwkkn65VkPtt8c1JMwF
4uy/oF+ZJxLNIUBpVP9fDIq+EO4sV8nvQ4GQInZJLH0cRneO+tc0gSDl+aAqdEK4PsB+4LsQiFlE
1pW4AwLch3nWZxgYkVYaMUEL0uHsomrtr4kuLz1LHtoEhF87c8PYif9wy38wW2sEht3IfH8Q5nq3
ZAZwQCRr6Mpijxqpaz8IjKqX9j4nAaAGX3hDy29W//teogSsBqel9rGyulmKdooO5fWEqaszNQlv
WJRIuqLBgCfiwg47IPvGMrmcDCzowXeERs7gqLrz/dSynrXRtXNs7Cdx23mgIZv7eoSn4/DgKvPV
KrhkkzTyph1UecHc8BvWpXvAdltTLIg9Vr5UcR+vzIo2hemzog/vbuALDWn8ItNRIRTfNh23TjO1
TbTddV3f7amEupsqGnEXmWICW7hEPdHzCkHkx9QL7vax3m0nCCs0YSMeNVqcLMZ6phU5KuTy2cSh
cbJm4Yp2SyPuUg4jmiIyPn4eh7iWBjql2d76y7aZICUPo/HanWrOhwoOVmN9UOBv8AAN89Nc1R0l
c9p8fR96fdMqxa/OaM4cGaRqwoPqJDywud/1SW/+du+5uXtzNjEXHtjz41z5es/qbnrRzOQlMhO4
knjv4LeulHcAo/1fH0Vt2AIjAVwGxp+o1f95G6zAWptPBG8tklLTwFZTgsJE1x8BgzxUiGfVbiOo
MbM/y+CFr6j5DWke6D/kCBSsN4iefCPOU2YIhytbdQFTKCqYxH+vk0+rlIYAMZ/7ZDEEGAQjT7vd
bgmdJ4Y/df5XrzfFZELiSu4kAuJcxVWnz95m6XBKSByWIqjf7SiBNXhmNRTc0SWiVId6zkTwS2p8
6HpDWC+sWKExvCWDqasoFeh6DOs//41XIeZHn3QA8JEQ0BFDhxndixWBrSv8ZqA7G9M1xACTVHUf
vagD6nRmRRc5J/7xqVVkrw30VtAqXjb/E6wZI7gaHvptNV0OwZaH7sXsnl7Lxn8zA+24j6Io+zUO
sJ4SgTYPgK4urigoJkJ+TGykew08494Objc01JI9ZLODuqBkq8YV2dGI51xhks6WqiDU4v/5mVEM
hMF/IT76G6ioXflhhuL3ETZ6Sm4xU0n98cIqAVJxmussVuS0iKYSHN7e7k+YHlejaQ5ObNxUInAG
IKqGO5QrvgCuv5UxONZQrS8O4kuiCetjL+r/Wbdr942sbT7yqvAqj5BKbQA2bv6+9YzHVXNshgXE
Do5/MnnLss9eBnhbDMGjtUuBgous5HrgRFAloo2bijPYSZFT6Q6tiKqEyReY2lYT3Q4CZ+qa4KSD
3UutQQRge8WdG1dtGMfmUewpOoUBWqxiG4xudL5MsyzKZy3wZ57e8Nxfa8hDGKjNdJVmc/efkqGk
mkvUHm2lxKoA16m9ffDmIpWZJ6wijt7HXD549x8G/ZmK9KbbDQiojcrw0BAxJx14I811FOARlMcK
RSDXtZZdPBa3j/ZPVZLXVY2KILiUVKtLBZ30IFHTEnMEgFdH9KgGTOJlZUtnNnqhSBoX9h+s79zP
6RszqR+ZTVhaqqKrBvb2fiM+//zotEf5d3Ur5z1C/XXriXbfUa9k8tRJ0mMIQpQIVu1p4q+JVZtb
SZOYpfY6sJjuvxdPjjLo8SpwC5+9gje6UYfsO1WPmxgxTkrD2p9fVhaor0jCWjpHEyHvQ1pSb7TH
M8X07Jdzl83xmF/qK7vvKULtSjmOFgCyE3yTjaB3SRwaQ0QFOF1ja75NtGZBme+KEWpXeTzNbrzU
BOwrraXe7AHcLEPE1x1zNN0q1mq7DwsHPMJ1YQi2whuUHA15yXO3fadu51FBVO1Q+Lbnp57SxPZQ
zv4P8Sqjfv9mnq0a3HOpCnUirjDb+iQE9tkC2cetUdvCOVckE9hspwacyoRm+KjxcJ1vFlZbrT7T
RMlPQ67Oi/Eek6moWI4Gg8y93dUoeWoSThKk6WchSe3SKX7buyoihZhhnHQcTduKkxBSQRTivFIF
3pUQZYIn4B6zDTHXtQvxHUSwz+Y9Jeq3fN/6vJQw1QyciprvT4RFtWogB8hD6MHTup8v52z84ylC
doBog0/qavqdWeBS+27dYV/jrcSzsom8/YXzxqk3li976WEw21m+tfCgBouHRMUkN9kdhOCWit3K
nhiCCOnZPlEdMsyWohGbTPTa/RnpNRVc/jGjkQb8+j4NyFp6lpuUHuO2zU5mw1FowsfsVzZCh6qb
eNEPpGlz2GP0fWeNfzjjWU+Smmyt/ySvmZm7My4rU6+XIxJjgMyjx2b587fuxHaAt9bYUNEsNx0B
9MZLn8wJGsL3rLMttAb0ARzmwc6uydXnW+IFO8cnjCM/R+vygkx19VYUWB6H3OTtKYMwTHKcwi4t
ZBCzeCB31QXRj9Vp9DLGotDy+cLsWAyNTeBxEM8ycVvbpNZD0jKOtNZPYA9hgLdouN8DKNZH3YZg
/vvcYegpTAouOxK6QSHTcFi/1FkWf8ng0m6q2bh26FTKxWJtdnbNbo2POd6DvkWweqUZqdz9gzy+
q1qZ95VdQqSTfh3aLXtWTJICsmV4BrcKS8Z6YihqWnQtBZ6DFyyW2Y5vkjAKmAxqh7kS1+kQGDdh
2f5OoPJbPNezzYMC6Q6TiIObi28MieFq2OWlP4eKqVvE8oy8XvM9kbFGA4KAg4PcbE7IY7XEO6MX
pZLHhXxyGrNDc+Eb7ZMThtB0JOw1Ke5snL5frNudL19zPruRyrIsBiJgSTeFMsfiwvvyIyKWwYCb
uHl8CAEuzyBkn/jm5FVDbvuYHkSp3thG8FZLe2JLogURRXVZoVhzKmNb3Nl4X9aL7qQOzMN2YNuS
0x06xy67Kic68R1xwUyGOxB1lJTUnyCcO8H+rHVo4RrEyLv1MhepBtkFCb4JF9ubPL8xyu1PiNkL
fQwrf30htvkaLdDOrSVZXT3tnVjAEMUnnJpenLx0NCKSMkf16c+ZrLlgi1CCXjfGd4vfDmUCaLZ+
ZHGLI6SHGZT9kLvR5WyZ7sLCQFItxMUueIIHuEaadpzn7n3xDQyFGa1/27F34LHGfAOK4EY4vfj7
hWDXNcpfDgzKOoGRVIe0dOtVGfDlA5QoJvaJNfCOrQZreRNKWgczam6OP/s4OXZz9lPnseTl/A23
sQ1pJxIrgM3gVmeo2tRtovqwgGr7qmLe6/6JmynLrndBPAmNximZE4yFuAWBjYNs/b95+Fm1zojX
W9Yk2//MHJAK6/LBRvUsiAZElAdOWh06FHd/Gk3auqpwqpCBN+XH9f2akMnI3ldgcn+BiU2pRC8C
Ua+giYS43ASc7r4lFQn+a7UzEFSLHAHi1x/T4MiDGLM1T0Zl1yUBlEsXkqCuG0A/Ux3qC/a2dtHL
pdMigny4se3yW6+K75PJwFzAqEHPTfzq96AsKoe1WvIN9aggtezluCy0LCYkzOpuSPJJwzL3I8wd
axXwnxVvIcbVq4cluGk/f/gPV1MIiFe2gVRtmhNnwB5CWs5C8wqt396tshSZCQW3+IFg91E+3Zc/
LVAkvXAaJI4yu/DKqI9bvW0wKLNgFF3NtQ42pAnc0CBxH6olVOIkJqv71HdXA/qI1CylYJia7fRS
dj0bUyMYUJ2NhYRRWPFNWXxc4rwe/S7+Z2dl5yDqlLtbfzMV4K34V8pK301EciDeP44p0+V3Zis4
+9xF3GJkgErta6YCbxODzga/Bp7Kks7lHNi7bDnukVaD1PZkdbnJ104OU5DaYnPVWEDOM4jbdhD3
Asu4o8UYwoNtfxIPim4EsCrJGb+1w2eMIPucAcVPpnqplkoN8v0WmPoQx0gDfp+QmM9IKpP4BMUi
36VkygDH7+EmqY4GPWjmYKrBGdyQPoKv8nMNizysLbERgHdPMtbvi4TWHVoHHTX9pXD6hBm/p1x5
nlGogPwJ6tc/1fRBS5O6G/8MVG3OUqkzSdNpb2x4+xnl+M0EBN+3Bydd+fgEyOziznep3zHJynS/
1Vpl1OjGG2NxlYTTOs/Ctm0756BmIV/hHXJV5g0qT+EfkQ8YSs+HvfGqHLXdT4ANBUHEx7+6KC+L
3vy1rKMaK/Rz6fXzIkwnJmeJrvTKRC+I7NEpK4jMK9AKA5l1vg57I9goDZFF+lV/OdnxZwlvvZQH
8hwjQ7INno7wxUUuhpxKcwUFQMD77jRGo+FSpqwM2iftWLHbiCsgyhcd94Gx3S5UyLfheOaIpiQ4
DfuxGOD6niqhm3/ZxZmpdjJb8uYssAaFc8iFmPjerip1sBeCL80QoD8FVSBjjSoTzgRApmB3X6ja
wPQxmYUL67Upp3iNR1Va3PzfzJawKQozNjvmErXXdt5ah7d9ICN+hnxAAcFMg4Mnk17vFbAhC2Kn
IN8vb0xcUgxvODvFGLsJMR5ycJqii9+4Lj193/Qxfac0swD1ybtinCWaljdX7FN5v7qpG286FjMj
a8dYCx/zduSqgrxYmP4QjlPaGYR9MBROcBzpme8qeJfqZKWWb6PDUJahDUMjJNO90QQy3N2t8Nfp
GLr2/ZM6mLFSpjT/YPWDT6nTKSUfwcjyeEhXFfGL4YCblVDcZE3WIZazOiaifpHlcxr92xBoOdKf
kzUXXagzcWTmkE0riSbp/smm8wVYmEE4UqCuIhOHg329qRwiSOxRwj++FltJZvuflUEWWgvAcUTS
hZOR85E9Jtv0Na/f1fWfRFsVocd274Qg7kvKzvhgF/poN5hrywohTCXnPEg77jq8redjg7uyjqMG
8YkdF/FzXblLKWWn8a6eA+G4uZLZkT83DWQMKF/QSe0xhwlU9Jr4VBoWWMFltX3lgptPk3YZegAP
SYEUYxtXOMfltzO9JWyjNBvTcsaBkU9OvBc5ARHUWhxjJL28MrdefN0T83cvaLrCQlWamySFY1oi
/WqmvZcr6QA5kKGrRFizrV1/ViRqsWCejGeP8314TetW7YAIWw8TdomAoggGQIbatsbhSCQMlp/o
/dxKIkUqwby56SpZd+ZOXzYtJhLWx3v79DoFGHhifkvLXaOksVnCNz/qJPGrpgm2+AjzUPKS2Rwz
TMq36JOqku2clOA6AbCnnXbQsBdUODQb5SQK1+JGzIwykfc/4LqH5DCrGrYr5JuTLRUnD3eujcgA
k/bNfrE5bpYG5K6tlFoth8jnvhphTV3X7Kv1e0GVKUOxaVZswv190ZvrnaMA5QpnNtMVKlaBk16u
DgpCGX+9BkICmbjL7SbbvmaOLTr+WJu1JiMmm8uwhNnpCN1ujZ5lTwY74YgyvecKwNe03eXIa13s
9NR+iRu3ZxSadNCR3wqxTLLm1rYkJqdWGXIia/MLEwWxfbWMcZSkrv8h2hYQjtA/866w+NSZ+JQJ
CFB5VOJmKVIGHRxA0PtpXwaJa00E98AdB2QY+qCaAXrONR4VNulkqxeEPJAvUezZ8MjjjSNQwsf+
Of9oatmHGJeH7QPqoqMC6Fgf1jx2YaGhnA9Y91MAYcpfQGH0PbsJ1RQoBpunbicI+Ftb7CXAiNR7
bTsaCfp5eWFVjsCwAQbnl91YVORnu70Wimxr4iiLnhsVMY5SKuZjF6AZJi44w/ncNttv8c9qRkP1
sxCZC94i9WvJEC9/n23oJpRVY9Z8AxRi7/qg96O1WhIJVe+O3aJBCVtwbJNfGnZnbllqRB/8s8ql
rwYZGZBdYTIOA0AFqKal2ozSsOqghFudTIQl/J6ncEDY6AGG/fxdCCl7jUhSoub+VF4tE4BicC5v
3Jd4x6O7gY9Rcjt+A/owMGucZ02vfPQmeDTUaG732AB452mGb8HKzLspUmZj0q/RUz0uxTp3Z99K
pPlUS0O+roA5tWUATZilgY7ytYBMOJskMXr/TpgU0f/yjrublBA7EkgtXGy5uMdjQQwMkO7sv2v2
Z7nmFI0QgnXSpINscUEU8FdwlqujHDma46PYNe3DqpNesDg33owMWTbr8GqMG7G+QA7/r4+WY3dz
PKWcZG62uc34ybAKKXDKYf00fS6JHETM1GdDblKRtMsqFGzd8LyffeJLFemUxPGwoecYJkeIgaEm
vYgHzhaIHS/vSqiih9NIEJ8BfWS3kbq73BN8pc75oDzh2s0+LmrxbXl1T0UJ3BhCgU7PFXjnajI1
ivyHxR9/moJ91vBvksMDjjID/fgsKOFtzn6aOQdO5LQLl9cMnX8PjCTUdqM+2KwQaKt7b1vXcpyx
VarPH8+KwRFT6Ad7YejS33hHTAtweiuTXtyPDtSm/jsTd1yfju1zlwW2Ck1O7MA9e2tuqNOGV4z2
Z1wtRKqJvIkE39J9sLzYEZWxWCMmIPAW0T1wE26lI9qkZ/bL9jLnRD1nPHsIgLL0GJb6xTygzBSA
ye5u9cX2gA/G6lbNCpxj3YlSnFixbf4nX/Td3Iw1ia0MkuI82w7jDF7KrA7GNoGIpZ6vPYhpNQL6
Z5vgtt+Np2djS+vxXFQHDaagIYSPZNharAObDNf18j9J+lRGDfR4XMhLzQO1Xf4HrAjzS/Rd9c81
LtWGPNyOLwOPf07I85Dp2gvLhuOtUZIYLKqBNl/YiSDjJQ1t2f3wncidgLexo3Q7CsbhnvqDaNgx
j4em3CBWVYGLw58e5kBH3PXVz4EY0v2xjC+pCLHOu3hkD68O/0k+GT+4Qg5b23ok6dY6DUctHS+q
DKnRcVCE/synIWmywOIU4H0k+Sr+gsLamcJJctdsoVIBPcqtfrkUdohJvpz4AB9p7KIsuebPwbUl
0yvuLJzYdDqcxPAywPY6wIym41XdDUiTTB9iQq+1ZL/5Glwc/9+3686gksYGUovTbrVBNFhGyjOF
YDxwH0+KyfeDjgDC01BuuVuIJ8UNs4tM2b9ma0NtIYpH2mEbIvocrYUnJTQDx+Udrzz26VfUSQg1
HIqJXPYkYVrOJnmdksn7yN+no6FW2BwuSMH2Pmo20AzERrOQ0aTxOjah64teE7Z8g+NZizgOFf+I
g2ArCxfKu/Hl4hypZTSwpdv8ZBephuYjPKx4u9rfdxjucojReODmCFMPuFSA2bzRD5KQPSq5eYI3
Atzx6b5v/41mv8yudrW9MKKiv5GLFXxNGqB2Dk5Nl8Qr2P+Q9MYFeximMLbu8jaOzeHm+OlihNUO
JFg5F21Xh2CQk+JTX+bn17waSi00ldWhvwI/leZT1hKvFHNPwULCngDPlWXl8dh6BP14lY/j/L4u
D0RAa68S5XudiUVDSPdnsvDR2FhSB//8+b6Oay8DwwiuiNWyzAAJPty7ikP7O2NP1nzfC4SvJXJl
nnIA5sZj/aPbZEa0UEyqleTL8U93tLEsW1qrTx4Ad6HwjRFFCNs1ggCm7BA89EM2dMyOdZEs9Qsr
tTUbaVW9vKLmlqdx13hDKUmJl4dnbpQ+giMo8gY3Y4Iv7Trsd3LMLP9Oj+x4Yb++9Nv7tayOCe9f
jj7Djc1+Qn6WU/p/FAl+bEyNNFfOhZfUEZQMFUP4CltWkAz/jd1kSaH+EhrLhjHJs1iqW7v2EVWb
mOmWp9vcWAc2mtfTAx8l0aPRIM2516lT7rM/RY02SjJcpG4JGNEQElSoqTU9+1QUWU68qLCa1g3B
fHz1700xBLjfSb8XIOqxNr1hatcKYuGS7U9LZ3vHSq+MBovYmlges9Wc3Elft8TpMVUvihqofZnC
yjX14NomBE2nqgx1YmB2VxY3stBH8o/khptdoF+tbO+BG0Bh2WU2V5Ur84PNvmjhAq8/DwI7b7Yo
b3fmOZQdUjwEO87BfaMXIpzia6nu/MDBCvyYspaJj6fyay195A150EyBI8nJGGMBhskRsJSwhqwZ
lNMXMMph+cpsJh7Yf2IduCWjvF5MKPSE82ojWk5VcFLAMeQP6dZOszc6IRJU9fuavCSsNxgYCpsM
fnnUEq4WNVlrOduO1NChI2hZI4O4MblYuqjiLTf8GjmyRZcY59akl7DAT7oAOEBt/OoNAxY6UQnc
/kEXT3/EW3NL/9BN8A/AwHCyGPcwT+6JdJfDg3ENNx8cRvliBQSptqkPsPWCtDMLxVDvr87+E2vv
yFmx3Oe6Lk6jTE5OnSHAZOFdl6SG0KgaMc8ti4tZ1eBAeZgaFWn94A/yW9TM6dFcf/VLuHUMzDmB
Iev//llmeujOu0OD62vFTg12LUrLlfEAuIvXJaxiE/HGyEzo60rQR/imcFv62BhPsW3LxUUWjbxL
kBEfi7KOwP1DAue9HRPE12CxxnCPSsTaZCfWlsAQHf5sUgBsyfvdd9YXgwOlm67qMY1D0/+q6Whb
PZq081IO0/ldIrzTjssXTduOJfopYG3iVDs0zEa3wj8XWC9r3Khn67QdSB24cD9ks0UV1uebQPXX
b12JwqK4DYLPvToO7JatoX5piMVbz8ngQa5XuMrWeSrsmQwT986Ht80PGzSpDvxRC2JmRJMhcTVv
c6J/l7p2jiVKqthtsstwrn0IUnmCjx7LkGL9quUO0pdzVl3KPmQsEepa3QJnd5a1u4gyiPHQev0q
hj+HZKXrFfy2BE+c8Dix4nGPABp8316HlJ2yyaJ6ijwH8F/DUlL3eOUcgSxAg+Z+nQXNubLrm0Rm
3D/qWChg3FGyPlxmmOtAcYvMD8RXAugD+6qYpFy2n5xAWiaswPdlqIBCn22Za0jCQpEupW2/6o8L
G8LvfdfmA8fdyRXKcB3D0ULpWT4wj+/WLX2yf1Zo3ZCIm7qeWOL4MdsjrUEZkiGfr/ft+uCrf4gn
K+k5/Evk7SjTRZGB4Km2ZBuNepzsgqNfAUD4QEfDun1wWLI7LT63ym4Uu6ErLmpZWMuP04xJxUa7
QMGUvXbF94XTvdbTTAlBTQsDA/yFoFQOBCwxsEyAQVPQ51yY8eQdL1uoIT1AZ8i0wCJ07ew+bV6R
RBVyGMzA1ZZ3J8f8KlXLB9S8SdJy88mxD87hB7fI4/udLAEcT88YpuUJSGsI9um98A0+jRwnegZ5
MD5bGErA7kYJx+rUfgyaVUyueXRjQfqMimUYH4s09N/lJwESLAHynSluUZJjLFvhLTN/zSTQwdBB
ou2StFczoAyC6g3AIElCBdVP5qGoOQMELlIHruPFbOLsHzIND8i7D9RrHPqQXmR4ME2RsbYZyGuz
n069Qj/7LHSL2V1HBm9aEmHR03T8K0lcJMGxZe0vWMb7yTVyz2WznV8frvgWh/I016IpQcoHbtXC
22ECS4sLlzcn3Fv8JSa5Y00tD5bGWkirFJtAhKvYIR9zoMFKFfvsH6U6GNh2H6ZbKsRkIM/oQj4O
OmyZwTc/gyGK5Tet//mniRImPS7nYzlNib45vkwO84/R4RjBYK+fbfmPTiRBt9jzTJdiCK1RaWyG
lz6r5+B3OXNL1SlG6ebRiyFF1z8rnC5vQURt/XQBOclmM5YCB+StrCCH3+yfyhEzQDN7Rod7fvh/
5e6hY761pgGxyAjoqyZKrOSGJMVzRWklzBvfBCri1ufSYULpxjjyWzn/GVGywrx/mIGmmUJq6oDj
hEFf7UAGGQgP9Y4/ldDvzFkBaOS2T/msCg9fVKUuu3+XYG0KtUrobQDiC9NzoS1kY15TUyTY0vOG
MhUm79YnjOZv+CsLlDt5V87eDza/w4xhJblUpV/ulk7fhGzbiJXp8XNaztarHUZevNpnuPVPG3g4
9vM/1l99DqLL7r5jcB3F/9/mRcDQS1fDJhj6OdRFHXQZWGiFMmi7GLJR5ApiyAugV/otd7aJ7H29
vQZQwUKtFaIPuGP/e8jTnpnqLDBAE8jV0T6KqLSu1hyd63tILDTLSdvWIl4b9V+Kh+2M/+8l5WUO
Zt9XLwM5pehObgIEFmjrsF6dy6T3rbzjJ68cZCaqVsOWOGC9kgtHAQZnrOtD0f8QfFiNhFQm2oIS
o1O6gYhnKYUNrHEiePtHy+/F0iPd1gcAONiEKDL6ybOMyC4UMtnw6LgY4NppmTvlVK2owKYDB+uT
YuMaIa+VmVjE9p/6+6CoByBb4dbTz++PRdhCMLBQe+bEu1Y87ys/oXlN4mwJnE+GIxibiAW3X2vW
3pBDpxzdReY/zeHTSgQxgbT4wzQEGQra5ubQGFJgSHhLwITKBuyMzWYbYjISo1aBi4TvDNSb/2/N
viK8BY94xq/KdiYYMm4lmIUkp9G8000RN098Gp1CEw3CYO8lFgrxQR5PXtgHbzGrTXWm9UNvCLE5
cVWI61uHxBaAMh7XpyGXfP/Wnz3shBb0Jb5w8OR9IWtmcwgfNhyjhF65tyPBGX8KLcUHahl7gK6+
9CHOcdOZpplLTBleP+Ice7zoO0cVgCO20L2kBWZqifNlOSLIvP23uPCfMpvbtCG211jvJzTpvsHq
6YrT8hvxwBy30wMf/hB7wg9XdZqaGyC1eqSCNZ61utdZxqHff2HUiB4szZW8vOOZNo4KGvXyDYvc
6FjWTeSc2nJ72um0H9pe3ZoxHsg6CIgnIK6iI9M3eKvD9nExwzo3kB2kbi4IA/jQH73XCHVwKowP
a7ghjgF6CI9VPdsYujcN++SXcE9QJwjfnU770uXOY+M6U3A9FDy6P+od7nqesUG5NNogSlqMtTzp
T7C8+NN49sypFzFTFyEkbT1yxOtP67yE1yI2k5Yv/hn5E7Uzj4y2IUymsOf7LRhmHOaiDF5ZbORP
Tl+7Rp7I3STBewDiZUVaO+FI8SJg0htcB/qgUwulTRNthLxLISeb7K+lyjEd7lXsuzy51HF5kiy3
pfKTwxUiqopxGzx+9kzyeMP94E6Ak987KitN1Y6jaGgcOPqniXOw0Iy5GvKbAd5bh/OFmcCL6OWL
d0yCe6QLt6tsNylEi2cuORehFH30OlgSH/iiol0whbjrTKBjg9as5V0YzjdbuhEG+GCQHjZrn4Md
Wp8lgG/4010gxaGQ/zIbBGlsKbvLXDNt8yCnj/60GtHrbHxkvqvRMpvshExZntCo2cdSO4fTAf5Z
1kvpKuFhfBhbb3Sr437tP2g+4IBdDk/VqTVJmAcqCCDs4Vvg852fGxYvcoYjIbIBilpYFN2ZRhl4
h9Hd7WK3zh4uDZUnHi3CHtsT89RMGWUXNEWfXix+sIfm8A1vuiDASIqcjT5mf9dVLWG4NcR6px8j
Vs51HwaURLNbGl2KMvCKUAhmFwQ2MxNQG5gn+4biZgXsxbtgZdKPJ/bcgZR7qLVe0t57+VP8Bzjq
2mO1nTXNLIz4cTfan/GH7CEiIWuGv2NnNOKdYcAmVjT3Ke5pXhEeQosq575IQWrD4raRt6ZpSIgk
l/t3hNQS7nJlISneXgVDCAz+O/Z8maIDHx78OAJ+qjaI3o4vMtaLTAAkzs6VXyE0+VTLX9Hi+JDF
MjPv+By2vU5RT5kBHbwoonfPC/D1QyAXKhsRPa5Qq0qVIWAHvQeLu+zrSAc5N9dLcWi5ZjM8iBPx
GP46KJ0Or9UfmghEwTfRbl6eomgkhpHaQamkv+s1WS7/nayFHY+Ai8JIeM4mrHJGL2lrmtU0RO0f
L2b2+eLgKkSzJ3AZEmGBSocDymKTHPuT5JAlv7OLW55Pjyvs8TK70C17u3ySyplPGOVpHNniFVYX
ONZZ31pd/bCdMas8q6WdHUTC1oEt2dcNref6njod5V1qDLM1IrxS402G29cJu40RD2p/JXR4T8yQ
a8hllOr3xLiipyXFntLrtcRt2FzgKo4i6eilKnmRKRRLoiFHZuf19uo6AFstIYm9d9/ZnqERRJXP
hxq1kRPk9pj72xSfrZP/o9rxCzNsk/5Du5rB3TImOhe+9dMT3q0I3gVdecqHUIi6/XJCIscFGxnm
+Qd73XzHAQmWbgo7IBiAvMrzL+tIRBrOtsdwaHosI8kDb68/QlmDRFDyIHv8rLFcE834tE6JsHy5
QCyV94cDx2gGNxn6OzkxF4h5trCgZpc9JhRgUQEiG4X8tiMz9StajU592kmrzDaOuSdPOc+dz6Hl
UktTlK7LkiFvaaTKCvWTcotVN68CcoS2mWQJd1aeUuhy6beB/VE3HAomPMdN3mo/xCN8MW5+KZS8
kzkDMgBLaeE70TjSGMcFKduCFY1EqovPlyYfUIqTdZM0Yr4f/lKqFi3rkS4l8UXtEfxu/aw7q776
eOcieqWRaVTrDYQVhhGTy+WMjrrEktf8hzFBR5IBdoSz6TuftKSIVND7h7YMULHBZ2zVNhlEpyWp
5sTSi7kafeyBe+roQCa/jzwczln9RabY10mPw3pvEKhQtmiI+DBekfTctUjBKqk7EF6ymWtCSp5L
51xGYH8YJSNRKdhWAUKMCAxepH3e8xNJW9G/u7FykPMWUThDNbRr6CHsGnGRXINmEx4ZqJSN+jDU
bLsbq1oTGP4EkcAa9NBhxIz0lS3/TJLhnFuzeq1QwYKRit+8NIqA3B6mkNXDbKj19cGJEr8Vxovk
mAnPNk9gMaKL1GooK21mFJnPyRdNLqkIkRX/wfZJV/pWQjI90DVvYtJrMek9UMWw+p1tmGXh+8JL
ZxIM5HSTBNZOy6zvmmY8hKOikb7Wp4Y1TyYUHnrMBR1NhkDSiYfo6ZwDcqapinmG6AUohI1UJSmK
wjU8Un05J5NiY38WnDIxromXy0X0IcHE/SaMJbYadM5drvrhBTst0JDYgkIdulce+QZR3lnQ264H
5X8lFbYWt6jDkyUze0sMM0WBoY/7P+d6sEJtW/AnnytJGsYW6YpriWxoHVcPb/t2OnjB79Ma0A4t
OhPHuwW9gXukHV5u/d7v/czOk8UZiMcAWvvT62lprFDmZ6qNqW14sxdAjXr1xLnqWdiAoFVq/Z/+
Xwelf6/GigGk6EIWwTkT13LYspmrx+PA6PpbBpbRfCWLwHiCDxVXwLgciNsrUWNlG7VdZg6HeiCq
IVVX5lm0rq26lvZzKGHwFa+pF636bUctRmgcZF/Yt/YzJDVNGmjILFIjIZG5gbEU1BmWE8nYEv3S
b8IU2DS9kMHus3fdJBXKH93Mq7ekGIRbgXRCFxhmQOJePAlVLhh1L/vfKRa1Xh9x0MdjqL9qOp4M
bOh0eDBPLKQ+0OCBUoUQAzqVp0b7Se3nv33TvUN0i2gtvCMyhKjPYrVT7YxXVqJuGRRXBhQAA28N
QmTmKWcdizeXpfnDWQ8xIiWWv2UTzlNN356tns2NJMlnoC0pZKApqqWU1wvAVQCM8VOKIIaDPDk+
pw2ZHo465pPE709F58VMss9P1UmZKX+0j40/y/wmWLTyN3cDv1icupVqKMMRMLiFMg0yvoOg9X9t
DfbYwB14IgPmWlQAGslnv3RUYJ8dd2nahFmCBiE745xKd2fVaUiedG3q+JvLqdE0bbhlrgBpnNb+
lR47ENiNcSlXBwM9scfIWTq8bvsPN/grbC/AkfXz5o7KdiECWBpe1kvhVAGg1zSt6DFMKFfyxTA5
tyncV7ncNyh9T+j9Ulkf9hzbjVoIn//mpu5aDPg1GWa7ZACe8a/1nAugK2pEy1pTYKLmwf45ioOV
c2lELaIH9xN6OWELljR3AJKDdgsajo1e44NpCZC3OnNcHAXhG0U7njxK+SSKrLeYN1WUet+SxaGc
ysbmRZ6RfO4AuTm8UvUP/uTebBI1ZQlXC6A9pK7moZGYNN2auddtqdefBRiqw0TsbdO+qjQwYXK2
jzlJbCyy4JAZuI9BP38D6z82c8dc8HERILLub9qIOJKcZ+NVxZhK+fmbPIiBgYEk22SBOOWi1usi
YUcnen7lvEehmEwljN4qHWwdY5avZ7/toWPj/xBGcevAMCmGgnf4pmAgLPhxoWx5ptJwCtfRalRp
nzahX4ZOR9FAPLKMh5KYoJb7bm6lLLIMlELvc3Jf3Z2bF1lE59cuq8E16kyutQAa05PjR0xqKZ6C
PxfR3wc/4aUUYSzzLhgYDUEVSZF31AGcsgEwNC12TaMpAmKlVQw3NQKQQz9I3NC5LI4mVKpS/1hy
BZIUg0oi7JThq3IUA8OOeBEhU5LfP2nFO4poLYkKUcpcqOtxOdmFDNCeIdiQiylpSJrr90SutHD+
ASlZWtTrphlvs20L+ZRrIlMy6LbxMOoOaW61ERo72AdE0Rh6brq7C2XpJRiDiuKRZ/k+zMfHJlH+
2bQ4GSxQOgSUl+zCR4pqCgvtDFaC783mygS6YeV1R2rXBd8HB20V2/Sii/qCl8aaZpJmAgYJjoIR
dP289YvwzyULR1bCXXIxmJDK15MiaSnAm5S6JevyVl48yQGZzN9r2y5pGaDmyv5SxVhi4LcwVTi8
RPqFNhYGe5YIpCLrwVDIbeneQcgoe7xjdErtintO+/s+jFq25rdZD9lXmJ5GoC7ko66IahpNeiP6
ZBux7dYyKqAXnwA9RnPx9CrOkM62dysrUPZZGbMscT9NokjYrI4vZ/m6IbgIoRBJtih+DTrquPrW
3n7UZ5Cb85xnOpDt4WNq+1+1l12CgC8dIy+GNXeDQwh8qPgW+Y/a9XZG/qUD/O0VbAxlntL/UbwZ
fdhExSNozez5UtHy6b97ZFvxXElYY2mIjPRaOPn4eaJo5CYrrvGUWyM15IwTcIr65w7wKiVyc8gT
jLJNmvMmNpDbLmbg6Ps8HbGTQ6dXHgVEAk2DIBlXGEgeQaq72A2E4R4jvG4Oc3Nu140DhJzjDgjz
Us2amT3Vz2+d2dNIplYYMI9FVFbfO3tuQRkYH8EBEf/HuRq+pUJE9J8/1jImLzSVJpNY5vhnnT97
WKDoWcHSbZJL11+GQPs23MV3QJhO2NWjelWEQqqNc8djs3TBXuGuTwhwdfLH5rR1dEquyrDW9yDB
ftq05y0f8Tj08+T2AXFVnSJaTs4nQlJ3mb3DF9Y2VefbTBn+ShUlxY+GEeBWPRZ8Y8icU7xxf/7u
WLCyvZkzZGNBkxjUmGsOAziNJIzj9s3rrYZRxYKB7sRWZdzqykSdmeZ73cHzKjJAF2xXqRxZkSvJ
p3RPSaamrGT9LWOzgZn4HP4lg2mTtqQ0KSKn7FSQYyiLT7y3/jGwDkoeeD2qiN+qH98FPrHhZEvu
jwJx8AkymPN3kvWJXpqeRucfvqFV3fytLWQIOINQvz7s3SYo42D9pAR1t6tsslijYhvHflOFr9N1
9Yz49LSlhg8/MaE7Y/FgcCUmzW2o8GFuaic8QSdbsjEK9l93/oisQkdKfJWT0NzOzNMuk7e5A6oW
esLXwWVpy/QxP10YPG8iVc7DcX0v5CGxLsLOA0D/TOTiwDwEhuTlppSgsz77WHm2x/toY7eJVGAA
DFiE57uyvOeRxs9We7Pg/5ILXIJzdn9NNgQBZdxqgqbyGDbYgXK8JTBvuDcySY+fkNFAjmPqun6m
eNaVg/v260+qJVTSKM+i7CuQrsn1BwJKzF4Y2/TvZ4478Tkl/6llcFUYA2fqfN0XQttiL2Mdf6A9
IBeea4xSQwF6PZyGMfSPm4kvgStcFIQLsxNwfd5s56OY7R9Y3NmEkNb8wwaQJQReyU/maew3/ac9
LqTajL92QbBVqH9q1Ju46wURYEg5syI+NyWp3aNmMKhHpH3fr/e1iURJrEeOtjCyH0dD/oDisbpF
gt5Gh3Z1dS4VX6M5hqumv7nXYldR9wmk2RhHn3rvioGQ5JarC74fDIjzmlO2pdZs1LieHTRNUGsj
lAq5Xzvj2RuK9H5ChtcyWGuZBMNi8rR2uclqf+GNTbdvf2QCpgNRnkrvOzXaU89BNkDN2QZ3MTGL
0Myge5yi+tAb5KvG5F6O26kDw2FFxORFsuT0K1dOMs9KSKk4g3uFU+0iDWYz7BxPYaINiDqxZ5oA
Oc+sNv1IKw7j4sAoos7au6UUn1hAd0CFubGxlqaTUH+r5GVa2sLGYI9AE9lRoLN3dYCm62O26Zfl
6FfSW3ngp2D0n9lCGy3Kdrgfx3PQNacd4qMU29w7x3/8hjAMAoKgZrPVkFLva/sxMih85puBChdM
mA8qbvQlMR8nQeq+qGeRAuuHmdmJwP8xZg4MyPEn+TlbfN5zrBysYrNem2cHUWFRSixtGmRx+ML4
oDd0EDfThure2JDHOijaAU2pj/QRhecKld5xpH+SAfeJ3yewmBRnVTvGvrSk2v+EL7a0+O4uyz26
0lyo6WSJIC4PS/RoLznjpIDsbnHREE1hGGTZebP30dPmTm/4EpoJ/hpJlQ2xLCvMQ4lbmdD7awut
Qi1lkoH7uHyW8N6eyW3H0f9e3hj14M8Dw4zXMBUoIiT44nGrTjlcl0VG6o/j6yksLwjeUcjKu3Pb
2jMfSbZXrRdpmCe/dmYEeukpqlz6844NLrSwixSMfHuUV3YTz4m1KIFk2OeP3/t5RzmQ0yh2Tjud
kq7rzr4HN07DG9YMS9vQkNm3+RcKHT9FeZja5Ym+k6xb9aDFHtMBTgyRA9yxLAb576xFsclJjZSK
MnAlKDKuu3k7GkvSQSe/ARRMlMN7N8kzAGTlyMC2bXlBshi1umrxloSJaxn2TW3Haw0nlWTl4QGc
2lm4I017R4fi3mqe6XAKnUg3g9zEC9UqoBMnxYAISSZpuGNr2Z7wDeTNviJQ0hoRUnwUVBKegMO+
8zCriWH35Uy8BWlARxNBTqc6PxBJH2C7BLEaMqS22uiHbxXhsUahf8igFdb273uGQgmWUM3gB8+w
9Z69hEuIvxpmaTziIFdQ9/YZf6TYObs38NASCNKgWOi6vJUs+irdHGOhmL0L50tA1tGiSuXK5V2q
teV03SJxvwGhQDt8YLCVEHae17aRH5glwuJPY+4PtCPmx7KOnvFLQ7jyiGzBDNG3mERbjAWKRLwZ
7sOQM13WYQOSdSFQt53FBkUxsyXffQC8WVbxHOGNonaNnCLw5VWCJZY4EKdCeSUVqE7WoQf1MRkK
lMK6KNSfSZq3/DXJiyuGx2/UEHosCd89bfcFh8KslJX+578rT0JXsbRmCo0OT7BNre2M6+TfyTlG
rj0FGQxCiOXXXYyZWGwfvjXfr57tP9WPqGdWHQ0w/KUCfA2XolDj1j0cS1YxIwScT34bMpJ46SF1
VfZhBIXyAFkG3PpsN1XpbmWbs+eX8sz12XMFhKQe9p6kQLfpAaZPakpy43EG2lEPi5QxwP/NRdyN
aIhQLxj/pvnvc9qLZlz693ce8CGfAcXt15mvhSZpO/gcOXmuR0rmChVtJ8fq3ikTj9ETLMqFPOry
o+AiZ9D8EM8MtofHU5CQz/tFxoOznxlINJLyGS+mbfibnZVbSib+Dt16//GYsYuXIp317BXsZV+S
mwAuHHlrvGO7ywX6H839na3H5eturQ02+CB44ej2qhd5lscTJCScxYg798QyAJxq250LrDmCUiDI
ry+0cvKwR9mXserQ2omhtDBsQfAB0wehlTvWdATe+8Mu+Wmdzib7EWH+MYJBtol6bv/Bxpsxpzz6
7Afs1Y0ez+OXvhjFUg++2E1LA9kSnbvnKmGPtzWaQ2BBQWhbx3yH0gFoW3AP8YwwOljIacrZGRY5
nf/utp3AvchM7lH3lWxKh5UbNHGA72o5wwPi6qq2SvXrfmp1ciFuHSeYlVgGtZOANZvx7qZBvUVc
RcnJkS5WSnJASA3NcU36p1kwNe7lImVOlR+Ls+KuqDh9lRzPDrz3HHa6Ngl2lI2tUjjAi/Wdrxh/
qDL/2T/Ya7ubrgXspKFptFJuylmRJu2Gl8IkNyceFx2gV5kMSsm+QTF9XLIDTjovMT1vbR257Udk
Yn+1fU1RxUYZO0tqVlxcPbnJIfGOJPkqUiR5Lm2Dsed8VLKLiD+j5RxSKw95+oTV22gXVrCS7TfR
R/ovyhv3kRGReQBKV6/QcuJglS/LCA115wNmnbFQ9Rx2f8B5oL49SvajOeaq6nmc+wHS8KNLaZbw
0m7zm1Jbc+inBQo57frkFHSDs5KBVC42LnsO+FjpS0hJgJBblgiD4AII+F9l/wvEm5UltVh8Sh/I
BeAzdts8axuTMPaofx0DscVYDUl2Soj1hBnnj7HQto3W2Tda8D2wa9zuizZsOxIak6q4y4Q02SQm
Zp1x3fScHb9i0S2r2pwC2S9k11HYMsjyR5TDLevxJh36qyLlGQBti2T8NcDeJO7cq9nEyJR3kp+w
cXfMW3xjSpYiqRK/gfuhHwyhZQjwvFrVN4uu2db8sK4/a3u2o1ZOKKTTzKkNeo5O6DT5Hplo2fpM
Y1J9al0BKHZSszbe6weTGgADtbrkPU6iJzJ/aNe5n7GzZudu4hSIiO+OfIx8BTNqf2VexYam7y2v
Qf5x//A6LvK8zJf4DnfkLo2CDGIG02AWYja2GvOyflgHNP76/SvqPXcEMjJn1t3k9kVV7ybmGHzJ
vkaxuKxUOjoCuS/UJjduuxVJVN/oarsWQhPc7Yfl2BO2mwUU+tFTth9wD5bBPARf5FQa10n4zQkj
qUQqss2IGs/sjrK3wOZj2iF5n5hriaAfpsIbwFt1/6t4oHKf8bzPJrbhkzxRhEYOUZT84BGQTV0x
B1Pr9YMU4fB6nQx1RbS7KKJJUEFTP3HyTSE5br2XEiFdgEnSUcDpVKVXq1SlswzkMWPuYQQ4MExr
X/j0hEozMWimd1sVtHGZPgK3SLlZohu6FGMBs3ewtVYCIzwzjp/CI2NjYm8llmOyafYx56fTl5dd
qc+kAwZH7LtIXBLAbSR53d9aeF3bgIO3m/DTUnDBF5oOhroy/6/aZIYkF/pLO0xdkceCjPm5CdUT
iyse6v/hcuWlSjnDJz4O8gpI2lEmDAxenyX87LQGfnA+wvNxW5AL2KCwywfnDEv737etTdeklpzt
upO7FnG+4hcqw39wrSu8WDzm4vOWkX/dChwtdEPRGXHsnthqCYE21uQx7M2WooDnypA3qTmj9NPh
6f3LFjF/x3SuQoz3JD0N5qQuxKKqeRBNrT3drVSS5GDlOD+okHe3BHVxQbj2n0k7WSbUfiRq/DWU
P3T3Vj3+zowC8SHQm7PuSlHlJwYrrX6WDLGJBqr2dTJbP/69xoqjrNPRfm0nKqaSQBZj6C1Fs65m
belq93nrs3d3RsmrS1sh/+ngZcnWf2Rrfd2IMJHFHrELfx/xPSVNwPHpXbrNfwovG48RNm4kZaqt
gg28hihBpiw+BPp5tAgou6wD8Hp2eDVlD6tow5Vp6QPwXEwR/gZaBwAt9W0oLbXTM61cEctKqD6H
hqULUW3vlQsfLrKh8+377ME4sNflIqGu4dVkkcGoDsFjNdfJfyhFrGhA2Xl8SYwS10/CphSHkQVe
ZGGBvkk1qsek5rFc4r5cddpOQ6L7c9VwJ7fuC4svX0+GHMmZvozxLkQnPvCz8kgEakdhK58tAfKR
DitVxnTvzwselL0//QiRmGT8xpR48x2B9xUA/S+lmCqv+2RjjMrRaSfiMtCk71gtKCoeacemmKPm
AZ+MnEvjDfQjvpBcorb6yECYympDHWYprwy8wMQFFrKmrdxeuQoOGqDGB/prbcOUhnyKDFeOpKyy
0a/mbYW3RtkA3SUiaCYQXHIjV7TNm5Xd4+8qsX4g//7vsINLGUl09pvbDOzer22P8je452U7ICr6
cIOvbrtoWpfWRMdyLLUYM1o03Jphya/YhftIcDzVVza0kTaoznjml0fisxdj6iWAXXIpif/wn2LP
ALZ5ty6yEfxNEjiAM0AlQEjIGaE+VKM544bi+4QymfHVg7LmuwHI+LgX6cBEYfdGoIatvG0z4gWg
PZORVLQR4nczcmJGPT9dHwjrS/rw7MqkKm/BLBoppFzyUvW/ALVkkTsGK9/ywjyMEcILknQadwnF
CU/LKh2VNOSjQ1J7wUea940cCRwDmf8jAiXNqrh8p7UNytpAFDgPp0zqs9w5jB6RfsKH8Ew57tij
FNAY8AH7IlMIvYJFF3vCBi1sGcKNZBQtj6eU8IhU63y4LGXVeo4AkBlHKIl1PA1PCb6ErBPhH7Oz
GWk3PALP6B/K5p90xbkPoHwasIWSR+Ps+R7vaj+A7e+qC9CblaBm1ifFqvNmiGABP8Blavz6b7yU
/WXUeOpXHYx/Ge+sOD/uiwMavhYubSdBDIqsOvrFXKypR3uhea2eQOxofpb2vE5zuspqRHOTfp8u
OsOKFPosOt9h4jLBge3fC3Y6xd2quwqNbRGQ1JnXbfr7Z5rK05oP4oaa41/poH6+0Y4W3FZ5XYe2
sSJgz2Aot3xkS+Di/S6T9p+8F2LI81lS4R24kPO0p4D1DMqMvJLbwvp2rLOwOEVLpOTEpoClQb6R
IPT2BB5A5CqWBlkgsQ1nqrDV9KSQFay/18VC3v3clWfSkOpda10M2fjfNjEeRXOZihFRvDar+R6J
NQTxH3Oej49CywRZvnb7pTK1MxlIZaDkengMT0sFQ47qKlGsFPBezVXDZZJgNXTUsg01lbTiCQzV
Vu74GjwJ9t+oSwgu+FwAxXg5OU50KlMr1pbHMHjAR3kvaN+c9r8rWXTueSLu2jQ74vgkq/i06Je9
rnM4+AsGBEtkQRXY3u4lSqHwClTY4k7rboly+JUkJLwdfePEHFrR+CDj1bRclco+ybcfyt9FsUac
9vd/DzqMvtg3Kkote3d/M8yp64uD2N+1S+/WDPyBGd9FXYy8aOu2nckiSH7/4ArTCeEMNcsoJMpu
605Lk8z89pc6io7WNJG0YolU3anPFNY/XrGwvDWLwu52HhkmG0ELU3bulyMlP074Z50m1X5Vnl38
aO4a1RfMdNLBXzWqrq4oZLZuFQJuL/Qr1S1Spu+voKxg5tX9AnZvqtKI4hhL2Fh5Yb7pwInN0E+h
93ItNgu0853WB1vKhiqQpOgG+cb9QduMStXlTcxx9PkW+PRCkl4jCO8/j0G82CtOe/vivxcEaaY5
sOQHaFRe8QUt8OejSDuhzOuE6zllR+X4uypmaeJoBhH2gsntDScO3IOm44/J7SJFH2c+02N5B2YF
xloNh8W7JNELHpkiViYigkJJFmciFE9g7NFCY9mutGw5nvQBjmzr2CcJ3TO9dsIW8BhR452HImCo
/TOOi9VsAuNTAyzUDGDnr4a1BtegQ25xJRwVSWpQ3lrH8kmlweUH1z45VxA1Mo9mbmvMAevknUvM
xvwF8/JLEeTdNPeg62nBJa25wSVYxmRQD7i0ANxr28CAn5e2t3+ebxkcZO/nhZh02K1xRarPOIVW
+Q2wHIxXklOFXDPNgjWo6RImHIjJ+eV9vkdb5T8S6PHRac4z+1UDr6mhCE9BJKj7VzvaXmN6neIg
BKTvQMx8LFEkeVaESLS8voZOBEnwFe3A8xhGukByA9eaGGP45dneGGGruZFKV2BQysaRc1jeWERz
pg2IOrceZmiKb5l5UREdnAr0Ws2/AB5s3Z5SfAqnwiBdpeu6U+PJIGHl4ejcv7KTjwRfDcwfWMB6
B0OGwu0aCDPcHplQUHaeOVan92TC5shPuuc0DPAjkhig14n7OniNSurHCZcjkP+H+eHJNeFYIohM
se843XtwD1fSyp+vYGaK7v5gIdVsihfZ2p7zmOIG2ywtkd2TgkY3Z1U35mLPvIxqnpNIzI3UqLwc
cC/ZcLf1KCAU491UtPBJG/XE+c6ngB5tsDhnGCZdxJV+Hoc8VHeCnv2A1PHx0+2zK6+JYQvacw1S
Dqm/wIs66rjLJxeLFPo8IDHWB4JjjvVCB7VkKhc8Mf9QK72nqr/3bkbswknIFa0keFM/RTEBbvn0
ixmMq33yRTAdQnmUXjoJxdlnTQFOnCPHVZmqJASAtkVruHkEJK9WxqnJ6x7LX8C4j35RDanoX6Sa
6TU2c93QiaYaSLZHK3daVwrU8GOAejxdsWsF9jJD+Yt8koYtsRFwelipv7elKdT5CuGAs6Xd2v0i
gRnDEPINsI2PPuIodSkUQI+Ojc0OyjAhmFOh6gPNW9cxKbWQ3+NleuQOUkrRZkcHDug6x1e33TO+
5QBloPHFW5xp3tmYfMDpeDdmHsQgTDHZjLAqiT/FgC2/+Pi+NDvn4+Aou+YGSsmzmEQDjJZGuzgg
lJXQPzRtI1HCw8mfYgLo/uPFJeOlng7iCUjf1AF7372ROxxJS2POCNT8PpBJSi2aF1zM6gFOU3Gj
DxEoHe0Bg1HehgmXwnCkR649WQytSru5C5D2LoQuumG6b7TbOKjbCXpEA9otWTeMSDYbX9yCPfAX
DN3e8vC29H4vcBdPPcEaGVJYPbYdQ82jTOdyPYemSZ5Y/oXCn2V/A4Yd+yegSArn6/NpfQbRDCFp
JxgqRdOxA8okcYSmppFtyydmht3aDUSml9CNUkbsRGf14ihCHlqX5ezxIqYH9RCduujmMGmb93Bv
H4myRgL71QYLZTwDqY4cL0GNfSu3pR1eVh5SHvvv2nZmSFU8hslxhxg7r3w86iigxcNxZF5Qt6Mg
BDgo5l3xK/ggnnR8h9Ge+WborK6EyVaz2myK4BIT81pFSkQfkc61VuOVRBXN8GBLwmFoltMpfKDK
8b5FgblVv2kXsmnsTScMozy/H9yRQQn4oRynrqr3cVX1CpVk5y+LO8cMFAA7vPD9/5T5AZ79j34q
hBI6Nohu7gQdd0fhX6DbmgyFaqsfI5sY4XB0m2zJ5Ep5XGKmHXnOlmn6Q+xjsGXxFOWRWkn+bbmP
6dG/d/8mt8lsbhIV01LEobA+0HJBaRvOp6Hgf+p5DdzJ/a2KFJ+O+3f/Q+xEBhvQajw8PjYzAU+v
cM+oWu37div/SuleBWTMPYjVxscsrcUhocNiDY9qkLqzRg4HBOP6LYXh/+Fz5L7CLE4EpXL4E+Z0
v6V6LNkwkzpSliAe/NUIAviKonvFKwMiSGgU4bc+1ZsNt1Ac5kalLaQ8Q3YGVyaOUBjuxHB3YPHF
AP8yAjkWpiDsqPCncrnaAnypUq83WA8/Tfi5GIyOVFIsrmQkZT0KG7uurAAg+ws/o+7lD9LkC45A
dKkPP16zpdO8tg00JQn8TWfAmu5JOs2I4I4zYMO8p4x2skzhffYxjMM8aRr4OidnSbkK/4/57ygo
pGDyK8X1t5XJ5hhHmHn3+9f49ogRkJLE6pG3Nhv2p74zaBx6gtyyINZw1sTBWST4HGxcOq3Z559z
T7m1m75fx+fLRlKh4GiErXxYazKgv/o4X1BIGO3eo0qfDHx5YpJUKyty+IVhZgiRtti3fZAIC6et
t0HuGMzUMZM7PYqZGzJrQTOM/Bq8niHx9Vxk6mhGBh4C8MhoVgtmZmDslLC80YPYaIGKQO17pMd+
7cDVvB+RNQYC98xhxoCVkhiwLQbRxTem44ZSjDQy3uQ5YL7cxYCtqo3olR6qIQE/G9P7BQi2fLJy
ollCEIiDfINee4Wdn1QWNDHNLofo1Ut40XdWRMEA6bqml8jQeQlOgWi+hzGXITDYYGHSus/EZFKD
PmJCJGsvFWgRbXusk8r3QkyofxuVRR13WhuJJF398yIH5ino0G3MsAsFRXQ2RQ5tTyXT6MRPy3IJ
ruI2x7vK3B5O0kopjwX340Jd5OVJxxZAqvhVTvHLxIh36huxomxgAYRwxsCA5gb1rTCXY6Jpub5V
NI7BRpKL5PHKMW+8Kc7Lh6D/nI3DRtznDSiEggfX3QCEdOaS8JvE8LdFdhto5I3+KzaG0yzghmRE
anQj0Hw8RqNNgR08LDxr0S4Lj3J/vVY5wrPB2N/8OQs/bbk4KMgy9wW8g4EzuBOJUPHT9wUFacUv
Yt527z1hi+L+1RffvdST3t81H/TZ+xWSTLz8ccXs2w9UBjvLHT3P4SenAc3eOe9EUXHHAaECO+3v
43RXAm8X5pzXLvPsMxbIMv+TUjfLd4b+vdGzaiLcVgR0+2VcFCCszg91qpT5aA7HYSROSyCBWc5b
mgFATFGsMQKOkWVrSXTqnozmAYRzQP9ZvvjJo+M6n41sXetLd+Vn7yBFPamdZOgeIs4gxUKEySzw
J1A4CV4kPfaDYmFZGfTtC24p+zq3a4u/98QPpTmInwiUb/ySbFwPGp0uXJInPeu6u1FBclXjsHA9
cfwVwcukHoLN0KYiarI/QQtPIYoExCZ+qQZoeeCK3WIkpZfi3jTLbZ9KuPcrE6860Jd6bELLv0qf
1MNTnOjm9M8DfRY3QW/evr+YlLnayNPSg6cBEgJwy7ytfb8UDOSeoeiPyYcMLl4s7vSA07M3NJ5C
zvM2hke6qfukAB6cIF9mLKNwXfQNS1XfkVuosI29Oq8+rRPqfrjRQ8EgzUlVn6EDjOqHXGy6Hf6F
jEcuvWcc4zG0AA2QJr7DXECAVpNHV3jrHLTyJ+ZycMeRM6LgeN2ZmfJV3Dynk9ho1D1dyAFxe/xH
m8xdzi1e5TO9/2I1/Dw0zfTkpzWK5J9LKiBoZAN6b2Vmv3PNNUDwOLaLi/k1KussR6LlrQI2YzY5
sP5VdstTmF9rYOwDBirLy0MoUsXJn7wc+SoYG3szej6MwABSBueWvUhLF4RZMg1YWjCc6tK4cJom
NqhQlnrVBxSPxnSD5Fhl05n7s7ERnWa6uzUP01VD2UlG+C3bk21hTtEJ1eV+X6Zi32TGKRWlPoBB
APkEswLz5YXn8GafZ8NWezICAVlynyPdAbUQV1Mk2Pxz76nx3hHPiThRRz8vtWDmIuFw2h91x51J
YKWs7E3Rv7H/h31qzNhruQlOn4YGNMJqlxn2XWMdFb+2NsSlGNJl6P9Fur44zeYEXmuHI0q+pekh
EkBRBTcaIj8MY+TjR6+ZxuwqQoqfOTXFlG0lV77rNp83fEpqUDmYuCgl0oOvuYGNeI03YkGVh+zx
CTH28ee8c13ZLjfCmQUUXfV9YhnaouVC6/oXlPCFKF4fQMJaXLhodkWscptuA2l/IKQHPdXQ3lKj
zjGEGs1BaHspW+D+w6gj+VshrCgUF1yqN4kco5+FgzQnDdgPjxqPWstVJJ60rTgX8+q1Q2gvFsR5
Ei7jinRljq+oSZH2laD3YjtpgbJSFIHs7892TKCgtj0XCkl9IGhMO4JvVHe0XgxxcRUpUzE1CXPC
iNRyMhl3zG7rWzhlFXjaGok8ECXzSbZFIxmZocmaCVdH+S8GESCyjsf1ogyq/DvtNHgeJiYgjbPY
9xN73qNJqw7Q5+j2Wqid7TTS5ioO7Qlpf9hnTkdaqdhNgLpg/0HZ1bBrtt43Muum8ZJG/6jO0nfH
Mbz3Ldr+g8KegqmyT9MlyME47PCrzfkcJlzkPzsiPWNtun0dJM037t2sisBcj1l54fXvO2YksPSc
nYskKDeq6k58co6NvMdqEBb09N/ijMOes//ZvxUGfpm5uxgpBkRS4La2a5KW/2clm4YrAs9NtnKo
BsiD4PsC7/GAk4wAvew7J4s02Vo/hySqnLkR659bRPYqZspLN5geM+50xuzsYgmNlQISxf2WoFgT
PT3+1124dEFqo7tzhQWVyt5U2akGjP1YXd1CVX1SlkcfJLUOemUc0wylQghdZI+uoraS50a+2uP0
SeuIZAugkcpanaEqbUSXbrfsd7idk2Rhu52yF0p5rplK8QkWboTp2jwUHlmyVL+H+/b/1YSG6NjJ
M+6/VNJRTv34iRH7o69HhgHeS5J7SWxfVb+vHiMvBvGKPXQwTzQ+z2uHPbFcZib6jkaPENJBHlz8
UgTB0vqjVNdEZCSDucH+oMSIDj0bs61+n4iDkPPP/JoZY4+bJqEblOiSyXaKd7yRtxRHV/FG1vqC
pY8ok9mYPCcex70zRrVk/OuDFmE7aBqamLggE9KD8kfxLY6JVvNTwsjyozXBo61ZSVoVg/kQbWOB
TBeFG/pxa2eKXXFygb/jDlG3QFuAm4t5l9IMB/xbrzPFpC1OiJDRlpg0Yw5HCYM+CvHQewTc5mYb
u9wQu6O2jbmk+0i4E4cAyxe3i4ArCkvZaJKyOm8vj9G0pzSCYn67GFOxBDzOQYpROdao6q+VgAGC
HQYMzVuRMXK8ob2QH0oP5mWMFdE/iq4sWxE5Koi6Q4XSfStlrmuPVXHZCoKYicPy2OHFN2A8zPIe
c6xdEGrNcMXNjLK0/IX6LXV0+u23a9qqAuXfnlEiQaSzHRL8Zy/quWGxMkBFRVujDPcEUdm3e6qP
OIdmQRBn/6sq7OeUzdQhArKYXQ+vMmIrKV0YRnOvwpZZAwT0pE/Vfkz1uwAm0egtObJNz7kV0saJ
sxdzYwV8iDfVq9NqGHUEeogfZXDpptbs+xBVxMTxYA5b/f1hHgKUkUrdq2ZOYlqMZpDmAlN6rtka
Nmco6+99h7oVCwjwJAAerQK83jep0e7hDIoxDRY9ErTA2s1n7EkIUzx7IaalWvPFtSAEVulRQXsT
OCaXdH45Goy3vbXngGM+MPgpAQbnQb8I0jura6zhT1EG6u02nfdwAZ7FVyI0FkiaAsbFk+uxCTUF
kSR05u9hNtidMtUsMixkyG0dgt/ki2iUHLLndxyqSmPHe3pwAJXmoO+okPDxiTR2aeo7TVJvrbVE
HfW7WYuO6UJsnMw6IEPG2G/Y3EGuM8S5BJnWfHy7HXCaRyvVrPN91SOwqeOclQGZx25ISp+CZ7AB
h1cYfUDuNcjSnLhqNPHtDk5UWnfM7VOTdmLBhV+e/twoNJ0AIiaW3pXk8pzp9CQX9dLSxeWrER8E
FFFPIk8QFGSZFu+ZcXijgB1s2om9vbBy7dUg5NsMlgS6xsJo+s5n0Dh56R7k/nhydgLxKSxkme7t
zL4nTJxr4AJF8BH5ihZpY355PusQVCRqkRkckzkc1EdAIjn8H7HJQ0scXGfo3AO6Fj1fP4wjh6DE
k9HMvN1XhJx41UZOapgKwbVp/d0fkVff0QgtwrBuZFr/NvekjWAEy97f8seW4g4tbvXuSIJlZw4y
tRFyXYjZJTlSzVYe74twpIoxSDUmtWNR748Oavn0xr23/QTp8+jn65003yRU6PzcN543G7ilqtRs
+bsw/TnEt/x8Y42xIZvfHuh2X98QpS8vZweNpbuRnlPVfXgece8EZqNbcAwN2bfsorBdzm5V5q9r
M5QE3Rx5TudiHWu+mRp4bY4t1nlSQuIZ7FBhdQlsa8acPKDoHj0Oqmc9swuIM8PJWDtIzYKH2jzT
wbz5qnO9t087TZDqFjeeRjruKpjhvEcucGpKPYm5fPPGc5ujX7jWSbOXUGiBVE9v6jMETuotWaka
2sI0gZ2coMStWmoXOr9QimAeYl7PhHUOt+m7SzkanYZ2bWUvNLIRFRxml0H8ZXP8+mNy781v7M1I
frBtX4hLIhL/SwDKjWoRHl4bm6+yOTDg/ZfDQ5R2eYH7QFo3VZQpUfh2vleLJcPeDmur6sTKDEyP
phaRXuypeb2vV2rUi0jpXDKDgcRAwSRMd6hAbHy0Wl505WQt4rc7U0J3M9K6AI78/hCqL2p16nEB
EcaYqSGUXxLIicTSd/K7qSI08I9BKJK61ej2GW1qi8seeozkCU8aSVzDiVQD05oialuuA4ZKGYDT
crJK0btKOet0Pquw1mP8/6JxKWYvt238Uper6qj4TOjGNaCSK55LDUsl0dgxoX/ADBbJ0MrZXy1c
7DOPE1RO4UL4fyKHwrAhRmizBUMLjPnqgeO1T6b71PvELsD+6tnrAxCTSNPPcvDAv18im8NSOI9V
tNlagdneupYQBCDr4sLo2ccvNRdCt71R6bQYUbgdAGcn5qAF0boEOSqaDmhOS8BKNtQJzehp+8Zw
c13ymlfjKwBt4uN6fqvWQKtr+T/A5VyF1iNs92dM1GV3qe5CzTAim3xouf+k62GA7ur3ZNkxMsCK
KrpS4JQUjL+LK2OLp8mDbtYfal4d/54k8J95mj1ku8ytRkgmf5LlQgyT68idC5QecS+dz7ior9dF
GbfkgkxZq+YrwGRPFBoBq2CmmzYxGZ7d12LMVK/o1GMeA9IyHR5EP0Li9wMt+bDm28pRivY/53uR
liOS4mjWWANkzBhMl8EhtjIl8BH84PwtwkwO0v7pPcuKiwWdulDJSxJj4u3Z93g7YchKC+EMhVLX
zqJDbN+o5f8XQlSbGDu6NtX3JzkkOZq5WJ3NEoWIRcIJlr7U7T34QfZeanqhqq0Bc+WAzlNPpd2z
nLg/m6bXIsIj6duWvFLRzRtlCiYaNnn3o/vgNBtsPJ1bZBklNS1VuorOgftZoTmRwSDJkKZipQ+J
ffHdhXKkTj3Rf4nY7DDjt5n6uMOf1w/lAaJZ388do3JDnJ/fJ32KAuDVxahLOzusFJxYJZfIGv+7
f05FEY7LXLoa1rBXRB7CZp2JjgQVCqG0rag5hgmARIShJ/RB0KTN/jlAopTxmc8tjuXEnkqasC5h
Jmlh34O0u660IGEahKRlmzDMqyFLuG8dAIPpIU/mnCCyj2WtZdM3uHZ/hWoV5mEPKCe9Zdi6hxFl
FA/IMiOKGspZnbifJrgyn1LVj5b+xRf20hvjQcmG/CQEzpzulEAenEIoneAEuVZDW1jZt6iCiTP0
lZZLJb7Ct/hc/JEkda4mcXrCCWGbjyBLtjyy593rcRid+1N0eSipSbemaISnP5EDyRxtgtw4j97g
psmFBjJ5c0ELy1Zl+BAHgfuNncluP6QaiTunY0wq6Egc+9tB234CdsxcJwNcUU97U/ufYccvFjvG
GwRuZ1NUDSpCgSt3MR2juijILKz7scOlz5MkO476VKFES5ytnoUTsMd+nOITMvwxmE2tRrm0t2PT
HSMM1nAjQuhfeF9ZtnP+cWjyCAWCbfS6dFGuvS/quOLhaJ8wF0Z9Nuhp/uXhZogXFWijeR6rybPs
2m4DzFhKD22xw5RuUg/v6LemiNEWdywVGFU1TjGgOq/+vW+oAuah91aB3ppH8rB3GsCtQyD7k8jf
BW+SxwLOt5VidsC4ogKLkVfKqaJ+fo724UdVjwYiVEzhgdUIpFT+GkOHvyV4dDz+AHiQFmaOZ60v
V2XabpbZT4uexziVpG9BaGeSypObBk12I6dqrcSdxVmIaFRSDLAJ36EuOGeusm0oUs47N1L43Uw+
z1MFyeUGDs6WrXXf0C0omhCieQ31brgMy8Yq44VAlct7mHleGZN3VOhjNG4DQppkLmPeobtK+TD1
GZn/e3sLodmi9Gp472iuhKp4crePO6liUlqj7H54tcGRIT1u40KUrcV6+SHqrFqb997nxL2rxymW
sFSv1CUgE2TvXEdvj+ABoVcsQ3fXjudDMx/gHMhoYQIPOF5hx2cl8NQGOVqB8txN4mDPKSUGiKuh
sehq+kX9f6W61Jh58EXTznpNSAkZvze78xeW2CZbvU4WwXXRGCI12lXqX0r3EpCY4+9LLtKdibQD
n/2NuHQ+F9k4byk57aexlKltQkzuYzhnfmCH27jpsFptHmHN97A+GH2ri6JKjJVyP5CoXgdD0nh7
Z4h7U5B/TtX168IK3ymV9C5UNDx4GVPMTCPbzWlBfbfNaPUdgff2+vC3XnK+wu6KVuYQxZsl1kJx
lxXmkzhmnoh3KoUNebBPSL1QS991MV6iML4XdMr7McKzAkCdDob430ezYkN9HSZ1fUxLKU0Qjddk
ICNbzJynk/0f5kCDNj38WJGIc5wlZIS+rO0E6x+Utidvx8aBjRGAkRYzhkv3qwGsOVQ+2m1lMiXH
lYMW+yDnowh+t7dEQCFVUkKt7+NtdAul/aYHtEC02M6Xs8Tn6o1fIluizA2Ew2Y4Lq/2Wr6OvSpH
0MCINiNOwsIEXVuvDk396B4ySgZtKoGRD2mPD47wc+Zddsn5c0GKVQR1KcxI3njNH3/M0z1+ClYC
BM+Q+aHu53J7d/mIHWBqFbfke0+hnQ2hV0MRLmMq+nWlcXF9Mu+NJPsYwEBs/UnFPbJo07qUEcaX
RvTJZLeJqeeYIgdT8XnAKlxYTWb5WvT7Ghyv3QEsqeW5HqG0rivDLFJPR3V33nsOasluoWzAi1IK
AW19vZ7eBlXQODGiaa4OWT22vOdab1OQ40F3M/n/YNc6q3oOxAk0gTI7eir6eJHAmuT15r1XoMfX
YDt4JZXd83JHWuew0+IOa4bof0T/O5WimbKjI2CPUZzM9F/1ihaR90v8Sbtc8P/qJtLFOpa0Sszr
tCQT9GfIYdUAEm7ONjaTnoFPdyIqVlyZy7H+fzksKVEk13rCOL3o8+E9zK21mbrN+OXIgWU1+ODN
KUNFWb3S51n7hgxVcCGdt6R8ubxt0sBJmYkYSWu6Go6nqzoF1JGxi3vcRvew8JUG4oBfBa/CvZ/d
eoiuu40TEWaBBvqfWxRJM/qZ4cofrwAInDelvZ6KSBFc+HUCY0LTrvGORXmZcB9lLiO986tG7ugd
F/XQ7WZmUO8mmtfXc/4Rsl8bL6jyzIhM1As6as+US9dJagkbKsYq4CF4t9n40CDZ5mbyUHqjdXdj
N7OO5kV55T40B4VoADvloGlMe68i0Lgn7hOjmmLFlWcM195N+De7p3lQm0z+I0/bGcj4OXRh1p8O
Dei70FaL6jCV4hs4D03L/+M0HIr0VsUcr5uGQ8S0PRT+oJhedPMMi8cnMD49wHF5V59igkw+Hi6H
JNtdrAQY/d/4ofpoTch36kJP3u090ltYyeYRUwL4ZvBjekI4KXQb6DOAguRWNtQB0SbvJJJUj7Ys
PWvQp/Bg3+SfZx6+l3vAjADysnhlOm6PwQQ6NzjhZCcFk7szKYfqyOt/Tn2S7TcjD2d3n/8wvz2r
3UPQN0H+g8jw+jNKuGlDBdknqGwarHJbCiFGeOCtMPXj1WG/+MKgAeTxkksoIYi3QhQTPQohgsAt
qs5El/RxcwRouuviY9wqyGH7weIX+pFR5n8WR3QovKaDziYjrz6l7KKXRcXJz+FmH7xeQASjTcvS
H5RDXcvHuytnIxnElgGqOM/u3J7lqHv/nmA8Q5LlKN3CE+5Sfngeqilg0d6YNH1n41IuEtVMgQcw
eWnQvA0CTy/r4lQZiTn3rKr0SvKVmkcImZGVZb9WmrPNWa3QZ6QKFswtD8maSzwCmYxyB6eFeD57
p8Pg4rGp514oVxXFgKuzBV6Qy294JWCefIszhiKl0QwyXOrOujIDHSR3fKiUII9zvfgllcih7lXe
DNt9AGLjY94Eka9ca+AksbY96vD4il+ba357YvmtL1HT0GKNwsvwIMEqYxfeKd1uL75rHeUmR386
pDXssriaR/S943oNt9r2fVLeO6Pwf6ocTW/KxgMyIaasVkvS5kJcYrtxt29iVYWIJnZVKPrZ047M
GszDYBhWnC4pR46+0Kkj24d9yrNr/Bt2J7R9C33kkNYqtJrq5zxVNirofjIsBbjo+zE0joJGTjpq
7SYe2ugC9nBLh2ktMQTXApQ7sigeRnxgH+kM04/xA1k9Ptxt++76GVKpllCkhyFerG7RYHu/+dgu
lmZVhzJF5+7JK1lL6ejQcj0B0iGmdyda6Czg7B+IWbMojWvRBO6+bsbwASzixiy2kYTtLP53a+vI
pk0wwsSoyGs0zwrRrhTIuu8wqu5lri+DeJwSV1KInHADh+WP5cjZOToNhnnZ+rZn6PGdN0m1rrJi
8S+TvGpdwmykJDTkPN8vl+j6BS2FToSf1v0i2Fvl8gNQ0fdY86NdGw+OY+ukMgPw6SxXDzUjc4LA
1L0JUAQqLYyBWSTUUUuv7Nt8jlJip1Y7DNAVFN+spc9KLkbJVYVmSPsNXgP8SFhPNQc22J4+PV6o
GHmR9AAqbVyX913jwHozZ9nVi2McX0PRklbrszh8AZKKD4lqVooLmXxo3gCZL/99xtpyHK7j4+A3
iwfeSD6xOTvW9Pbz4q3q/0HnI7bBM70PdFySzpC+hC50WDrTVx0HpvMqkCdCa+/ao+PygNkKejPj
q5ljuBzLvE+xKkIqLBWR2TKMYOiSgXQs7LePY3nKp/VAt/LpknTX+ll3mdGMiiYpXiYTY2HYfKB6
LFyZVEMunK08J0iH8wwnoNiI0aSzKMtVPzkqH/TU/E5qy8JJYiZu/kfYYoiv/fEaeaSrrAvGJ9fo
WvJOutDStvnvjgXLd+PB2q9uxf0ZRpnVsO0YDv/Ka/TYS7hED5iFa+CN3rjOZErgRF/ZLPOJgiv7
ixh6hnCd143jgP/k7NmovYC7hZi+VtncIoaXgDxj5iBT2ssBeffuu5yqcVraO1lPbDStdWfwxTNt
eKh/x59OTePkrrezfmNsH56jL94wXo60sPt/99NZNylHIXP9tnUDkoNT8V5PMiPjQJBR3LIZ41N0
9yErIigcF6kIHmWXMgn86JWWKf7SDKrDgpYTdr7iP2GDxt3vzOIk0YvBn4KdiOR4kG4DNDo1d2OZ
hW7cRyAnap82wIWXoV85nmuQ3mhxWGOWHp+u7G7Zh/zXaB6Ot7GAPklGBRolQzWnvXonAs6xh5Uk
fRE/cOC1Ajn5x987OJwgZxSKUarzkZMrSr24kc7ZdTYJotApabuIImglalQxbDEkpTyjtDYQRmRm
1jwAYzRYcfS8ShjgHTvBAxDNonBjruNtyBzwZpM21jqbpb1HnAWwG6ONZ3HWwkGeSMG0NDQqA6up
jmzKlyDvxwDg44op3ilCI8MPi0wqEH44QQfWNy9usTXdjtZ5bXxulXAuPKy6hfumeo4HJGqSHPO3
0igYxzvfJT5GwWVPygqmuJ9d65JXml8l2X1ShfCdeGUwe1qlNwJftbzFt322OaY5WIEFbQglZUmO
jWmevQglPzia66b/C6SVez2OEvvp3I/jaaTRwxqQYavX8KN+ZHXl7diV96v59arm31bjM92Nb/gN
8urA+3y4NL4npDyv7DLk2rgBuoXx4I7s/i+xkhl7L038806THZyyEz9SdMYmxDLMZT6ddHnCoTKO
nFVq4r+JBsl0SOMvky8bUi1NS8ouXFN9C+s0Af/Q01d3kaENVh/gM1e0srZVtrRKf8ipVOu7zV0t
rIdiO1ok1V0seu0sgO8852nN1GOF4kBSpvnr1fNK4DB6TPaKodOJc/zgFY5ky2quO6+lhGBOQvHr
zLahNOkFyo3eKr9k/C41f3kin15jAdp1M6kUZv21ZSqmdKSnrFa1DqYR0CC9TVuhdF+hkDET+do3
wGbxA5UG+gWoy+NoRNF+sbByVnIIAM9caMWFCiTXQEkdErZ0cnJ+VZZj1JcZJmHzZ78g/dl8tnWI
twFqn+5Woz6nafFcIdH/t1J2koJGcDophmR4beJvgttRpnUcqcphRXNOoc4/7cPMQymnKv9pfBLk
0LiED8Uqb/kdltLf61+9jANLAayiWnILvw+0tsu1a7nwqcJ4ze08Xx5P37BcS49sJI+HtmawZ6Ar
iKOUf7jkxZJQwe4i6noLdvHmiMjoOqh/t0yxb4DCqlNbWNkdlflphy5ZdJ04o/c5dq0Rf0P1J+XY
nAgTSVzhKR0WfxnJIak3PpJpZh/iFzyE9q6S00tQkipEsVeNpgoMRr0wARxvZ6BuMe8aYR4j6bi6
pEy96VRqi8O1UPq3YYUaSBMMnwKWqUXT7DUwupddS1cu6tI5tqPQSHaD0qcolw6b5xHZ/oOrKztE
kiUl2OiY13H65ogUxn3lNqukeoDFGfvMZQZDow6j2mQHcotaIx3yHi98hEXmkyCegrY2iKTl60IX
v9FBN30m0sVv2gpHGolZoup70kJj50BNuE0XblpaZeOrKBJHANs0g0CfTUJLSbPqwkV8z9b1OjZE
2RmWY+VNIV/wRPER3fKR/z3eKUWBhfuawbntcfdUlHKPR/ptWDzi8+VpuuzK3OHbKe0NvTus+Un9
Vu63wEgmtSkCIojJCZPrieq15MgGWHr7ByZYqJNS654kU5hA55/4QU3S9ZWj1IIxSvqhNfGIJk4M
KIvzEvUcf+/O1/rGaofOlHh9U8rEVEceU5liMUNsCdJQYLlP658FLDUW7LZiTg1YLDS2buPMqgDP
OUJz/RNTpkgBWz+F7+wmOeBWFItLa8zNS182UtZ8r42dnKk05AAIT7M10DMTb+7138aU/0pP71ao
d37r18rbCQdE0f7ADx8MSl8fxWxdU5hQ/rIMz/NLxD/6Yi4soJN9Ft8LezAGbuKaFu/4HKvrGAaW
+agp3uEzBrkD0afQTh9sZXZ8hkBRE/0Qc88QM0AkUn5MPc1cfUahn8Fi+lNphzYUccCD6TuOU88h
SkfeFqtl9QM2tGAmdA8SzixIPwsGmyTVYLzjMupEuhTfKp5sJAQrKxnfAfzK4QkFTRDmRhwDNlMP
Txo1Dt7WT/1PG9v7VepZXk+X4mvcZdiBbxoEOuU/MXDz9FOe+4CFCP4Z+xbAiiGC96wYvy201XXj
ttNK9lDFKZ6dQSGVMW3qDiYveTIDAD9Su5k9aFJ2Qiw6M2WR5QSJ0DqsW0GI3NsMu6m0IiIzOFCM
/XH/l92vQx0d6GDE67Zwv6favsoJG/MDOzekDo6qiMiZT0lEIIKdxHf7ZcxevqHTvhHrlCnQsgyj
lIo1K8LzubCvYxn6tc/IfCWqsXk1FI8js/l1gDEfPkh3QCnBB3zuwll3ZGeX/5bz0Z1ATJxJ+cO8
20fHV/Qz0lVikIbMJEw0U/ej1hMPoCgsk+ytvGjkEZx+7A2kfltK5u2VQ0ny/2ZlEou0mq9W1UB+
W3CsYLhquuSNtRX1ijcWnxbR7DobmHmFs0Q6yf8bfvAvDL9yawpCwerUBC4=
`pragma protect end_protected
