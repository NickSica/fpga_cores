`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
R1WqgqFekyFBf+R1EmSjRCQxUuOx6MT9aQyodTNNebOe0CK13nDxh2Wir1luIC2E+1RiIa720P7G
30ynEHVRjA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KNMY+1Jln0fE2Hw6EJV59uwRAjQ2BHIWVdMuSpeAltv11pWP/JZCrd4z/uZcVTngSRY8jZzhCZTQ
WJ4MxCfVaXUWBZm7mY0qLw6qcMnyzincQFakqwRdOx84IckfsGjNGJ3OEjUVkf7dW/J0o6KJvGRq
A/P9gVOYmGcnWb2CkLI=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
sL7gG3oizEXkzDHancu7/45cwKfdv4EnXAdeK54QMEX/eoc5P95Q2IxqcI+tnVljSH1drXWj0Eb6
Of0W/iXPKZ8OP77HA72GpMs5rDnQtlgP3rECZlxuTJ9RMJVfJzzO19m/vMWeqMysX1t8PW29rrsf
0Tqwcs84OG2uxBTuyDEWCBSCU7Yk0aBYU4VmF2rkELqh6jo2Q/udlKIUXrwoYSdX0O9uon++5ahv
mjzu8SGK6zkA4uqzG9ghLIe8qBE6KYXQuzvdlMdTVdy8eHbCbzVTNoB6j51Qlq+S5oMMSQvxBaRz
DIAN76FuevwCbX/XKHESsvee5Sen235LJDeW6Q==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NTwqMfOwske0aroynepwGO4Lz00SLylJkTISN8LAcq5uE8ZoeT6aFHS3yIuZsI6EEE3s5mQQ8Cob
RXh00Ler2BvOA4K7lNGJUpMzGqJI7MZao2GijCVpdWL1r0vSvaacAIY9nlusgQmU63NqWs7cQx1t
7NMmVlpgPTHr3KxO5lMNWR2EuXJ0I0zOxQbbrTneEEip68PBGwJFyFdSjQNe3iwSj7O0u1NlI0nF
01F/RGHelGngznubnZikT85LEu94GTbx+WNlMlaxWaxuIaRvhH8UG7MPhsxH6x7sS5ZS9GHBkFDK
gyo/ARDW7a6331M9HUgGOcgw3trs1/Klf0nskg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
F0eZzxJQxbI/Xk9S9oAxZw5Tpi91CrcqL3BrQB2lyqn9Vl25Garq+8JIOwcSUfEju0nEdI9Cvd5l
ooe0NMs4K3iY8tnE+FiNZhFGnmyV5djhXaAeRPiaySzeXAc0nSnoahW36RgdEHyPbHBrMfq1pT3d
S/0aa8cloJNV0EZcGFq/QrhQOhscPpDi8uk4IV75ihx4K3Y6D/SPBsIijokh2lVOyPsWt72NbpFl
R1J6iXczzSEND79HNenePfXgQ1Sr+h8Z2ujGHirxn/++xFCAHxWZmhGcFFwVO7AI15b3pfNiyQF1
2SACCg7/b/5q/JpHGBLoFY5e10UGMoGkaXNq2g==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eShHfvBzKaZ/Wp/QUxGlK7/6Td59dAgzaJsrKOgtjc73r+sFOocLpKUK8YR7XmM0pkfLOBkjrXYq
jGiy10qSwBo8l2eE17VZo8T9nQ0IB2FFGgVl0zNGiZaKSzE4a7K5so8c5gtUyyVlyHWXKqYAj6Ro
NzUEnqMqJPppbTPQbvI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
VtDvfrNdg+YlmytFZV1nO9Ch/hNzGllGY3c+wOLUGxBvYhloxzDDcAB/7/ljwrwghZilvxZm/DJg
2fzdltt6rugwiyCDZPTj9bYqZhAAM0bSdp5YpZP0gTz8EvbCxUo8+Op+ufZee7A2QX4lG973f4tu
FbV42AkOjECD3RCU/zC8zhB5kCMonmYQSEe1sGWBe2+Ga49sur53s1VC1GSUOY3PQLHNqtwSq2Ra
owo+cSlmwu7mHpq7nDvHG8vWLm58VKt4pglBRfC9BYdbhmSQeWT4IcMsVz3wzwUMY4HmFkj+0Htu
JAA3fKLFH4/svF3ilwX+klAmiEhOn+ftw2QOyw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HHgo2A7au8S1PE/PLf9TgssZhqFUk1LyRHoBPoQd7KZOhYH8iTwJV9W8hjvxzC2Na0peqSJ5zF18
7DRfKJ++XfNw8OtnyxfjOhMGRjIzpk9/xlZOxoCpZPFsl6WTW8CoN0RLlh22HuIAeiFQu4jBiY8s
f/eG3F7z8aDUIS222+2y8Lc0ifWDx1YbNoJritsavlDA9L9WOwq+EXi3pvUCyXszhqfkMn1JVCVR
qUhUx37i3M4UJEKXpk5rfAol3dwNa+jlOtqwiBj8/VnhZxY2i53S+bX3OP8N1Zx5wRoa1UkpaXLd
9XQOggc4VKKTgU9CJZPlRk8FrwN41qv2G8xfRQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 236256)
`pragma protect data_block
eeCl3Hcc/V4mGRBHBrnlVPxBhqk3ItIYIjgE8V8jPs2XbHnEUogLwX/TbEnpNrebRZEBMoeysfzj
RG7bl1tmXvDI9vMC5FglPwWlSuvjTHCSrXELYGZgFZDaijhdoJR1Ht6du/CzpbqZkYe11kbUQbEE
vcJhSHzw5gf4zU0LAda7LgRybXZB4WaqogBOLsoBE+sMig+EUJJXpvEGSNgVW99MRXuBbCk7++B7
fsldI8QdOcNbpOqqPSRLzbAplxpxF79eVwObXRtIZq7dAsv6cbDdSObFwI2vtqEQEAWZJNC8Sf0p
U3AcG2hKmS+WO+whAkjrfeATQbOESusmf6HqgwzNPp2ebe+MucP70be5KFLZAE5BaEqLNtdmI5Nw
XSeh6Zz4J2oz5396AHcTJTbR5UvzbEe2mZOlpGakK9cGaBsnrz4EPckPjKGesbs6VwT6qCWwG3wJ
HliCxmc/BuAH4MfjvyoTEuhNO1Hy9t33H5nsZuwsiUTabpWGX/7fc8O384hn88MW+UmELNs8UoJn
zbbmoD25wemODuFBXMuCaUjEWbFBIjg7zNuOU3HNcDYyHK9EFceU0zuwidohSCaOiOrCX387EfLg
cZSwOV/R3DXunHj1sS9eeQ42PRObHFw3JGOO6R1XWqD4WJkGIYXMFLPbuqoOf9KCUOvOCQt4FVVI
q00rvPgEmKsvwXGSsl0D1AArIdELox3TLAQNDBLyjGlVyQWahXQnkRi8f40AKS8y/xSgLVmAK5Gz
ynPSkMKKatM+CTOdHLLaZkJ9bGlhQHz6CD1rdo/8iWb6MdelzKwhIm75rU55KycXd3fZaNSEsyyP
F1kWykKL2IgiW+jTOjGUJy2KgskHRBpL5nRVwHCUg3+9hpnXecG5qvPQWbi6CMBEvtd2qo93cspI
ohq2JHEVRp7bzR49fYhrA+8/TYRGhK854AoPph1jr1sdqjvvRn0lYMZsq27ugeuhiIHCehvdGtfm
5c0+O25u3eoEbhpgprVOgELK7l4KsmJxs7n+rPozkMInFMk7pOmItAWHS93zOAD2L4fBtov7LUwW
wCvACIW6cLQYq3KNmvG8Q4TuQ2a9B3aZssFsf0AkGGld6a/tYg1G8s4QcLHgZW7EQcfI+x1ok5Xp
gUO9NiSKTDeLFZoOraItgR9uvZlN0p1nc/lkd7ZIBxRdz7C4JuTmT79hu1K1pO2hR21r3Pg5zMS3
av7eWCTEASrv0TMxMcV7Llc7vj+vTwenGeeGKp5YMOnlxJJthHNhJTM33ym8tTMhNgNSVmSsmlVF
FvMzCF0zs9IJlpcf2KA0moC9x4dl0/sIXddp0jS7W2UYeZ3IeA/yErmA9s4ulEaykHahMCMQaXo0
5S9cKvqHvZSVZhT3ayENEVEYo8dCptFHc0sislURc/3GpukF0MLMaGwX2qMKKzGs+G5qW3ZH0yh9
xiqDasi5tQ5NiPTVTtisFuRRmOSzJDk9dTrVMOnGyqVa5IurlokO6GuP1xryQ3+6eFfjUKemZz8P
BeZ8AQwCZvpv7ohMCQFmPUuswe/kC8qEmrG8DKNAu38riteKM2ZNnYfAjXJEb9/SmvRypgTgq4HU
y8MIRi9kt7vxw3BPiPFxHc2/Q1QGao+r9lmNONGTRrAzHXTeIme+O36z1gLQURPb4dBaROXeMo26
3BfXrAdgdEfZjnxVzX2FUmtnA8tOXA65dGzOk1V6Ghi3leriPWcNu0g1UEB1qcpRxww4W3ePiw8y
Eurx2bzrz4kBEQ8utT/MGKsqhdKb0TDmHkfnmta1+i/F6CAQIxSWC8e8UfQgG4jxqQmoDLQvnM7R
6kI/xSHA/knlyVj3jLcZL5Xp6woN9nNC4rDVyYhOPVHhZ2nCXheq4Qd5g5xF6SlVNE++qtRhJU4S
3xlgG94G9t92RUD28Z/gFoi16wY2MjUBannnCMXW9j/cRc584HEhuzTYrkfisePNJuk95Jbe+FNY
t6Ck2N8evbZL7WUYuuEszupkPIp0qSAjhj9lC9zVYqvdxUFgg2+WWd8kP1ebUR2bKx6CgCz1l5KI
3yQvzG6mQsChomnw569ts/ma1Lz58VtJ4ITciMGNWWubDCQmu9ZMdsFjiI15I/fKNPbMOIvu1Rl4
TBFYqAdZnYII3mdWoiHmhBw5Jm693ajPRX260wmcb0QqndpKK4okLZn3+Xbgdjtv0Xf3S1CzawH5
mUAfDkqXjwY8ZB3JnIjbJPNM+hppOYNu8ZcaATxeDQdg7Qjc0VGK5qJ9CCCrwjZUDFGz5uO3Pd+3
SVe+pW51mPw/1Vum4NAa0cPrLJXUd+KRv8e0JMlJHEI35X3AporW1xmaeRf2LhssQ+k3wzqLfu5/
oWPw1Md7s1aeNU97+0fXr/p8ezd/vYve/woEYamfvwKZStF8eu98Xv6BKQfkBy4r9PZPHxBCfq+L
OGNui5sqh2q9xC908CCADdSzZwrEBqFRXqoq1PqAtmUuD9Uot2AchhISFY7PvKxIfUyXQcl3tCN3
NTdwmRriNzfahpTGCgBN/+94OOxO6bHhkgNaoYWuKKkWaLRG29wt+AUCemzjNmkItxAucj4PPUnq
OVr//SokjsWxEPTHjE5PTSslA3qCFSNmWTQUH6L/AJskWztT4mcBdtgAz2NCls/x8iPBqnH4SK4L
n7lKzlOI8UzXxvfyto2bcQkcOHgwKfyZuKqsLuLwZphgRCGuqIY0/SRNe+rMuNmfcJycz8j8kvrv
XK/yF18KqUS/aG53zie3ukHB9UBdtyc5ALNGd1Y90FNJSU7oHE0t/4kBaaxOBiACPa7g09D8snoq
hX8YfqrtxVHmyBp558DEnWy9ww9xORwlrFGPnocQ/d1DgZbjfaFTj+v4LA2ySBgn4wYjBZXKge3E
HqrGaMYYUGffIjyFq/2q6jwQn+SC4KsoqipHN/fv7W+TYokOLRd4cteASoFUgvBtyvbMGFesmpEp
8wlYP3tuuDn3Xlrj9UsUIsVea2iU0HwOye+e4JEQ/7n2nHGC1kn1dfF6I8qKxr1S8qF4TeMG6ifE
AB7EM0PofKdl8liiGteiohOAYtZ1wrAyXo4X8vSPQ4jeEWgfc07Lwgtx2752js10sDJz+cjPr7gl
ELuTMKBRTMUjDeJ+bPl0RQeGNcYk0L/ykDh8a9bBWdm+jXSkW+ubHmM6Zj1ia0TYTx98soUG2VMh
yI/h4/kYWBWMJv8OBqG8Whe5svRVNT0pmt1ZSH6cTeYMSUhyhBas/4w6GXVGFhuzQV+TSGe2/sG/
pJYeJo/xXGpnoJmobGuLUuN2auEnFlim7+LLrzxguTbxvME4aEprJlSh7NyY27mZBqJoVWBCSnMJ
8HCWOhhDm4UETbVTzInGf7KWQ3gL61Dzsw647nrmnO1ltkoeA+zvo4qWxvo0/OjjfiOsnhKEXndp
8IboUWKiZ51mBIVrpsN/a1+YLXwp3cOgaCW7IBjBvzkRU5LNtvG/lrTbLWf/ClUu4f3yGh4O9cSU
V+amz7y16k+abgQBLnzSJZpGL40/OSxhGMH3GmsjzWCKlpPml5xBvQghJG31+eptVh42BPewnxsb
bA0FGWRdJX78XuCIFA/dcRS9lxu4y3qcscac59hF0FKU7bCcrJikhO65/+at5lqwN1FadsHQCYC8
gGdTMZR6LjCgscP9pvvuBJSBvheos/Zrr7sOEYSeK48ieP0mw9487aEv5HOjvfsiZHOx12DurEP1
CFr8T1mmp1y8PbbGfQppw3VsyNfYMdiaLAPylXEhvCHfeetbUTdUZDj5eom0VY8qziGI1yl5U7QH
Z74AueZAYAHwR3Qoxq8Pb8QFwTDdgYO5yl69zOFD3Xuvy2xfDsNhF6I0UbcRnSrL7KwXy2z0P38L
/mROS9NRmiMDIFlguBevw9/r/EnTLmSMVeKl1Z7dlRQtGJAbMuau6PyDNK0dEG2/9GnG3I19mHhA
g7h3yzekLMckA0tFaUX9aNkQY6W+1snE9Y7WAiqsD+shd3q514jPgA9H9kS2IJGLId3lyZJNJ/L0
HLVtDLgrOEGfxfB6xlP2AmlFoYXQmorTm6Q/Q2nDHmWGY2G6mga77oTDzpDZxlDyNHfTpDJyg36c
7/c9BbKFKSE6/hoSlphHzqngAK598jHwPCrqB1qWHQfKq6D2YdrQ7qASvfvChTEHGteRQxdUYjni
2T8FTlHcg0BmDM/FybXK2MhjWrikdcFCytzrGKm/L4zVww70ulbzkAkr8U2OkqdjZRDif/aviLHG
1lnSlIs5qiLQ+R49qi8YavzwnoQARX+moadaaoMZXftkF+Vqy/6iuWwsF/AGaJxF0wfZ51W9pBsR
3QD+du5pNVVC3YUwrLXeZ3IlyJNqJq9M/b6Hqlw5Ws4Y7uDMkkUuqp+lAUGdSK/PFpv2nDRPFFDb
gozdebHaJZbMht+UBEWvON3zC9Isiv6drm5K0NB6GdQhI3LMoByq2thJdgPOxqRmBmjWpOA6yL/d
vK3rHW+RAzpQj4d7wy8yJGZtxBPWw0kAQ7RBWMOPInhBmT5Oj5mYVcvIdnD2pT5TcVqPaMk92mJC
ZqNW/rtJgsAv+T0bwMR7Eqapp8v+YEUwmslWnCDQ8EX2XRstNnry7XRgZiU3IlWP6Uob2oGSf5GX
qi5mB+ef0UvfRpyexXG+28gGWQyWaM9tVi5vZ8go83yzRpsY50IP31EotMFgAbwoTk5iJ/BiZOAp
+WMxjcLspAEN5BQusRmNv5TOc9F+KXeBcB3tZTo2ILOh8Ya/RsrsB9gXqmRXkmU5ks+RqgkMjfFf
TIrPogtJWupECqMMMHsV/oDSdKm4tkwwiaVp5ORwwwVAQQisB8UY9z2RQbWX0v1d1sTovUOdoMNK
JptZdUNB7/UJ2+WPilY+87JHUQr43S1lOrQKskb9cZ5iLbEQi0AxvXJRZBLAXSdl0Z9EyWdd3J+j
p4tjsUITXIGIJ4lJhj9eBebm7jdGnfHJ3O280cOeqNe7rw4oVt+9wnvQu9sdcZ7aOzw4stZnTIx3
dgq7D/pu8nmU3vg0M9GSbwzo40evAODl4RJBTvglVF1BpyHTbnMjLgMzwnr6+WlcZb7d/QjspTFh
WHDU9zWQ1phHfJNEmRSHvQtvP/fmfOVYArWEGl6Fp+BrenHpgA2SyvKRppEHMr6FpBzH6wrEs3EG
zV8I7BogXw0ajnhd2C3KpniiGdMnLKY7PjNNSoaj22KgLznak2IhxR8r1FWLv9xYZjIRqrI6janl
BONXE+Dd8dfF1QbHfSB6OzexPKNgn5blOiKWQCIisKN4Ce9VVfQCZX4334crbEgXqJ/2GbjKbVHI
tObGNOzyo4wzkV0bYUj6qtM+Lfllu0j1yFf+JrNX+yXykKzw+jJpWkjMxWzKhmyugTYdGvUR9T74
rq+WeBhPxjY156WbfePofylsVrASjuZ05q5rGc6h6xg9u3edV3poQpbuL7Y7zsep4bu/k3sR1sUr
DpXD9zBtNqYjR4t9E20m2pip4z9WjszJpBwdzEPej/T9+w+qAY+qv1L/7mCR26WBXTyvPwKKpW7Z
u7tfrdDLMCPzUEpiGzh4CsR0wmv8W60+21P2HyuV9Icijzc9Ih/2wqW44+QvpsavfVHfk43prD33
qMw4Z75290qe/0nlXIgFLsjTcbsRDZgGrpbTKZByvSEYMjViKX54FwtuRq0g5iNrKaMsA1pt5LhJ
LWkgharmQ1+XYMmNM+R+O9U3iix5Sq9WZY9oyjYtMJY9K6aPOWNxvz9ArNdNINUxZdXNP61frLvt
mxsb4Gh4pmxHA6fKAeqG7XfDMOnlDNHSAumCXm7puRlM8rjK44JeZHxM40g6gWOyFHycp0Fa/QcE
Q3bYUPybGv8+vT6TlxyA/FkBKzmWKAlNi5e5U8uHVqQ4wdwmgxBt5M/8vcyOFfVEdCnD/BEANaIy
IFoY5EbdnYXRl0OnYZqb7TU+a5fJ5dkEL0KBnrsvfcMnkIhrl7Cg0mJOaPUQGkWBY9TSC9S+AmwQ
JAdTKtCKMAe68Too62NcCZWxsQMA/dX62CkTa9aMW8IRmNviLLySkaWInuj4BE/9KB/i6i+VPBo3
SRvSZhWqh5XoPTLtRyfaouvEKDq5vZOZywEjRkQrhW5Kf5o5MIFMGRpB7EDnrayrIke2Qk52lNdT
EtM1sigWUV8KaRAvIa9YsQFT5L6GgBz2Po/uz8kSFu3/lhdD1BX03ab8AcPs7zt9Gq6W6kQX8qyj
eGRjKP2YcS7+fJRiHe8h1ibFxQGgW0vjPH6jxhBXMCZ4OdSup1cV0bUv7ptQzAQcvPoCJPiGkX2k
z412BachcImGEL2qdTNUQx3HBcAPp/ECb2CZamv6iUwwspirgoQ0p7pcv0W+FfaBc02MtnBhkPuD
aO1X0gzPZmbMNU3+JlGjTzHrwyosvcKgU0Fni36Ta2z+TwP+JgnjXcEEdWV9ZzLUXG7KAuCmAUkM
70IMDndZ4iKsc5wJ9bR8aW5WKhvWMem+sFKghA/jIdV+cs7x92wPBImtj7BehEcKmLASRkqQy7M9
CdFjkIQBYQB6XP6+rgc91sNED1kYdGhFtTI7v/iRHDNkB4M/GiD3cIbrTlM90fZXMl65oRGIPBjl
FrlHe+htQ7VYw1iYFNRa1NmJVJKrt3FlKZTY+d4P1EYpIY5W4g4ylUDTOgGRoEWHgU37n8c5XAMV
vZ1wualbG5qZpVf2yEJXmw5qYJhdW/prk38rVX8vD0pgRTl2x/C9xi59Vh9FEEVD1gX3Hs8cw8eM
Yk7ZUVdmeRV0fy3lRGq+gfX7IYbW2hoX1piXW4DqGKYE3vPwW3/io03gpi5UEITUDPQTEL/UT8ZH
Bxi31Rs8mJrHH8FrlGPE+gWXoaZLDdLVR9gs/xI4Xjgqh5zcpju5xv6Wv+1Hfd0L9gjq0L6UT+1l
FrwcNDLJTuDc8qDB0JuD71lVk/jPgoyI4PmeC+VoqutdGLkExWchxl740CkbilMgpcByf+d3kxSn
dWoH1MGydyh+zNrJuTbQjG7H4jebikgd3RWVued42aJtGo0nlxaKYQ681BjS6e96p8rW0VygL337
SBmyj3Wx2KYf5jUhsC/UDapwYsstC5QGDFcjC+2sAoISEtNQDQE9drof5NWeAkeeIQv2wkmt24uD
MvgA7zJQQSSG1/HQ8HdD1upAR8SsQejNtLK4qaPxapI6eV80zf0YQJbERQp9WJ/zLDSS2UTrLR3j
NI1Zc1w3lo6JHPvDmLDoIw5xEv697jdr2a6nQGCHD2weRhqDAbH7jjz05K20GzWGNSF+7TiA3y/C
FSrZkGlexDl26P8kJmJBlVssUD1dcG8vI+PGREjpCO0U1Mi1ipH831ZSHD8PUGreCtpkxqYsxymw
M8YsNc+Nlx4Y2cfNvZLvECJs5HsQ1WS9ZbNREB35KToXtziDFN88eaN9BThOtse+/QkkTnQans2r
T09te6z7puaodShB2XdebyK20oDJ6akcXgRkDlTUejHFENwDNP7t6uu+ibaapRmzNcQtyxnFP0Bu
yhVEjgzxVrZ+VcmHkAwOS9+DsRgqIXIdT/Uxq06jd1ASxqDzUFAUze01ERkXCD4K9RGZcanQP0OY
WsHELMqbkJWjClNhUX+eUufkiT4/WOTZ0o7vHImyHXsMJDJbDCLbHyN25SC4OIYkFMfHRdN8efe+
zERck+DTlI7SDaOTIGV3+e0RWmsH201UHwED8Gbt2XVnL548Xq+5/K17JwyjeWLCT8zfMTDy3pYs
3TQACMRnTPgRE50T7IJBIkUmP+hQiUSM/wFylmIEwjRKMxLSPEmOC9BtMAa9JIrpXRsxBzsxZpOE
2byxLTQNwBic7yoLekwTE8G6/DVSNYlC2YQABKHbURCbI7Wh+SshWqWF2DT/NDI4njHdFxLHpL8r
uWzhbBuuHZA1yO+u5arCbAvHMSsNhmzbWXXxIOAQcBENy5Jz23keCoYPIwvuld6cIOoOOF2eJ75I
VSGO6rKgkJd7b2ZIBtFfkp6//7dwcmYT81WT7WloJDI7U204t3foxtOLcJ6mmlkEajryminnzt5I
PhoyWsr7Nt2flmbc/WHWJh5mpxMdZxFkXn9jch99LUIlpfT3sXLjmc3iZ239CPypCroEMJU1ZQ1/
x3u7zKB2qsX9R+v3l3tXmaxXwo9Q0yi2r6eTTk+dGNzvMGjouNUlsVddPnHPO++pP4cuSzRAbNlx
4EHoLvtdCWzyPxLId4qFqW0BJq2DikGDGViMDfzgTr3N/sGwVaKwdDa78JF2o8b1Iu8LX5hcIXQe
euxaHneDd4nTkf9t6fGm3LKXybItVPPhIiOw5R9USceJMISU7zNHZdMCpiIvigTXa4rzuMy5e2Gi
EmGD4MhLSMVM9f/c3YjnmMhPeLMcMFZ7Idhxefgd6iP+0GPABLERTogfUjpC8uZHB9Tg1QkCLUF+
dYVZXkPlUfVD0VqPPKsA8sarPm8etq2o0qKXq24ogV1+jUONMjpDI2YCLRtp0FIuydzY6PSK48Zv
7T+qp/m1FLiomwrMwSYSvw11aUDCexGVfsmSvH54N+mbWf87P7AyJf89YPHMFT7mTS2vU94ZqgU+
ACXWCX4Xvp9lJhPTKPWI6XRnG8Z1rMY7uN2srtPUj5wIg855bT3q6Sce3a4ANUJxKixrgSaFfpYy
n1kQm6H9VLIJwH4CRVCZK/YwcYAzl4BQABq6UFF8xNCGzVL5QWnz9h/5H6GpmalEKdNuIXNkcMZW
XJHQEIorUidOfZ2GxpHZuShOzUcy5CztEOQKnRJYYgm+0areCGmOfqv8HFmRFWczuDfB1TvyrSys
k2Sg2UpAKMmzIIQlB0Rkkm0t8fJavvx9YBXT1t8NnBLCeExX1Skm2QvYy2OtuIJWWyM1/1RfFc5I
4W1eNE1YBCs2vQDBjxcZSGk+++CpNMvdkIDUFwM1efDzA1K7Bn2SEZYXjuwkZXR+2FUhyH8t0ANP
DWFMVcb7prG8V7fW9Aa64EIayvdSBJiXeo0V/zB/VtCG9Ov9quvySghzZ+sprfOdoxKLqZIvYWQ3
lSQ0vFCQjb9BcxWPHadCq/yRH3GD+rhrJdHsQMS2vPYl3+0Dt6JwpN01PiND45sljBDcxjsh/hCu
J/9eO2Ie0OtVc3C3Mm7pjrL0t5I0kdeNFFiyATRtS8rCY2Jl1/BtGBCIkAdzt4L64wlE3mi1oacE
f8MfPYPwgQXRTMxGkxHvOY4YluS5myNcxkyza54rsiZ64AHaPxDe2DnWQNjfMFWLTCO4YQlO89x0
biNfa3a37fRktSu4Y6NBDj3Pw4VmpmZg20O57K/nNKsgDzcK+D5hQqZxTvrukeTVYBoKZKmEU/3P
8yjcaACBfuk5F+WaK0YaZhb5BmS2QNXCj2Lb8Od7YjizCOMvf1QmA5Ir+F/iAjyYnvno5cZLGaLD
DjFtE8ogd1/w2P7XnbOp7qMyJ8Nwp1QJJOwon0uD7MYzeOECL0+0MyP1BXLzZnHqk9EX5gUMBZFF
vHYZBWg5RORSMiQwruUKemPIGy9doU5WQvi2hpN6f2Ukxa4+vflrAgmReXGptlneKA3BM4yDkIhl
aMVdG3Ina8/vsre2iT7bXYjjVsgQZKv9Ofb6XEp9B37sR4k0bdrWfQ5RDh5Xu0RRrOZmlz4XHkNY
Y0OdiJ8CbZ2lqS3fEz6qpdZ8jIqzZy6fxkQwIil0vRdEYxSmizRke/xk5XI5DqMLsycuaHUclqxd
FGscvECKKOp4x/jT5NRtxRznbiOeRk6B0hP5Tk+as4m9qeqC3mXgwf16BpmdkXVX0uhr/VW0Anpq
fwRf5sNTvz/Lk2+L0Ik2a7r+v2h9CYERuGfk0i1Gb4W+jVnV10zNL9wymq4dk/olNoOFzM5XFKc2
2KDEat0bmZS3jdICxuBpy+tGwV+u+wa1r5g7+k3rzl8DV0VGYQBNjTmSDxagtYrLLDtfX3hHB9dl
k3ZGUElPK5IWVaD8Se9LnxwLavWbCmU7z5KPFvIR3Vo7x8ezh4gYBQYqwsJCKbi7UGTqwktrTJpd
AO9N73MCoRKGa92Tg+TvJKymVWV01tvF0zVNgtAZXPVRkBtCv9S39lgLJ81dJex7udOq9wRpN6+j
J6XMTAhklM+1IUip+NA6omzYgqJ8e8iCDlQH/TjZUgu3j5ScsRW8cE08kSzOBUKoLniFd9Fn05ma
gVwNifCXzzpXTZm9tDp4wloqXUkL4FI9fcqfDtMCLbYqjFvhSd6iGdclGCCMAYe3sMaCYQN3k8JD
GYwHbHzdaX2prOnhPPBsoe0eRZeUlcRuO/QHirkzpbrnTudjd2EcIYxi65PI9Ie7s/aeR/rKOdgJ
1Q2KybbvOs+Y7KIhO8xoCkkmdDYQd5eFLoc6i9EVnjkd+mPimmUYUrmHXBSEEbrP3D0OxlPNO2qm
C7hIzWRjSnBGE3ogDIF+kCAd2Z8CfDPT6No5bQg4HU9wz0ao110yhjvkYiFWYjinjs4UqvB9clE2
O3242FH98LCNJcmryNxOruRHNxrDdXIVWQyx7F5QypeIGRRtzKzH8F9dIeyymdmvZj2P8vIebFHU
5+I+9YixM6Zg6SHkzg5YGedmlVzxwiAD/UEisJWDnkmgmBTlxsdf5N6BG21Q3JA9EAn9ot45hUNj
PWNPygCB1bixhIu+9P/NIhMXkcyWV4TKbJzVwbFaxm4y9GRJ6Y9Ke9ySdKwScSQthA7lvrTVifZe
hmg4ASkKDXWag3yW3dr0DwvCX2DZfUvFtT60Iay+8xtRaEDoEeuW40jVZojShiGhrMMoxRoygsW/
vTBi/Dc77pNI0GFNaCOiUo8W8Z3glMUafhb04PSXixZwFgggbszJnJMhyPQzF9aIFdGxvK+5b1ae
wfagS+y7mpsdI2Nn9drN1BIoS48dzZzsnFaGxiTAv1Y76DAiNIrHA2d+Ux/6Lb2hZ4ctpGTNuhqk
ZeDH2k/tnyRFjyR9VI2WhT2+4/VluO3aUdHFTPMBxB3KWj/JDIRGjjNd3Q7SkNKV5ObXFQ6B0cb+
1VqeoO9JNboqKnfnolJPAG7LwS8LRFxiOFXWysKPlxpuw2o7jyX/t7bgrXmajr7dLwPVpG/mYqXz
l9dlTXpiAGRd3SGj6xxGRjJ3Y4awP1NNnYMqxTlWZEbAYC+58nytpBupe8Y7PiWe73vhMHUbZD0v
b9FbB5AoVs/o16FavnOrpdXlkuP7H3o3FROJjrE4hfYqjfw6IoQqNcdhnlraRL0GFLaM/tUKdXAO
9CtPUO9hCREsioGVcNKF2JeuqM94ATK8X66ePWBbF8WNbKw+Lo/8AU6ZbYNaAek74BFfZDgt81BG
EdSW1Q+fl4JprVyB0c40n9oWKlEvjbkTnsG7GT2BPbe4YJ8OgfQ7MKKBOiXvxk7c4kMHkdFDgvbm
qR5wC/3LW+Kvy+AmvoFiJVnFLeoz+f+dpEUTPjEm9gMRwVuBf9XmfUfXVIo1sYPAorKdku1G7Mlc
SuFeeHnD03v47nvHCd3m7Is4JU0ilc9sSlPOA6mP7fPqmshivbS/9jjvkNn3ZHjjMjyjtwGZPRsn
mFi+qdgnhwvRAgxdF7of+OHaY11M1H1ciR3SsSQF9YVqOxhXe0uqRAmuBxj6fw0mJouLeirBlnTR
rJqbL/kYjU7BZuHbuXpU1I+mIBQv2gMYPrKxelC28Wmvandjgu6wVrV86EAmIY9TRFKb3afS0v3Z
lECkrMC7WG8EEECjdhO0Blcahvazlt1UWzyGebRhCwz8bJB2E1VUKZq7ZxO7Fklr0Os1nWfcNB1I
TdYTkNTj+UaHnTbQft2RuQcnaLGMPj9nNiREGr7qFUPHj2fyOYPpbrb7DaV4c8f08ZmNMTqCqXkM
CcN+JJ9r9pKp7lw5NFmP1JiE9vXYFPDJsNlQz3Mo6bpRWFj9PmhsMy2sEtLauDBwWm2JrFYkklYh
jgNeM7Yc6IIIZiywRkNDM9DV+oO6g/LROTB5Uv9ghHehkKzlRJiwgiajK3XKwBvk9vLG7+VzWjZs
HHXuPqzckFXEFPUfyu3sGhnk/7tgHAgG8JGJCXu+f75SG7y8m9+VZfiw9zpNEXFx5QR+VcBcOTiy
QO3NBEV+p9C/On/ZQkjhQ8QLuA/8dxKYZx2piRuAOT/QJJEiZiXxmgI+CANsQPC25R9YW+WlP+aY
XtcemgIFaLcOyyNyRKBIifJfL3i/jFWywm+xXRVTjFdHi4UR2NO7Kksf57z46OJ9SEsCRQyt3EkF
JCVkElnxSTLFrsNV421P11IumJsyswWC64TMOQSfydwMS/u+aP/d6uw6RbeeJx7YwGmFBInKLKOS
5i1gulFixkxBWChhXlGAinN7eXwhEvc7KQazouzvO7MKZbORBP3uiN445Md8054TLIsLPiRRx/Uw
lPzZgxDZiLL1S6Zf7p/AGsfnIY40DAS216DyE6+sx81s9hGFTKx3KAPYFlk65x0LoAyu1L8y/VZY
H5VffWg/T5hcmAAu9CQfRPbfTfGeHU8TPS1Vi1AvrQN/67w8HkXkk9+4o9zte7keFK6qWlD/SQP2
jBS15DdBfcr67fbjyFvQG7fdRDqU6vczA0OR21Ag9Nf4fEluASB0mjz9OtBDc9fU8NzdKBxVrNzf
rVvfi2LRfLoT1fL2SrI8P90f7MOY+nZAOvnt3IAooP906ZJNj+dyBti7hiBvxmnEDC1V2lS+TPMc
m/2N8W9vazPOBktmmArD998bzSU+s/Y3FHZ4DxB73mFVsHQhr5of/1V/j7goGvTfRM0hKwl6GjqD
4TFTRypI9YaEyLqn1nF8HFp+I4FuWDdwh/7FT+WZDDn+asjhthWI5YxfwjhOqKYqJyorN/jBIsmR
9RV2WXf938wdyc72ZHOmW4YzO8hiHTPYCi7MjccWsLmMCjl5NTppK/28Xc3bc4lZwFe6scR3lxfm
XVcGeFui8mgfTqSHXEVIGSygC64vsk9QJ1Vp1c6iAbc0pSg+btSbA2sWh64Xs9fLKfxoLNmqtvkj
CPo/RxrhiE7GVfBeKC71ap5NodRPmvSTTmiBN1je2aBN3YFUiOa5QPN4cnF1iYo+9VuFpeQlalm9
Oilzo9ptZVQHc35IKURo+8XEPRBMvbaS15A0DPgWIh9Paf80HGACyO5W7L5sbtcJ26WzN7YQOyHd
C5VQJLY1XWulbjMhTE5pdycGvma2fJsvDvD8G9XiGpm4DTErJZmNvH/5r4+1aZA3JoY4GGCeFvo+
59n0hd8F0NHOhDvs7KpOxXQx64ICluct8UgwQpCJAVfJoDN9LBOeI190SVdzAdXYqsoTEZWFWAV5
cM12XWReyRYU3ecGT6tkMmy3JttUcZXPJjfLSkCYAlP0+LVu2teres+RrFjrh0SRgLmX7Q/7v4XP
mgE4o8EF7zK9OYjPwdwsOx9gCPfbFL29EzfxyTYNa+/HlHI9TPhItPxEEaY/Kvx5wM3zhqeiMQzy
0PfvK7/cyyy9CXh2z/I9qeDtisBoLieb/dz8eCm39FC0gSXYnPl33chvdHzNsbhSMSxYJWbMse9o
FPWncmth8tQGj7FPSToWmLm+ExAYN78Nmxm9hqy21CDT7/+RVGqXrGs5dRL7eVmWbiGUkj/lVlU/
DMMkWt1RwuzIC623bKQT3dFCg+l1AQUNAt0C7TMIeO5dL+GZqah8x87w/zPZGsOSok/BFWztVwwi
M0PCh0saR5SB2FPxrUU4m6CEG4bKhno58nk/In+gWYANOVNSG+QrWmXU4cnLfZZcBKyYAk3LlzPd
ZwXwuJVnnFhKJxH69roTmw67oa0jPf5/NDYmLVyLdiyJauVuPyMcCn7Yc37P24jtoZ8rQ8d38YSB
lW7xBo7ZQr0BeDx77ccgsjbCuVX2zd4RQ7RDVa9gpSWqJ2VZiA4lA8zr0/GgEV41HcSNQfttIG5f
A8Ts3qfGwr5Kl3D40k4fuqGYv/oKwaNVnxAElJNY4pPUp7JPI8zSS3M8GxoF3X5m8NWg3Rzpd/6G
UBLYO/jVVxqjuXJW4HJDNnoQOC1Tz3OuyAD7yONz62KpUZtyw+frUbkJAiGE3iift9oJ1/NQHhqe
B2v30M75QlJwDWOkB3iDQojwQiiCwZ8LZgXtC0b5bOmpmzRF+cZSc+geK/rbe0/b5EsuaW3BJWs5
sXYIS4j7m/PGh2GQqJYa4TIOkRt1TH7drN4vgg461q3UR0vpiFpoO4kTABarW6GSgOLvPHRGZz5w
NL/mzft6wjOKGy3CI2P4YeZ36uEWd+dwW5N5V3D7wKw+hcf3j+edMOerE9DK1dD2rwmBc/voP8tG
A+gwULftQknYztF4eYB12fxSbHj93Rwt3XNCeI+BySDD5HxCjFptabP+WlGbGk55vn8s5p3i2IJG
pU1bU+V9pAFLQfxL9ai5MNrfDwa0VK7fOwZ5GODZTJKKxiWJaiJsOHRKJ0i+eDRsxFUktQ38xbt3
nFh1/lGBJpOZNQ5bOYNMyINwxTfVQExI94LVGSXTwACKZdYreMQiYPvh0ibqA8ZELLdoLQyKwrpu
9MdFF1H8/mUKC4pjnMFwsxbMOfzLBi5QngpUUeKde76WJ/VBaR+gB9gzpTLuv9Bm2VLK/jHI8p5S
CqNqVwCrMG/H1EfkLUCBwm659gVxq4X0eIV4FyHNtxQwrNko+b0C3Lgt0el2mO2HizMl0zNCIU/z
mMoQrfBc6eTRmc1KHDQcl83iTCs1IxDzGUOWJS5FTfJpik3nflj+vZH8He+Myk+IupgPSLoJYHlt
DRsgdtC132me/Gy1Tr8hqXdJu9WPtCkv06qd8pFBMGtFt6NnWcc4Hwp3usYM3EPCrHlfHYRUp6Oi
WQ5RjV0+Gq4fCHoYwB164NWWDcqbK6EP0IaY8MxgrmIYA7ZVlet44OuX3wFHED9ykfegA5dzA/HH
89SE/DrJ1GaUWJOp/jmJNwSFlW+QCb3KgbCfFFR+fvSw/h8prtkRa94t6t6cz7f4QuTnICaVNYah
HlaCNEQt1VgixylRYPHHEVpfeYrbEQSCAl1KOd4sl/kR2J7ouKZpXKDxVZTAsDopkN7RpFOEsKnh
/72yLaxJYOF3p2t2yPCoHNFj+tI0cLea+S6K0G3dRtTLQGYDTqIZdC+1jT9Gq0N8ibIKTpPGgzxd
hWJ2TP6UtcGYAz7mIfufzoIFkiqiDk8B7bDRBP3m1FyYP1T4DPnmbHcHCBXslTgiTCGTlZXyjGsV
sGzcn76wMsWy5RgPAOgO5QBSGhdtXp1F3VGgJkoQRhNM1N0JQ9NnOedHtVyZjAnoSWg5ENkvkenW
+cShiOtxr6WfmrpEggxN9nVQQOgw+rbsNK+nym8ncpBfvQImY0W6D98do+9UAIkDLw8ZBnMCEShR
pdagsZgJjF0DTOlQOrHkyb+nyo36gM/SEtHNxdBapA5k+XmB4+xZgMerIzPRfkmU9B6RYAlgd6Wy
4+cDxnudBx+a1rKc4lHvRzP+t1hf6UYFHbB4A96yUe8E01iPhgYVnvMYIJHf+WylMTZeg/DGRPT+
mzGDoBP6jr45nFqhqSbbnJeohA4r3bm4cSLAq8toPQEQq2CvqEb9KDesRyWUYFrZ8GbXwy7WUh1U
vsz3Gn6N1j3rAMCBSVNhelkfAHmMCUADAdHrftCRP1KsquEsv2Z7/a1tBfOdpzl3203Al141awzM
ujZrPOdvUP7B7YA+q1XsGe4DPkWa9rFiJiGxLMMguvdrq5/uBE8Ll/yeexyiNkPHZWms+7OhOCl/
/tRhhpjIRTRXIn0pUHEDBeCBfbpuqICONRopcSD4fB+aCe3fjHwsD0qWqQXGnJTG6a8O2HBjerg6
xfUTQRbIbxkDHuDvpZzG/PisEPWbcrnnWHTUf4LXGSKG2h3jul7B6Cfp2oRve0hbxOB/kHIbvP0x
hQNyGug7j+gb3WWH7LgANpODCW8VuFIaxL7pAN5J0Q40czRulSYaSH5+ZFnEDgY0Upujw3Ou2ZiZ
uZlaL8QRRrBQKafMipOOuuEL/jQqqs8Hd6zwQIN7XvKZ18VuPjT913LBKgcnSkqQtC9uAw3xmRmv
KvmaZcRufmH9wpe88Dd0mJDcJqNzPKGx8PNrya4D83QTlw+KK+dd8H6IvUof50TLt5FDCbyzbHlc
AISXo2LBjfvpu7f1fJ3oKunNPCJi3vE3qFOb+Z8UWSGtb4/fGspG2lHsdaVYVYsOPifjh4LLEhRP
ahyKwpJFWouxsSmGc/UDbA3jmwy8yhQsPl8Zmbr5NsEuxVFkMOUC6nooXN0OS1QKFF5xoJnXulzo
AjxOesovVkepXZXAsOyrgZBZ5f4uVWVhXt90RlsOe4dVgAXWW5uWBCiqlHKww1Q/D1Klgi40Phpw
+r+lOeLXVkW/oBlQ0DNNToHRl/knuWT7ikOa/HtYS5UY3yFbQ+KagHObPMp/7kBQ42iHIpeEhqdk
2n+2Ky9g9YPICeZvT/hrUbdGmZwGs+xHpY6j2PJX9dzVOQW2zJpbQuz9LmoJQXIi8/8Oo4jyelOa
vEVIMAI4I5l8fHZhLz6N5E8vGE5Pur6Ucrk7XliCdSaisJlotBxO3q2mOY1n6siOxVWB1SowCnoz
eb9HCWppa7WCEG2IlhVVebPgL/EXHcudNiHR4owM9eNx6nSXnz4cXHsP5iJUYWPcbIfdJ9MpkZwF
HYGaCirPRbhRCMQgkvoMCJGNYb/Z0y+zctmuKaa1j91APat+Kf9GuCnrssE/LioU0k2u7voWcwbb
2TaLXrNhpf4jjXPNQjSX7AFpaVH12tdBgfpPI4OfGx3s1aTnEIInoWHFBoOOXn87C2eZ8Q3yLMTn
8OwYWhTxUed26EXUWVF2M2FB5Z2Zrvpop/uteKrywVjds2hrfLqdfKlSJHhj9R3tqOd3pyeHyX6Z
otI+0ESzBUYqGyjcmiVEq4UuJeR5dLW/9igsafJV2p3/0jM3P4xgVSwc4Qoeohv5FdFiJes9MCyL
tTkqx5Xl4xMaZNv3tFmSwnlfMbuzbXAbYYEHVRsFn10YTorYGoP4XBV8y2MlXjGUIrgjFRAElJ01
hD9onu9Z8PYtVCdTNYFkY3RGyPJ+EK1GkFqxzX6WcYZVJZrpF8ZBPHr/MSl+SsETCXdXhkmiG6O3
k/c7UzQexbPj2aFf14l7BX1J0n0GmS7r6/falfSh8eRhmCQyyMGoV8hCA4y92TydufXjkrw0nHLT
2VApfLLup7R2+4Z1CdpGFgDy/NZuLL9UMpA3jgnolPMKaPqCWM0nOgo7OpIaGGqTDfHa3+7kdbjc
QAds44M1G5BSeRZvV18exYp07ehh4jiNuGyoCvBKc6DnqKTKRjMD+MlxQABI6Vh3x/nrMyTaz3HL
phKWza+qYr63ViOgxmZ0oPDoacCNJCRtLKkHfiQB5prdpKxoVZh8mBpn+zi+/LXH88RkhSNcvwSR
Ih8lve9jIH3sWbyd5QSgR/QpyaXSsTbQv0qQJRWR5Ssk5jIrPDjxGy1i4mAyjZdfpZ/glNd4EjeU
274ja9SIj98dfYu14UJb2WN1P90fPdDKdswsy3b3PXTRNRyuTq7Z+gyGP5JEuBXohx+5UrhPD2lf
KFYDqjG17WzufnYszNTWxkQGu1T6Ws8mAqbNCboPdMkQ/sEud1Yg1bglyyogy25n5dBTsubmPt70
vKDamCnk0OzIviAzJ5OEBHsCS2f1SbTzgnPCkZgtriwyjoWC91BHdXHqiwrh1wpW6UwXZViR34mC
ITbpdBMNAyKfsmTGBgLwQEYFqBHvlXSom9dcvl5QF0vc0OhQNv6SG580e2OeHKPEbc8fJUEPGT27
YKiO8ZTXwqwJo8eCdh/LDGHGay92vlnFC1gdnfUbIp0IJ/MXZeNQK6y9FIPUniaZvr7+aWsgZzyM
k0G6Mp7ML9c8nKXJnzA7DCpwqlflXuXynYt/QIX3Nz8eb99z2h06hj7yR8TgjruoYu/bUANG4Jhv
vcX3tcnecZnq/sHViwLgM4P08rQiaktXWHKLZRR5KgN8SrSN8KYmRUrVLXrpa8oZGFv+4c0gkbVu
udqWUr9KKmrFQTdhBM6D+VZTWVvnswxkf+vNeQW+B4Z1RKU5yPyS5EZjCoFAbJr/1gt9wmaVWokm
6l3PmxuqZOvyySfIrrZX7W2d5jii+t+Z5ZM7T/lJsldzRDRmFhmL9Y9VAMLEhhzleCnRLAdo1T/e
0+N+i+mBlObUy+fpR3HvYdNoHbjIq74+aNVnLH4OlVjrQ7g+i4rUj1tc2frzfwYr/drqnzF4LsFt
/5Ovmv9PT3DYhZK0kf0Hgwt2uKZRYVjm+8ieDB4Rek6q9aqlYGnAEEi2/p+MflA81cb9sKuWI6RZ
7rrSAcgRC83dk0QNyCQAjS8VGrA0Oh0H/6J9wta4VCOWjqLhDfYslh4PLxwAuBVE9+2Wy/EpAsK0
oue5JBXS/rSlKeZ9M8+pxveRuwnnnu65jYgL3ca0QTh2Ltto2DSbZEgLLwjKot4vP5YudpUTxaUR
EvYOFTsi7Bnh2msPmh4Mrk1J5szjCWqxOJ09u3sJPjXj5hP74p3Q4x5Y/64ojr5o4Votregwp+a8
+CmUlKi+5QV/MB9s/EKqynfQPhPSR26/+Sz/fMGrKpXfCSB4rkgqicOYBwpbwL4v3UwjHFaCXJjF
jaJYUXUD2nrA9+qQgWcBJ1zS7ulK/dH8y+C+jv0ARasUE5z0XWPQja+ahYvleAbqB7/13fMToIGQ
fskupVeNkkr84tQ8DHLd0/glZV2TpSofnBCUyAmp8Ad71HzAVn4VzOZLbtsUtOHqVLCCMlwdqxuh
si8rzcM97b+CkvqCFcm+Y4KjCKR6Mavyg6BxUwDnZJ0fnlJ2/2mrJ46g2aTEPWDUSSEJ8ExeqULM
c3MxWPbuCTmwspeayCQb4StnR+l/Hk4N/SMAU1w3ajsudsOOiRAqZrrqiuXUVJyU31dS/BruwYx1
hfEdE9w7bw932o0ib8tEwv1BptW2nsx7g1ZyCV/IF7GOy4Kwa9r7BMKNRw40qlh/eY9flI6Lt8OR
07BMJU8AhCElPXFUHfX8pp/ZZiOXzlpVheVx5ln2XjB2xYnYX3TOMmz6HwoIdr7jpZkaie/YnhyZ
P3TSF9aFXTC/CYDE3Kcac8CQtqAycvaQu41z/kV9PS/2kPbYWR9a8xROYfP5g7FI28dH7CE9XVB5
DJSIoTHM4RZPBEQs1u/5uZB9IJOJ5A9B4q3FwRlhgbkLq9mXU7qIzRk4faKcH+sfGIJx2py5/8EJ
fv0NRrFAcTejCa2SfnBgD3mF+jok2VhaqUKqgO2RuIOzZEv2Ozg+DduU7dScGFUSSmx6upQSwkgT
FftXv84tUIh7DPFYs0JhN/TWrt0yvIuO6+bD/b739imIWsM5RPuvHw+6q8QL0rD2YbeTohPqBVhT
f8giOetRG/fTisUBawFsIAlfPLT3b2IR/xgpXkOSua233hsx2MFyp26fQTZvFa82ixraeUxPI06h
Ppl+2438SIvotYQowN25RhjtiCSMyQU7gGRJum+7xMZp/vxX6+gheQcp8eYije+ozcDWdKif74Ip
phY0VmS7pEYsPISwcCoUqcoNkTroj1yj4jcr13Gr+eByFD+PSBn7Pu3Qh62hRUojraNv5VnEw09a
hguXqggQBAOuDBg4JYzTO3CsgpOtVQOFuFAhfqHDDTODRpX42jRea1nzUXvRQDoAdtMUdiVN3qZB
GQs39Mpq8u+hMgC13FLXIwNxynGTais1d5Wn75Td/O7CiUGaEx7h0yfRIy0JKlHknNSFJ1m/qjEB
HC+5bgm34qMJkGlWbKHTwF0X1cpAuuFgkDvl/w0pD1E8Y9V9KEPUfJ/+nB4bkRL//1ogoXwsiAEE
B4jdOHGRZxZENX5gjh54hWIR5jhYlEomeSGSpCNKAPPRs6bzzTG+hORQ9gPsZ+OWrVix0sEZnY7C
houNvZ2pW2VqdUo16ucMeDiK1J+wN2W6vLD4cwxYhnEX5sy6EXek4TkbZRAnLEQDoKD728RiaWWD
45n8q4yF1YaQErRvwpAQthA0l25Gim3SGrhQbWhCFN4H7HUbDQCzzLjqQ9/RPicSzHLnnJcXufCt
57i1kvMlujHyMTbH/yDw/LHHrtCgc3sP2VuQVQSlAGVcE53BKXWQ31yYHfFMFSLyjNjqc7TxqU9o
Y5JqxIcrbifgQqopT/OaoBE5QTmHeqBqTko18g3t2KOWz4MbfIipyqNE1sztXlb5oLGSsxhXDQmN
DHBq+gx/+4WrYFdgPkPqABAe9LvqvcfhBFDP3vvO+o8Zq8NYdINjbY7VFWi5V1S1NVS9XA4GzEUn
jMmW8wUsOnGU/WC42TZLXkXmKsulCuX0W0XAAKt9BzWEwjjHKsyac09TypOenPfWbA3xpfrCG7Dd
wjMNo38oDEwxqg/LxSzq3kJ1z0oABxf2OEqOYqms/YdgOyfaxKy6QfOVWxZua4hHIAMHYuzG+snG
+ctetm6OEpYoB6zOs+c1IdoeRozMYQL7NUg8CaZW3ekSwKoz3ky+BjDz3qR/sL8aHYk1b4gskwQ/
Fjo0YygYahRM+/x5bvEHfAp8hn7Xhy4tJJ6yeLu7h9ooB2Ytm6DQeytI87DN4cezz6SnnVchknkA
ozz0/cIvBTrymQ77C71j5iSehc6sgi8mGI/ZtCXa577RpfAQtnSENUvZjY/ToEg/HGeiB/ofaNcm
dBsyaZSpn4zAQNzhDqPqBmAlqoiK7Ryp2cfXLUR827KVibmSlGdEZB+ZH7uRx6NIfKfVinPuKtBE
9OuJfSL7aVXHouZCiPIlHfYRDXtg6e+yc+saBidKh1MjCAvS0ea4EQ0zyBuGcv6WDDyHOr6SU+jB
ezvU1qxJoywkId8jdR91DFtiJI+0F5z72f6DRrpM+6V7kbCUU4GPY6iB1Oe/E8RRarzpBjLmc9MQ
c1K45aq/yvs+/P/GfqTx8R6QgAT3q3dSAZ72BKhG8J0MdEefftfaQvFscKlBFbdRUZ5gqKs+vX+f
ojOAajnvFhD5qLzcw19kjNK0T5Fj0ynjMSkYPg8fOh50s3dLEs6KYzl7qge02dnTuPxGVn+gbZD4
FL7RoChaQAncmLQvnUcNjmPZOqlDHtQVgW3DWE4tuFO3RusT0v7qz+LcaRuAl60QZRlvQyVLYUO6
apBxWfWng/5w2jn1lgjgCsxoMOrsrHMZAFix2Addse1AvJxYsDDJadLrClzTXcX/sfSpKS1TvKs2
kQw39utijivdPR7tlMtE75bZZq0uWzthVGXQxPwshHAT53S8Up+Rh3ltrTxUkufFWZJWidNtErQY
PTU23RvZq+JSX3ojGGeGBZsjHE+M/zWquk1P0zwq3ji6a3KT44av+STlwm570ImUPl9o2+gzVw4U
bNVvdUoSH1IkLvjQrrZQBS1YURhKgGOoHR1iac6YuKcQX46g6vYP3x++YjGDJCm+W+rSnHCC+TeE
dsZpJALxgMrOVYog89n4qJ7lYeDxwCxqjnfEfrZ5o2tf9hd94gmTY9b7OxZlxDwHj8f/ZOM8doda
zCiR/X/se4ak+wYpao9fUuQwuNsL/DNMMGZqwLfBbY1/BgBTeWRYHXDmp4stVzGXV8vgLHJL6u/j
aUmC45jKtt+DAcOnBHJxa6udkjhpHcuwTGtFyqiZmneT80TksVh7zwV3uqQIYXexJwu+h8dVNDA5
ErpznBo4JLdOIV43lqPoIpOq/jn+CtEe8Ey1RAPhLbcqZXiSiHP1HxCkOhkLraJqI9TdXANgrL2c
+izUNiBED4hmrKj8vI6tD4sdHsqNnu85vAnk4A+IY8akKBFOd7dFlNueR85uajfx/Mv4z8SR9Y5o
wiljerAGoISFh1mLenVMymPaUUHxYXVeEbI65AszvPkv+EzhTtGUUe23wm1PjsSaaaQsnHPfc/tB
v+IIY/vQi84BkinZvDE7+t64SPfWHczYCxVBca+Onuxy+shKUU7DyfsXCM9uVZ+uv6Rhkjjey+vE
zt35rqEMz2+0yVcrKrkCEFubd9uQb8NJ3TZZ7cxULyPABVAk/uIvUWSxRVSzTFemYhDeCoEFilTU
MfjphD+wUUhagbkravaM1Vfm7VySSe4dGr65sBy3OzeaahVVGju4l9ij+0lEuhexdDsqah4EzzI9
7kvy6INWTOqlafBP6hlnki8CtgwQrwi5Nwh+5AfAGJ/KePCO7LbQUNOcL/+DiyLoh6/jnkbcPWYm
sWZQ+PsnCitx4FgtEh45GK9EnK3RSL3g+sXuiU5hyd0J++gaTvanoLIzRYSYvk9OpnzBK2zlV88Z
Y6dRV/FmUg4soz/nLECW76bA5vGHNpHqDLwUY9LmQSwaFDSX2i6jJEn8vL4HKYWC+jwYSoKcyMPP
hcdViR8DiGty2vtFFdG5TAyH4wtnRfp7Ixj++rIRBl8TiVoWYZysDSoXJ4mwIt9SiZosdlHTXUDR
1fvtZK0m2rg1QvUHuP/SlHCjJOvDeKM/2vxQAcWwXahMjJty/bcprZv2ue11KeJoUnDfgskiOhV/
wpZ7Cbcj9bL9X73/fj79WfNyCR0GbFjoshDRKVUut08EguH67aSdIXXEHAiSpK4XY+r4FpIFZ6lK
CoH6CJ6BfoGTa4vkiYHLRmPiXRaDJpzbK88HDHSDAQTfCI/SUuQ2BFQVfc6hNBqRgUxodfACNwHf
PbICSIjB3rg8Tbmunj/pcYLu+ar2BJTLcfzAZcUTTiBuE5yryBtmOiX6/rT/ZtSt/4PCTTu9feDu
Dmw3Rve9BOjzcEAnhu7W5S7P5N0+I8f2PYrtxi+KLQGdwMSsjbmXcG/SiyKeKlXmFVZG26DCw0Op
vPQnSuum1Z9FsPbL2sWceqTraxAlXCJQePCM/Dsuu3WLrLiqtbz/5NGhQAPfOZsw5GhdovUSJKHD
wK1De+rXRAFsR0AU65XRtNxWxf60oxnfsuQnKBQg+mJ0onPt5mCmskwzKlOiE3QpIGdfaCZenBzM
s+cEWWiu6ouJrJ6xUSbxXNDH5DjYsTKche7mEDHHs34M1lFBandWQu3XyZWEWJmiHQikPSRH3SPc
ADYO78SJkZ2ttpn0XeAsmsiTN1w3LXaiVgLyWGIPR1Ra9mPY+LbTWCZHntFRhi53u/NVfaaM3nmr
x5P0UqYykbl8V6LSEYg9AX/6urTGKxmT4e8q8YDuUvmTtdcqvJzdsTJga1nGlW4XMgg3ErfiS3m1
L25gehQ1rXniXlitIy8Z/0D0G01tNq60vTGijZrpQxY5EWfjYD41gnSfmecaIP8Tn9Jdw2D1PG+2
3kOYTn0WGbHb2mu1mQ2ZiF8FKvNodNcb4SZ3DSSInsNSDDm01PEmekpVaadIAjQ0I45rqRTJUtOB
5eA0+/+P5GY1774pDZWeK5XKWhrA14tAjTrnVhnjpUVqpg89/iVFEaWlMQvWO4CCRiM0b/IvPaH+
hXG8ZSx+8kXzYiYIV1qG/KknxF1i6rpRn96kJS1Y5v6USQR1K1zK0XpKvUgBQZJ6vOY6yVFMf4aY
cPFiyYZ2aDW2wdDYaH6sBZ2ZfsJ4MFDWR8UXP1ZTed8xUcZ1iWYfiLGul41Dk7M6x9l7EaxxELjX
Eprfor9Q3y52H/qVJAWwhLOmvwgkM0Sfcs7tDApmkQobyeU9i35rH2dL6FC9DgN4uvkzOjNJmxsz
2ue9Dkbeazp/2wLq7Jv5FXw8lU0hyz13ti0UTdTPQ25eFAXMnPGyZyCsb+hiIRJbL+1h6EY2P93g
LKVdRxe8L3lMFrR1xJEc8ADVlJe/Nx/OnDQ/iHrzpnHWKD+kc3aOwNRpSAPgHMmyhEoHB/NjCOcW
182ZSzyWOeetQBVHjFwXKix7qTA9RAY0RgAqLKGaxEEUTQ1G9kz8n7gtJwD+u+g5V79KX9JqJ1rd
RCtyhOP1Et63I01zkgfmskjynWRLzsLBBQvYCjILaQ8X45BgWutLb2Vl+FYh9YqD+M5JGv+QcQrM
DOsxdO+UldzwAJ1DWC8NMYtmpjkrqQNV/3QEVxqFx2667XN0phdWNMcgJTVxoikzcCU1B3jSqluM
x3naRy5uRMqR8XO6CM6KiyUktKLL/AtP1MnOCEVbEkBPcmpLCZSL6UzvAQRJ6TAV8R2YkZpBmY3Z
aYfDUHGdKfLDfrauNOkuMymMnJXJgM4ak+MP4PWbBPoV7iELIatcaTckdWjnoM08q4LqzcaaX+p2
fTrvNuO1e1rxq6woIHVSjp5o9YxUXDHJkq6sQtZwWnokEuUozGru/ZKX7TZ6MDbpo+40vCqtUS/u
uH8X76v41bmvpyuQVzK2K69IWKaO5riefzWzjZmfSM1xmmcy8WiF6zDDu6u86Rk4BRUuTnK00pv9
VQK5OR3aIi1OaIPc1CzP0CyNHBK8iuq0BnB7hwvPTF2ZExqP6bLk50NLSrqRpGeIHsF6RWMOpJh3
5CPAwOcx3dm2YM+hypyASvPo0el4OEIh4oXdQ+88kS3WHXjvOyKXphRhelo36Oz9DckTiHPk1H9x
IOvEMizCBj734XSgs5Ex1DkaGxI2t3uxp22RXNKLB+I0yRym0DrsTXqgT0UjSTSjfgIWWDxVO+/s
e9INyFpzDBI1XGJf8VW6DF58m7zY16Tqf2QDoo1D890YMp6ECxG1nz57txLuL+cN3D1YpZQmMQiX
YUJaFoAzkohz5a/7LrNwG9mn5nXs4m5LA2wLehPyayGCl3L4g/wqTYmBW2wszrRyzLJSEgmdkGOP
sfos0a5mBH8Jg+s908iSgGCP5VuMju+QTVritKj6MmZJuakLjiraxWyubRuHlJn/gNKsf7aZ4rkR
teof3TpwvPE4TvpaoA1hghBHKIbKHcEu/lX1ayKGC6UGf6mvCi7ySRNuMPumIhLH/mLQSuD1dC/O
zd+/FmY8VlCeoLEpiZPC+UUsG552MAnZaOTlE4bsbnLEL03vcbz/9UyN4P+nWuk0mqL1Raey8/8h
XIwL1TYu6HPTPxBI75kxIKhtcST5ZYgVW5MPCnyYfAk5iY0w9+odt0bdOuSNajyMlsGASAgvVCZl
mzVWkHlHuIdr6tlLxMYNwhYHE+dKB0ycPEIrY4Z4I7bmqwnBMYlqwpa3HWD+RLpHQdDmjUrb0VNI
O3vjLM5NumKfgfKUVzybgnnOPg8tN91lnOvsolA7iQGjWKAW8Rr1iqre/Ertd/LjtUkoHAIyb1dp
/Ha7/YCDBUMlVEfoVfeDFX+Ai2vn1apDlKsNrloLpB+ozu15Sft+CDZ1ewW6Iu7yXAh5RseYIlYA
jqo2G17udzjdtkWZAGiSCbC5RTPWK0NGbpz56GPkcNfB0GlnzELjeVgokTqND9Fp10mcX55s3CGS
yvkhhE7zV/z07G9N//I74F9o2TbpgejGKTsHaTwTFXafObzJHmRs+P7I1iQ1rHAgmg545uYSntWe
loyP+U/Gpp3QRT5q8IaNljcbywZ9I1H5mrhE1gQGKfow5F2v2np1JJ1nbGywoJNKp79Onz7HX/xQ
mKMGvHV2IKc+gj43VordpOIubVKQd1bkoj0guY+cF+MYMnHxIc5ZimVOJgOoeq3fyVC9xd5njPrQ
zsGF/QyiDexHN0LgRFO0ra9BfIOvP2vZRBOw4QVw7PPXUrndy5D9kkpCHXaGHDj6Jju16DBo2de7
cxWrGqIv6zkzNI4m42BZwY2LEY/ZRbnUQp2L31hz70856ohQEjDztEQAbgQYARg2M/QrXbiSV1oO
HplrLfO89mx+gA3PgRaSGW0F3ZUyDp8giAnpuv5bnG9NCs9XGERVjHEkuOSVAbL7/iYmX2d55w4i
wFaJQcDODaHqlMTD+GlxTMCRaz+XPdmZrs4nr3hhpyZMxgOLNSUHfmkD3sbzWDNKVTBTOd2s81tu
/pI/NrpzaId/SMoSxuuT7AZVEJHnwdpOX/ycMEcyh+GsVxkpEf2IHc8uEwsfqhNIx7UMdzpUjjVK
vehKQHK/tB3JLfpo6lER3o+kZwUZDd/e9PmC3Lr47n53L6mL8/mqLiI2UX3SEDhb+Zf9dWspyaiT
1ObG+HZ/icVXru7Loa8UXdVHlXU0u9LydhiiqXA3W2UYg1jqdsE79u20AoGoHC7N9kcs+oGPxICj
GWQLNCySngbjcW8wlMKz6VwOLKyuOi95FSTBkQQoXe5IkqJmTyLNRtpf1QLIUkcIHl9Pb5uqFkBV
J3/tpbiXHCshKHgaMeGAj/Py7qstjQSSx3bR2o7+vqsnfAPGTWfo4K3h6Sen0OvoVh6Yo/R+uy83
I1Kj/0FP1xH1j1nDqgI0va4s+bpE5yKod7+HAsUxZ6DmYVzAXGzW7uIOdCnH0v4Q9J82k/SlIf76
gGXpCIoNhQEMM5RbQdIylUYNufLmRRMQUfnVAFMoORkCufhbZhILEye+WsEjwuJwGS8GFML+lBrT
r8GK8XIYjJd4tGu3NoEYnMdBucCXw4SK9ksalzYHKsCgtE+W2NGeWzfLdUqTSKVfmfFYJ0ZwQ8Th
ljSPc0SRiKXqbMndpocZf5TYY7OOBo2LaEPJffXKxScfxuRDUlftQ6bMsCuGuzvtDaD1fmGfIC5H
9S7pS11tuYcIesjpQx1TB6SuRqxwUj7KkJJz1gCu74n83Wk2QTJIy75Dsi/jN3j8gfUxJ4VVhL19
lqk+ADDpxO6epRpm4AuoihLlnSOtalV8lsBtSnmdTLt3vEwX6b21mFp2qg4kRYcyETiCIdeH9Z3H
bIr5U9mYst5oJwSo7j144LJOZB8KHYMpvdclRKcab+g6PC7v4Tc5CNcQDvboy0GgnWs6WMaPkYVv
bLxKPbtcqwaonOuzkCYtT3gzUabCm+o88npnP75lQ0ytMWrw3Lo7DjxuCU39J/R3BVAE5PYUs89O
zsleaITlirUXjmUkzPECn6JifUvTQIuOs472NxQA9E02lVNlCyEsxj2PlKQpfAdRPu+pqkIzduLv
dqJOQvQMrM9HaO9E72BRuk3Lq15mJYjs2BaixN9RJmqpRN04xQ7eDArUKMIwHKDembcCaST7wrZt
yjwT67yTf2Yvlyb4Lp+ntmfxQxF6C9U/qE5zCkRqXTTuDI4c8D+UV6MOrLxbu/kexTBbtvp+kBRB
QbHshJqzvBJaUoGdsg44FKrMdDqMaTro3SHd/xVqlTHDA4kwtoXD5AaQ7NALo55PTppzxCMXaYwQ
xvPQX25S3Q4AeSzTuFu1QY6GkJb/AUS3dMvdnmZFzI5gZHdzA3URs+TTHyWryKwR/YB9QT7z1ktw
9B1RN/X8kI42ffCAgHGW9wyeVPk3nIdXlUkF7fSgHbMjsUA+tZFkeRkdQj2wXJy1Jui5kSaFOLNG
JSoPYoTeYedUrRi/Rnp1n0c5+h54k9IZLXCTDCIZI1fjTdVfF2Gnqd1N8UyTd/vb+WhGHWjKwOrO
x9oCEIKGPpDMeCnE41G6cGb9kxr9hSYkyQdHvoP7RuzjB9lREoCAkb0a/fHOw7yHFMbs6udbngiQ
x/A1eRFshP0PQLUEB1v+CICXT7MFdfrer87h/KvqKAGu1VcrZrb23NFwrON3hzVWrKam0WARLP+f
JSMRQ+9hJe6SUVJoSIJuNQEqeMrOYMTH5YSczXOaXMuGrYbLdTQBeTkXZQk4a49dXrr2LZxn8QEO
KhzF/AI6ptvLsJz7Ys4YXpKfbuf4n4FQhT5KfraSfh42lZNq1mlnMyqk+rC4yMCHQ7qwsnBNaXLK
0SUWgzkd3Z0wkjNFP0QHVs49B609x1WZ9oIx6IlXfNbTKagjt4+EG6/nhSVN406CgRRWoKoeGgcY
eDTsqW/0GRAudeydxj48nY5jpep/H1P6HnRa7fnHCLLKMl0h+3hl2jZhmlG34IcBDYWdcti9Uiwf
aOoOoTZUNvH0e36cE88oe3MzvT1zGvz7UCNJnhJlcClye5EgNBc28zgfB416u0mrelOHkRYkU2+M
+mfh7F82+Kua6Q7Y0LzVglcjVxp+rW3/LFqBqHLkfXLBoj/PczLof55atkTp6ts/i+YUAzV8gzXb
E9uKcXj/UvQvZX/JyfEPCLu9XhwcyLvYcluNe8VyezZolmmDdGTqJO/bXp3zI+yS7FSAxkNAChLT
tENoUGAdlM+cE/WEHdOmJVNj+x2qPDRf7dPSfjgHL+ZJ1hWuTLLDPAnW90HZ8QAb68jkdcvNgHOJ
vBl/BakUWcnKBuGkeRHr2XmIrLqAmnLsgc7n8Xx4tLYMWp/8mHY2gVK1HaoKsP19gnytvQviZA1w
s3Mle/xGHGpsKUuPbI2PEz742lO9iVaF6LqTav6xHjwD7un5it/2ZFUYdtkMC5SfUDlmK4K/y1ZS
j+Mm43TOWu2fPTHuEE+Onkz9auI8xiEYW4ppXTpLCZ9qJ2dmIxpYDzTcktGoqZB8LjTMSDLPCj76
CMBrI7n/0S97UoBRAA9awjRJAtEdcCI6nnzOTbWBWSVAB3ogBYC9sitnCYwNwaJmdrYq3NO9BprO
iwNKJeMaMH1D1wd4JaD2E+RZMK+wVz/AeB2ynAL+FaQp0oDtPt4p2YxJT0oyfjzGngwqSwV5tznu
m1hv+mVDYHUEqjpspUZ2+J4ahU3y7RjadJFeDUQhBZpPyDfGw7uspSSQlxJVlgi+ZAZlu3qm6ZGG
G4DkWzYdYChs8x48gUAMprO+uxGGQcRxLrEt1TJ0sk6a5fwveEz4cKulthiEteQAG+GXGLHWUDT2
eaf4BCduQVsQjRqUQDy6lMc4v64w3UnfkX1aP8GVCaCY0rrVAJui9jCEMnUM7XE/fzE3004e39Wd
eGySeS6BvAhPINp+RIq3hQbkQaB/Vb/AlsJkEYVFjz4IOA37ex7qSJ6tKewEnWs2VBBEeGVsPxk6
z4xiM8Kp0SBJm3h966+ZFSUZPY3YCLe1baZqo2elGqmzPDt282zopqDfVICKKWssDw1SWKk7eVWZ
872wSgnKxxt8Kh9E3YiLaZBsO4FAtkXD8v3JEu49ara0qcaffumoYiEbMJqJBQtLgwrkQLxP2a04
ey42icWDmBTmrqctpaFrO81VTO/rTr3tDufJpbG10fBVapoRcHzJcbjRez1Y0MYLESNlsVJINVti
KiNAzefqa12z0qgmYpmiKsZaicCM2hEUnMF7CzHc541yBpAczxda49NV9moDAhiPrmpPmBcUBe+R
HECzn7eVwNZIhVQfbMmaOjCFkw176sdS0dR67oBGSP/vVSiSF8xkdT09BsHiNw6Gnu4VYSAvdHTP
po6FYe3YrAnea/HDyOQjboOxGez1p7dqEjz+3FURtsz9wqdN/9yiXMQuatOewQEdFJjsYS4jdXvD
gNGnVs2UICJwlBd8hul2g3oM7EcgVP+pgDm/ArJOhBYp5bXD1ZJcrZbniSeY3tRn94rMSb2122bR
/VifGi5naG3DTQQN63bigG4c3vngRcLKoABTE3xqVuiJS/zE4bYv7SAoivUaoFrEqGV00CgK9P5c
aaRH92z67RchhoXzBTT77jL4e+vrEMCSIsmLRgZrgL8AuJX6+DFBFE3VTFB7AF7sBbxb5eQVd+wC
y8QGkmtPltZFIRuKVtNbKDohVbr4pw2b+ERXVY51CU7tZJcH36VmaYmV7ODX0GWgCgTNXQRQMoNg
uY3+zNhSOwmluKPrdU2D3PtMT8RFn5LHqlt4gT8fUdo8DhcDzb+c7wbHAyiuVp/M4V6TGkYkVxJl
xkVyyrR7TGpGHULbK4RxIcYhWaCY2ai7UUcXvwrJD+EY26SNtR5hvKKqReSETTdNP8Td9f2bw9rU
KnLQtJ+reMknsjkzzDWaNd+6Vq2b1pizpX37Z5rerrLBCnvBdPxYIDUd0MtZoxbH6RGcwj+CdZWk
BxlUFN+k6XScEhdv7GkP30JJp2PctMRk8CNn7XmIT45rSM3qZbZOL7WyrvqetzXDxrm1Vqt0ijVK
P4l25fC2UVr0Nc7JVJ0JPuoPky9ERFcSJqxF1rjb0ROzfMAAP5Y0bPES4GRA/ayA1s8hV7PGRPt7
b7oFPuQTBqtFh5WvFV1oh8NOLfv1NPywERgywFwqUQSup1JwSb0tj2pZzYebFAcBZ216zYwMrd51
WhLFnij7WABdgqeZSW0bb7iFo2d+hI2Q1ntZR33X/dvBd9bpM5/XvHUOFDVlSVgi6IJ1/By0h7Zl
YBxrlZ8z9V/NgU70KqSxrp7FhqSt07kOhsuwPp/iO1NGLNoJP8FnTHa+LjvQWKAxRPJsgSrLMb36
Ww2Fk+IBhB0cFU6AGrw9PN/WLE0vAwHvbyrpfxocEQa4HtkikdxQJr5/qlOk4vihV42u+Yuyq6pf
GFO7y7k7QqN94D3m3PgjcXRO/Obbg1zX0zEioqK5/6sIqW6Eg/i5Xlo3Gj0G76BkbQLKGbPtlRJ7
yMhndjrAgtcdDJQ8tJ1+wevGlZUovnDNpLnx09gspch/xUQpurj5zudN9wUo7ba22Kl1oI3hZc3c
WYoPJBz4ovqL63MaD/9afePt4XwQuLqH1KZmuuWX5lJg0iQUnutxrR+NU7CbDmhb5K/3zp4eiet1
qKny+YUJWgWsIHIR/YIhPuX/RAf9PYbXCh1huVmkB0y12/XTpk3GYzXLBnmfXuAuuZ3KvwqFMdUq
Qx4gb7hg/8ZTGrd8umRRNXpz2JojQi+k7n7FG+hgc5lsjCWnwAPHe9Kcs9e0BuS1+USTMFlNwzgE
wNEJIywL8LMg3ooU27rBfaRP6jdtvcQZBl7QblNqPuFtD1cHDajAcLNMdRYAOjV5THQU+Mjxz1fx
pSC5JrCIjVOICVZxKPfrgFFl+XalxRJDMLXKZTYjt26K23lTbA3qZOlb+TGrTkl214Kis140fSY2
pVQ6JBf1mdimoWelxVkn49IhRbl2LOYQ1ouXhIz74sMpiu/z6d5oTtfibwF/9RplMw43hdnvUl0u
0ZTyMk6Fy240UkdFKESoGlZYxrg4nNRyIeNPhRN7Csj00uRb1Ly/0aQeccee/gLhxcOMhfPJUE3H
yMfVBIX1TgEGE+qDYz2S1lUmDC9E8OZxpsYvMpaweTrjZKxOT7ZDkKr7bXXeSK5DUgQnGdyqJQHN
c1cDcIkfrcwUdAd4WdNp1z0mldqOUU5wfQBfpjz8UMBthihe5nv0prDs6ZpaWzNjYb3iSwkz1DvH
fe+O0ChIZn3dPe+zr/PqtYBPaTuUo2MeH+w8J3S2sxdjpPRHMp52EBe/vkQH+/MnjPNVAeuoHqhH
0hjaNlTKeLs/tLM5lZUekP6voI9I1GV+nAAFCG+TCutEuNPn7LDHjbwoVjhkpiStYptRnA/6DNT4
WrBRc8yNf0gMRPRpHjYWe/O0C9BhZamSd9aPDedHVv1LnWEp8EJR/TMymD/tv0ATVifrzUk+kYI5
ondD+GeQrwRBMT7XC/SLA4+yUy6ok6RXzhskS96WI0Gf8zG470BALN9cnuGM2jjuPZupMs/MVpAz
QO15sR6mxYoj3zNzL7jYzfk0ruoaCxW6AZSuQr9g9kK5vB4601yzPQEoO2PsMPmwmCzr9wCtC9WC
WaDdg1sgUvNPwgjentg3sxivKUtwIA+DtSPoCykmHaKeCT3dnqFfW46WISFF/6fmxnud4vHecfm+
8v8Bg8QiVnL+2EbjYtdY2ksN0sMzeFcsPv2Y1EtTAXroTuQMBUvQ5bDbZt8gwDuRKL+1KwelMlI8
7cXkwlZMcKX/lSC/WXxRqmEQvTD12YrYKDPUGA9FrLJQlUEiPweMpMupKzBZLBII91/0IKvVGyKC
hWI0xqX0C20rhbyk3EVHeNKUGBh2rvpPqaBIafsU5lcagE/RSmP3+8XY7sFqKQLD2AjU1S+Y8wgJ
FgtC+n9CPaRPBQ9AM8GdKKxXwk6Z7++/M+Mc1WLcuj0n8d+0i/c6rGUNScY5TSsUSBQv1xpkL2Cy
6RXYvQG7ExzxXAAQ58oz/5L9SCsUA4GGvLyNCq+vtkY6kD1fc1JiHFFBgJvmjH0yUrv0cOZVuGoE
RzHPlGLWZMQ5lFza0YE+2cnTMHMz68XvFi3tdkq4HPjkIYclgKiS4x0T7HlHfXtRm7NQdFF/QR6j
uZ0NUeVuq7cBp4ydb48nD3JnqLWoSWi9/LZg8vJImvj8STC49n8T7jAH8VuiCrWS5v5BI80GzqO2
iu99HCzH57DN47fK+ffmTJJG43Z5/7C9xMeERkqfy+NOzDfv3dnmn5l1A82cooaE0aynrSqkRYpV
6QWgb4OZuqla7uuaTByIuUrPFgJ3GuHU8vkWmEQkCwemO8W0TcimeW9JHGTNchEqmq1deGYBJvAq
abIfZ+cSCtmiIgovdusJTkdV0P7nMhQj4d5ckUuxnUESCMkQuaMS5jcorV19m1U99JJ/Ho/WL07n
fFLfCoYDdA32n9dWZg49sPprLw8Qye3wOhW5elCKc8yWowqlINg+aXmjfQhx7ERx4fzIDzGf4+H/
kpZSJnt8lbrN+Qc68S7WUAFVsF0dZoHbYlXisE6jZQjLzI5LGRGSyXgfQW/1R22Bdcvhdl12zFGP
SLXxTdk9l1ro+q2jJqvo/yQeGxlE3q/uIQx4JcleMTkeSX6bcUsbOiI1737oS8daVifBrHrt7OpB
JTmdG+owpt2pR47Og7EysQVwgc7nOS1vzaTUW5+kMmn0IfBA27UKwtSUY363MBHrEAeHSdwteqI+
p6vmRVEoI7zlXRxs5DR8quRVDtRaG63RVPwTH70mp3wZ77JrlHHJhUbGMrFw9ghoLRbFmHlpcJko
TYVhtyReb01dFHEwyTYL+rjlNnRFPA0SxSjKdnLIlGzjeE9RJofBJT9zX4tyJj5LimU5V1GGqf+0
bi04c+uS7JTj8/njYcjnXnciltM2n9OxkwfWV6TaXyiDODtvz7LV1b/fEFbUtsGLjdkePqRRQmsO
a9+muge/EnXTQvfIcUos7zyV6WpwqcTxyfHDK+aiV/kfvSHIEdzR8rpvRzoDvt4dkFl2pFCBqlj9
0GdnWeb+E1DiWfbhxGWR+p7e0A73yh7Io/2QGF+gJDjuzsd/rn4jOx+MHL6yTm/rnIAx+3NLh1/2
VNUg2VzQ4gVRhIXDSqh/zKXSsaBOtqiLz6wg8Em6vLC10kAngCBs9gOr6xnhJHzZI2UJcH92+C0l
pBD1s11llg44peb02peB69QcA9ANtSsST6ONGjsMj2dKrEIhn+DJQHWdRm1vjkWZLp8lj+X2yIMV
sux4Y05lymvpcEWF8aD0iqlU8n+vADUT4F6jtwV/CG59ZKsHyLMYIN8KBxWqQix0wGWj89gi/OEl
b9/ticKKWn/zCOehp6YUW+y4PduAPI3jYft/NWf2JNp+Nj/DmMMtu6zMB2/wWSNlKmKj0nXlNuFD
yQSWVu8ecCi2M6KE8IIKrS1yftceFM7+5h9j1kjVZsRD0/NEzE80QRt38l5aMlRu2v0UAN0NDp/R
IIgFkkGu2RwFXII1g8Y6h5MUJTEPis3iqi7H2KtawZ1ZRx9ZHy/AjQ6pQKDMroCbkXnOs6MkT0na
y+sPPgxy4FvAk7SgJxWJ/6q1GJ+sbhdg9IYFbabhIdMOc2W0DjACB0MC2rpsqqng5ZzVPcU84fxL
do0BOZKaT4hIqQRcdyD38C7wQZMg0jrVMScY2jndUZ4P6o82F0tPmzLeIsyr1SFgE1gZL4LY8pbn
iMoutVyo1wfwCxCaQJbn2eW3z1jelGUiqItfXbi/Dd9dMQv9M7P/MDEo62Q0efNFVfPsDnKpFDRH
6i/dRJGwTh5PrApykpf6uInHDTBGsrEjjuJ/GEZBsYux8BBvVQIbAIWf6X5EH/JZR94oYqUC+y2e
jJXNHYhhElzLw93oGzOIyHmeDIdJC2FSnNleeB+48cOfcod+2HybsIStW2rv/19YxIe93v6njQFr
I4aK2kLsocFWW6PXgJ4wVG9e7lzfJ2BGg17nnf0+PFmvRe8JQn0TxIP2bQuA30O45RuMAMvB/Mro
Bgop/nJgWAxUM5C1fqDQ4WlSN/8kPcqHYN7KvcwEXoG+RKmXW9cIepEDgwldp5ZJHG+9LWGN1EWV
mtUKdJ6a6+19yszJikbOL9Y4bukgKFtrrtuw/QOOW00fandfh7EOGzvas72kX9BcrLy/t2rYNQ/Z
L2uGEjUMc6PoLK9BgNefoboV06CCSmWWsmOxmNh3krSnD7Ju1zWW34gvjxa8pIyTzeeK2+Wl0Nkb
81FsoTlMFxGwBZEJbfmzHdEeCQQ2a0tvJu9BJZb1gzzDCS50+k4BH95aBHDGe4KFPj4FMWZ4Wkkm
FrVuEyahMoPDtR2VVCnOmqYVzExypP8M6svsRy9stbZQZIEGcaN3p9rzZ0pL/duPblaMa1dfPZIs
ukmZUBUEeC0TyB9cqEPwDGJyJcz2OMpXdeQmCbA4SHkaXHuZWY2UyDGqF1NvxL6kNzPe1+4s6ugl
BgsQYu381rPK89S9wxW0Epu5zidX0pLvN8lmKE4DaCtJwLzMG7dsfgPIPsWU3npNMsljmjBty8IR
GkeFT8pfINj6JFY+5Hk7r0NIVYiHrkNSnrEntkm9tn44Sb3tkWr7ym7ll1POCB84Vkch6orw/UgN
MXJ0hNGkMYTAq1JoBnZiuYwvnV6xSo39X1WYI/GWQCV7Tt+KlXgGPKeYM/GwnJZT5OneWe6sg4So
cK4Mb+m8GaTWEn83/02kmPQ7wsY4QaTZbkZEEgDT7LtYo4FPCdelviKwpk1llkmhZ1hl2CE5eZfc
yoW/I+uiqX84FIh94KErBYcwyW4xl9dvuuz2DXkRuH91jONqcekD6x3taXNjrbMqAagf5cocU+a+
hLvyQK/keJztIvxexjEH0NWaOUyjl/0u2YM33kw9pebzBpI5sc2Z54fv2AylfeTztMhIpz2Bli78
HJNl3Pl/zVknZeBU6kf+3l+e+eV88kKT21Jy4LTQeKWXjbObp97Mg1CJehJ4jk9GIWXziY3PfE1O
MECIt9PMH5vWbtjzrQpphnCk2A0EPSU8ZrB6MVI4B5l+C3YAHfhP5Fh0K8p6eUKfm1aU3GlsyEm7
zktCpFONAClHQvwEi7dZ59a5RlONZtx4csmaOLfKoENmzSxLamKl5uv7R+vfvt/gjfQ7DX4EGqKh
paK1G3NBldKPrjApgw2I580QmfDwvK8Ttmgvh+lepOVM2kFfgPK7fbIQTVu80XwbG1EdlJmAMqjy
9kCw3qxKM1mEaSWyD9F57Qnb/j+0xcy0tAlQPujU4hKmajt6LxJEyN+k6KF8+X7nw1RiPa5rCa/2
Z3LchWjlPFyDBqHjagRoKgl0nkmdARMCBD8afqKXN5PGkGlEV7GLmfx+35qvomZxOHTdKKpI5lqB
Qambdkg7mZxJbwHHDUc2S9bYIcDxZKF/Q+wNCxRrE+HtR8nmaCsrLpwcTFKluZNgHIrOE4khl8r7
y0yiPjblzGk7kWZur6Tpifzn81ANoUBQEOavq+vB32wFDMPvXiAr3kJflfat+mabJ2hTCsSiwcxo
OJRI8lft8BLOsov4LR068n+Tcew4dAF5qWmbjlTJ5gJ0b7AmBD6XMmYDwPGaLOXPOf+pWRy5myoy
snsNGTQkBRRhiemT03OXc8Drc9wHuc0gQB8+hZKhwiU4Cj4BNUrsMQFZMu2dJV99Dcd94ohKYTel
K8ScMq/HjSbqij8urLXrya+FrpX7aMVmrErNATCuqCwU5cSyhS68wB3Nw7KV2dnyRhfZHQ2ch6Qf
Idn+yHh4hJ92dd8omP7o1UHsjtjquxI94dySUqd/GSPvNIOG/vs/f9vszvMdxUnMsZt7AM6c7xE7
CNqkhvb3GD1zeUDiFzfe0ydJh9gk72hiNd4H9qw9ENsAWNlZvkSubXc3ZWx8dXuG08quyklkV6j7
5My9GoUHTXH6Rv5VBolYmGenoZgQaxFb7SXw43GlC+s+tJMfRFM6EC9f8t2hE5zP7xpKGY1JaEZg
JNEenTVDtC7sJErDFXZDayBRvOxo5Rec5qoo3sAbpcHL5xbHC6IdgDJ7aUPGoO/+CjghxkXUQxRO
KlJF5qBECtCPnlbsGjXoKjRyOaRzpi0BshBAHefjWflAEXOJ9WpM4qKt2Ju9bLl6xBqq41UifwrG
37AhgcxxI53ucwnNdDCrYJGOuGgkcWmiIjS+77yyhxAx0LJ9/zXaw0F24tQ3vDFBwPPaTtkyYbsX
u5dcizqWJJ3/f/ncGNsSFlfz1fcCUxwCEHXA33UWi9r70pcjijI764XbGVGkRwerxTpW2XNGiNFv
fM6t0OvNuB31szl3FeTVZlqwIkDku6ZJkeB94KLYpqq3D9x6jzOvPFYJs99G2D6JhI2hxkRoD/6O
Br0SDfYX2K6gb8iIC7YbIduBAo33pq3XykeYWduVBLH/CVyOuRZKy7RYmXeopy3zzSuMnLOtzatO
IoXbFlmoAFxXvOpx/EcaiVoUm7lBPEtaguIuKyDzp+g1HBYLCBudSkJlB9SrXTwgqisjEkH5SB0P
wMMav5+tsiKx37TkimSUPZ11IwAl+QUg7tat30JLE8M/J4c7T8i56Z6WhIGT7oTEuL6LkkkuA6MF
zC96oP1rvhshkDaquBBI8COd9iLZjntx0FeA4fhrsSRnFLLHYhCfjoHYwhDaa9VoyL9d46o89tEx
nKRD2JDB4FvJwGzKPkJ+h8XYhn7eAC4LKnnNnaDzlFQ0As8pKkNv5BZx90Uv+Yz/tDo6e8tkpRZu
AtcBw9zLhT6Bo2qDUROxqqQXwEBSLFOC0vuOssurp3RvoYMuE8qN3OC7qQzl+b4jIRTBQFY9QA95
mt6b5IzCou+UdwvAcYnhTIaGCFxPB3eV+Io9Mdsf9SLtAH9MEbZ+Y+m5E8YNQpIWIDefeY9tJheF
h1aUkxoUEovw1ssziuXePL9yfd/S4vP0UGVeAQPKH8q0TsH1hQnToG9/JIEFRaxkt9iAoBBPKbBK
LgZTpQtKqy+Y6mDWeZiN1RYzWX9wPTfC6d2KBC8NVLySi3s3GncGso7rQLazsoSqXBKOrqDG7Y53
RBFmMZFGk46X3JuqMkrIGGvOK/E9GnjXo7lyxUeJOeR7YaVEoSattVQdHyGsmjTQlfKjoRDH8IHC
v+OMOncCBhNw8hdygj8+ogX0n0u9BlpX57u9bIukzK2hElnkP+PD3Pk+hTDChSo6BQ9Wx4y6wD82
wJviXLi8ddJ1UWio/3qdZrIdJ0DgLguzWaahVT48CujBOf87fWajaS4aMfc6mtWdpJWP1ggD4khU
Hr+v1LziLjk+c7kZlNyxbpjBWiwDHzEGsrDIPkoxW8o5+PR4ybXdKU0AN3eMDUawCXzlrVjDfsXZ
u/BHd1LK0P9lwg009j0Qs8uj62+sBj7Awe8JNgfsMP8AcledQdC16sMePbjhBN+a9i89Nbeb4yRa
7c0JY4oQQhXLSmM2r4TnOIa9DYWyWkLOH1Y23JQurOE3GOJVdrwJM1Mw1ThESnugwpZm6QbDcZ7K
0RU00N73EybnKHCxrvGhjD4HP9Q+oiTBwFD7Y5o4XHtKFc/+5BBM1+MQUnq2Q2AJFUNPmv+xn4tr
qx9a6M9rOvCwc2FsaOgIaFZF2x09/1z6kdMjahZdiD26pfiTsLkcnHHXOoEpF/yMkkYz7vej8wPT
HkWeM2kIS2QDXKSiiMT2K+DDwK8mvCz65C8UxjiOPOjGeS935dCOlXmignCyi8O4VDqxFpsaYhY4
uWEyKMAuWgg4K6p2rDIgxk8VaQxEMyY5iGx2Eq8/ymIcV+qu5V2mMTYX21q5HpuqlawCBKBBqsou
8kemnJ3X89SstomxZU+SQSS0vAKv2RZpJr8wyX0f9+ZPffFTBKI7PcFJ6wD0tZm96bAuRlXbbHGl
WuHM9wveGwsFw1HUUy9Z/pydJ+00dVKs6x8oiwRE2R8vC9vqjlvHYfY/ESSNNrVjzpN4kbxsXSh4
1oCYO9BZ8lJVEQ1OfprcfIP/j+zgETIinz3Dt7iWJg5NVk5U/3uSbPlx2gFhZ8O2IIyl8LcUYZ/X
/OJQdqHsYN2rT5gobUb8JY2/DIisSLevTZRml9ZUcG9hOxKPzeuXv2IOGW0zJzxZBVKklEaV4U9V
C1gQZ0io8lZHobEhyYV80Mq6MKlStRKrZVtY7X4POYpFDNEcNj4kDAaKo+Pua+7mxub4b/q4jJXP
F1JfO3Q0BOBf4NBzu/YVk06/AC6bhI2hKcLX4vOSfszdAqazaEElul7raSwuH76YWJ7s71zn4Ckx
8Tdm0dayNnrm406d7Z6BdzZjsiEoEPu1ZPEzAWljEchz/rlhy6fktntPWdNkeTLbYk235yTjftJg
uReNsBLxda4sTHfhoTN9olX6ZIqZfeePUHhVC+hC3LDOpvDG1pH6orO/mb3eT5EO5xw5rXBwQYc6
maFmftoFLhfjTR517UCs4MfYqI4+X73+Xu03mI64wTYO1/9SXKC2y17HmGtHduKymN/h9ZSn+8OU
wIDSdCremWre28tyPaLTf17oS1X1EIyOuC13iWrxL9A6UxOUHKmLmHv01fiOxCLiJOEfjOrjzlSK
ajIPhFCT0PRrXBbrBedK9jwhfDeX6cQTI6LJDlx6lxIH3srv5YoO0XWGPREe08ibj/E9T+2gVmts
J05kS96sDPFoh6gE10I8RtG7/jEr129qJhGL8M51VHkuddPnLUgbSqEzE7GHQYn0S4FrJdtttafB
3XmJuv7UyvTLEmXMHLcs2sDAVwRLvmBk/oCqakJrvIT0aoBz7jeRgCpZCW2FAntRP/exzNxhGjA4
fzjdA+S2vid5tQT/Rj9LJBRS6PKpmkRfPX7Sl6Hur6d7It4vxHmaPwNHLllmz1eXFFWwOm1pF86X
boEoukMFaTv8MaQLa9FVCRrk3MqhbPgk1Jic99FM9sAj73F51wfFJmWXpoNxqsYQuj/yPMxiFlVK
xytBYAXQdnLPuknQfep++2Bh5yN9wEKmT8p7mdc9275WieTUDNyOIBbaTn/8bJrpr7IkbIYuQS+g
AZmYec3+pRrJWreUeCXSWdnN5LtA5CRL6uglzQ5GgnYdJb2INFv6Iyk8DF9ZZRl4RMKeiQ2meWqt
p+6eXD0RaDYUnnkUxnbUD+UBR4eAZkdpeFsvovzcqSnyEpWGFYVeNFdeRL3nubJd/TtxPrKWGBqX
BeMsmYy7S1TY0UH66ULPqCNyTrKE/6zLkDUaY8ckJX3Lf1ArrKTNCWO+jm5IQHn1hpL67aowEw8c
UN+c5tel3FjoMmTnRyQRS6s7sGhQPPnM+/9DMe0/5xvyjd2aaFh2G9SD/F2lagpkYnnCZ3T+d+0Z
ubBdtl1sk8PBmxF3ZTFlABkzpmdzQWkDWoN1Cs+gyCz2O06p1fTKekpn3bYikngrl5dyoGTimb4W
UOSWkcBmC4nlp1nJVDqjvD3xPnrtKcHkMP5Y9fKDFnudAn+d178EccONguSXOYkQ5Jk4+sm8M51V
vN5YjYJ4aQ2MBIC84CQMqnxQTMnTgGeUY5gHMuqV4T4QPRUtWciC/tZdX9bnkIlb1ZxptJXq9lhG
QeoAjvhkj1AJ2Ofk+KKkJT9cGO6cPSvrV4CTMhi9xnSH9Ha8jIpa3Q1PRGEIj7yxGdGAUNyVbizb
1UyqtOUEq/0vJKgYBbDlWnvgZ7Mo4gS2E9lkOZCXS71jC7YD1hzQ+bp+W0gm7kHH/b6UQMrLUpBX
MiTuGDb8DbKoGrjOaJb/qkJqrN5Kk/kybgJb9I6uSoQcxa/okuC42BZS+t70y6zR+rcTacmXnF5I
lPs/jn5wUKjwzf/Jqmx7895mxhSCjsG0rHrggiCGIohQB7YAufvK1yXcnQmeHD8SHHIK86eydrAL
P8rTp3A1ErzD1vHcIB89BbU6pphcMf1qFBWnsKW6sZZOxwFCIxiZywswIU9ggxV7Vt8uX8aF0QvQ
FmzLxgmfSYdNspptYfATPFOyaE7nD810hQ+mC5RdhZpZRs8C8dpncerQwMeRnZxUWCKHR1lXU2Ah
Fvdgkp4aMM+zoT1mAbckkz7gizDP4JVt/JyJHT4QjgMCw0R8kFymxqoAsk8ziBMXxJnKVnrS1ZkV
OI1nR9YWNzlBuoigM/Xqv3MQPgGJm0pUQ5NhX2ZmcaTrdBwPDvNKnqKUgGu6rqipBZK9PcpfmnBY
WqlaYCDVSXhw/Ltl+2KdKCKTpreLcIS9ZN6a/HKgt1fTKBDCFHuEGS/+jwOcich6z4ZElVd4SfX1
TNAaOY2FoYQAFSGlf8qQmeUKMCVoqHGeXsSLWLEczm3IoBoYdcKyTTN751ndHrHc8g9+XNqWBd/D
cgE82RCPDRMgPAgI6KRDCr3FcHX90w9t0nzdy27+RSa8IYtezmiD4oPZT1T2EnNMCTsaHtyvadq8
ji/V3A6s3Ppu0gTSSvXvxWNb0ssoIDKKsgtUN+SyR+HQ63CQtnBmaXycamKXtjhGEPRxKEvoLBQA
LyJAUrneIXw9asQpvKVAF9LK8457x9V4HajZ0yLQ0cYgMSnfr0P5FI4uyoQkRCFPfpAn/ilwtZ+J
kQ0aCqA/RGphIuRA2XJym5AMqq5QAQgzahEkhYjIr1hsovj85/rvuRg6NKbUpbZaakvXkodWCT3x
AY4xF3O7m5vfz2rqZFfC+SCiFl9oIBEKSH3jh3G5cAAOt1/uA7atJ5mdlmN7MG+kFfF/ovRZQwDl
URWJgwqRR4m6k9fXsd4iel08iJ/whH+WU970bxQiC5BH3IEB6HrF4dSbbqmHsDOl8qISZQapmRAi
Ye0kzNadFO0FzmW/TJL3s+kxJnbY9WfO5MAB8Lay4pq6SDbnAu1qMRTeLyWBd5M2aYqPc2gQQ5Vz
/cIp+P5T+7rrs8tlb1azdNle8njvIA2KHX5HMkP8gq+Grl5uANJuDCZPgbaXg3cNQWN9gdqv8o2L
m6rGYGR5JFPkLiiHLx/VtLiqN9C/P2GFX9wYv41ZByWDw165q2K9Rz4dXQV/GHFG1/KNqRWiBclj
5XONSQBsWv9jYEynj8bvLqigHVdnYoO3Tu3UJxzCNjAnKg7ExN7G/Yt0Bx1WNxUx/HHjMLH8wdRt
ztEmrInjENiGfQ6wJj0wmMl9S/v93EzSht92iX2/vQqcBYQQ+sR/qQXSKKdc42dKzFT4WcWnre6A
eP84FME5ZH1vO2IrSyjQdK1JynoGZJO9ZZVb+g+HeNNsCOSfq9X42+k+Q+5mGGi3baa8wnaWrFlj
Hu/EnjczAHUeNaabMvxCHVW9stJYgmhAWdmqyYfRVZcMMpN3haOq8sktNLsInNSSdqwS2mOhckPz
VJvnnfOEk9NkvjC+lXSEtbUy+MQcRN9YGhCaIDIFimKLGhjpQt4Jyb/BxEKVfYHX//yR1fb+htIg
gaLyp3/c53VSuis6chgp+Cg6GbX1ud7QZqMhV2QEgdpFjbAQHnXN5czyK2QdKogpfHaRa1uQjnCN
VXnWLVgp/0S/Q4CM/BjEtDvtYpumiYbyn/mFLaGvC45qlTdj2LUxhu57EJMPrjpiakCnQKc/F2br
ffuJAuBjcjbA84QwJIhREC+kTh0HN1JB7PlVAOOIk2F3i8YytvydsF9iZ4BDmmgB7J42t3+oEg52
GQpZx+G3kKZ8hZH8utpXplIm6DQDKZlQL82AZwoFHMQpX8TARSf2YtESMk5uYuHsI4wbQAp2hxwd
V9sDXmGvp0GZBjtlz+0k0R+avgr1oPOS6qqA4SbRtAiG/J9JKjGJ6kA4eg8+gbuH4ykKjdn311ol
CNXicujTqE7Xr8mYT3ov1pWs4zvekMDQ7ezfNRaoNskTkAj2W5JttbBs+SjsSczrWUq5kxrRaEY7
iKq2LDBgYq44IFYEzvpFE2vjATIzbtJF/LoCUDrt8qydZjdnf8MpXjdFvLVV89DOioUgQMF0udF5
kI0pJ3964zGSclmKzasYzVMKJPTqNxJfRdn3ubQfUk7wp0JZbcc78xURfVD1TA4OEUL2B6aNQ/35
RwRu55Tflgf2TcYYp4cyvTWQAqReLlcoH38k0aTohk7NFNdTCNdFTLKqdOPkXR3vc+CMab5fht+S
VQ0T6WXAJVfnBPvsqeGf26fhlMkvCvw8PfQ0dyzXSONyHRwwORX4/PiqhxHvkMwjV3rqCBMLa3nZ
bXgFZmKzcvhH5IR6Sy/3xJpbSSe6oKKRjlnR4Y2S5nrCSgWzO87xElu9OmW5X0YMRf6hiNWGrLYn
Ew7HKIcHLxfj5OGkVkKWtBQrX0bPqK9RjACSipp2aTF8sk13BNfJtxszTVj20PcV+AioOjzn3lZn
MTrNtRmvqPM1CB7oFej3sMIeGihh0NK/ShN/dBncsUv12dnbxyTxBVugtgkVhSzvicogLWwhBKjZ
CDIRInbYkFhFmic49FNcqDeYdXsbbkhOwa9PFI48tYGAmoyCbcRmXDAEeqmcWrAVGiTxvXYn38Gv
I+NxpKdW436lzOMQCGBIeTizEC/DXCdaT3NGQLPq2TxVlPKPTK4jUaIoHjVRVpkswNUX7Di1atXN
StExi4YxUwBDdjyrduMVpeeI6uVf9lQQclUuVeTyZ60t1c7V55mPS0Bsaypl140DRTr0eYd2Lg+A
2FmdpN99C5eIx8pS88/V1Qv5IWZXFnOwsv/29pty4TUXozqWQF1NcXYpeaRPduo4t5t5fIZ+CqGv
b1UuBbajkyCzCr//LiSVh/ipPZUMLlAmmI6z1kwY9mIj/FkaAcUhAdq2XJ1IjgI7MBaYvTIrBAZ4
X8cgqF2jvTLUDobtS43q/GX80jppMshqJleYb7AvMeQi1ODe5vUcfCx6p+Sg5ifS5fH07MOUecAg
sMvmxYsP6uoZ1n7hdIdT5ErON5nUugtOk0OwMxu2jMt30rLVcbvIfsenQDpzDjgRHwkEl6kxkehK
+F5ZmWnfuKinxGtFKd3PraidqqugD/WSuvuXQsRLSYpbfSygoNemyyY9EQOtFa6Q4p723CiTtRy8
PSfHusMCWUSp8TWkuzIQlYi6+/fTkFcv0IUlqu3QDOWdoZbjhX/xmLfq7BbOd7JcKDGI2ChV2a5W
8RFDhbJeGPlE1vqG/Zu9Za0ILbnjPAY+vTD5FU/MCxW6Adk8PZAPlihxW1a9uX7pnyrUQrKbvX68
YYTdSFFmwizKRPGZCso04IhpztgmCQIQ3qD4EoFwR20axV8OpJAOOA3t/32VEZC+pQMGwczlYOR0
qkgLtgKOO1t6Wy9MshQ7ZZLrIJfz5KQCXdLSqbvPy/HyhudJNVAzMJm8wE04EXRk5rpqymB+r0py
eEa2eHDaK6DjvtvhuqlYMR2efp+zx3vVgCto9ZChOGFZrppTX0ZRAXAwTwDPr6JwOijdFfOEMIlX
v45gw7rtUUBb3ffDPths+JvQ64+tYgUQ3e1By/EjfuRdXTbbvNwSxcuRu9xKlcXqjv/oEb8m25oA
JZBiR6JmEelhi627yFwUqQ1/P3zXHBXeqlInEWS6ftpYtxAxvFkY/YJr4wwvFv4zf0Wttl+2cKWd
XzQoH/On0Ot6HYMTuVwO0jLUqxCGGtXrgLVVfti6O00ni1iZh8EvBkzflyzSjMGETNaNqDOaDt/Q
sP42RBQHeUxxPZy22HUli+GVnxK38VT1xMwp3KnaN8KsHq6/oZzbCGUH5ZbiWsUhQyntinWW9G5o
gJ++bXCOMmBU8ek5OCwQDd+bDeD5egeu3AwBzTGbyfUJIh945G8dusho7XVXKLSioESl8i/E3bjt
patTvNK/iEi1Kw7VIE/ojkI8S4Uk6WHP+rzyQKP+ZPHjczlZDGKiqj5cbhro29lLlbSsd7jL7jBZ
r4u7rrf5CyEBFkc5yX/MS2mCRGlVL7r6V9ryCgyFokRxLzG7xVeu5Jucf7M/xHs1b01nV3MnBWRl
gfbuRKsT33zrFlFn+viuqr6P8FRKkD9Qpj6sdQUskWf4pcH+bL/OG/kkcjBZG3Y1GQmStr7bP+XN
e4ZrZgUPQyW7pqn1L1odiYIGaMfs/RlJeKcJu+4Fqr3+D+q3hXlL2Iy6PAKUxE8Ua2R9V2XVEqS+
YuUG3VABXR5iXt0yMqiZGhY73oDOUtQE3A5huP2rnFKPdC9IXEbYEeDwkVr9ZGZ1e3MsM2KxA8r+
yUnp9SigO08USvUSHNAyp8QU/qoaWGALcv1Kipp7pk6KMnUvgYNXy313p47zkAYM9lepB2jNuYpi
1w0GlZe4fCRBWc/N1BcsHR7/jQnOCqP8KQMudVsDaKwcVebZzhdzghhe7CAsw7C5qqfNqsso3FFg
Ju8g8vgJjWx0KjJBAlMQFbtSVZuAzeNsKttyqtMN1RrhA1aqgKa56+4qu8ho5IirqpnDlpuHhgEJ
yTNjkUqLzNvCmia9+MwYwxIJAGPYWQhyc24wHL9HnUqM9fzhqy01AH8mcRbFpBBjGwin26pPzWoa
CWHQr91r12YW8npEVTz8mdgJRm801W7afMNftdWzJ465vAHN3aDC1L8E26lYLl2K0xBAhJZGShCc
wKgRMC3g9lmAwVYMwtxg/CioMCWlLPLPIwqsb1DlQ3iKTp29FwVoKWR17OtUmaBEoQFXbTG4r3sp
e956f5/IHwHymQ2WJRyruAtO+tNnFoZ4dovDSu8vV93ql4UxIpw+jmBI6TlYF1Xh3RP6EoSxHnsn
rK+yb5QB3cHjnzf+H9Ba4EOPnDkEN5UcRxTqoaQ8NrY/fiMTe7CymLQxxe1qm8NJ4+1L95Ho1Sd2
1a2TdPp1X1MT1l7lOOSK+MWojZI9O4QAJJOMxGcfroe4v9TfAed1jACBzy2/a3SNgqwDzw15eSl3
YYl75CPRlnwM572XDHiXIguBdmjA5KBxUOX6F3/UMa7tCBVm8zN9I9tBe5aY1GhaKgHh6cnCyq0L
jEh+opXa2RupGdU9cpRq7Ncbt5LD1sYRP2DnhH3STo0kJ/Sog6OGrFgGbjAxildOwaEFGsG63vLz
FuAOukp7tMfDe2+wmN0set4cgA/0SA906aaGTzaIVGWJLtpHNoT0tWoJedz9kLJz14sOE65wXQd2
WSFZpvRdreM4xp1MAPGP8UaBk4vNYMM5cGBhtJZ+uJbsJ1cuoXnR66yd7PPpwElXHUX9zo1fc8BU
/FrpMvKGVCI064RXKMz28TTzyvDEMsj4aHojenZsjPnPnhgmhsVpY2YsA8FmicQBKLCbb8nI67li
WObv+6Ca2NV73bxSLezB4qUy3fhebAf/yTsmBn2RVhVdNtGPTUXf7+HIuKYHO48ISuDxHu6Za6Jy
tqC2BSmqdpIzJZo/cCwIaWO34pbH08yH9gDsZofJCg1CRm3UlaoI/mTUY06qylW0SFLWaD5qMtLx
Z0AoB6Tvy2YppEq7dA72KAbMs/sLyeXMRzBpBbW8MgWJ1RFCExn6wM3QHE/es37sNI6Xuy1OQ0oY
teIegzNuIV3nj4Aa/ZXFcj5dKQoYwYAxd+iS98QOlo4t2Q5OXAFWzR7u3703Ic4fxDs29IeADv15
C5oeEp7Fc0lAfHdSk0z2o5ccLsgb7dGgMuiVafY0bZ/uXAdmXDHz402TKH9p3yiYxnCnq6V5fRvb
Ri4oWGCQS52n/s6Lk2JwkdRoUkM9+b1n3LU6wpjGDC4Z4h56JnSppnE9NluKWDGxwH7xXJDOVyFG
vrTesXlLwKSblAtReAOgOGkN6uNa7l9R0ONX5iTjOsEiLK9SjZRVB2OZJkEbgFnKM0uVSnFVWazY
IXN3W+7HtimSYqVFE8mAXq2/r2djpS6zPaqbf5Q2d5yNBsluXk9NNIjVaiFcL/Au2wASOFJ6uHTJ
b+mmqNegGw3R5YyWwttZL9fO3ag1cdWvgOzXrVZCZ7ht0JAywNJCXkPWr6f7vlN2DfliehQ+lYEn
SklTY1itrlLbfmfVWPeDnHIf0MFBipvVOvq3HQ8cPx+eRit42nhyG/qdUkam8yUXs38zThCOO1/S
sgayE3UD2JFctlTb00LB/s0ZE9Ru4hKBvgyr00EvkpiidsxzBjtbrIhsDuw0IXABcEWKcbUQaBTT
z7btfc1t9Kl4lXqqh8I9Ce9c3XpHB/LyYglEDBQUHneXPs4p+XFhRr18DFar6ztJjhZWDGG7HS5x
lRATYbn/jsddpstSkoQe18SelXjIg6wj3hLhFauKBQ5BSeBaRJ9F7oaCffepZhJpvlCRYlUgMO3C
zYROx/rx5GWTJf32m6Tg18F8w4thuV/FuXGEfjYWsHLVFSBag5YHF/Em0/HgXKuc37EbbaHVxUPc
Z2Ozv04EJ+4BUazdLeKO3oTBEjM3fqSmMX9WoefbGV/NMf4dW0QfQ0c2ndQsVfINxlySQPQ2SGxB
+UEziPbuKEneLVJ44K9YQE5sITqqm8sKmY+UnJpoLcX0nihLxG2XJ4wxUnSy92QVOpHxtQEK0yRu
WfNcvbFOXjF5N2AqUS2dgUEv26CQYkvF+FDmPGHz0EY2Vw76LUmvsu8gtWVAz6nNq2QxAl7t1Jh/
mKvjDK8qxYQy1SxVWnD/NtvttCAVoFDTxNTPkZUv/yrkqUVfxFPxkrluwuBw1YMsWnTMo3CuNdTR
HwrEFBxY7if63JrLezAKc3xqVzqTkXZq30b1zJCorrqp/B3bwOTaqqCdiLIEgG7kB5Q/WVcEO8UO
JTeGL+NGMFuLz7KiFuDBJVls7RnLiDbvHK7/eLr8QFrXBNw6QCKaiN9QKDbJEfWZbV1Ncbn+/Zjj
5IrynqKmkA33ld8QZGE4/2mk99PNBaHzfLqCHZp4i3gI3zIpVLFbuRQtr8Qv1qYFhii6Z+VmI4F+
232fUCpfKJkq1IgXp5X1ngPSnJKNmwdlmqCgbQzpeHa2VtjNozxdomiCOlNnLSIdU+19Hpiwpfcr
CmK6JSpUwr/ekPe872yDe/3IpbWSNmUbKTqLYzIOA/rSDwHvhtoJqWsRoXciVe64uHwNJQimAsit
h4m/oDWZF+Cdpomq6mAwMfxLCRxdrxOvFTkp5S1y3vrHbKoRy9EIdmd/nWITtXMNWk4WOAA9H56J
2cTc/+6aa/MhNoNUVnQC4FOmIwHrS5/yfcxiuqA0RVEArfR5HuwAcalgDxmcQJhKUlM2II0dJiW5
LbyTsCKX8iUoeKt4F7vN0XA63chprmhEq8TQnUyTsdc3AosfetNM2F/9y+yw050yP0NjFmYbdSgV
gZTa4Ae58UapERQXxWG9KPw4UA3PXKRn8P/6Q8qOX5qgjX52guCn0rHhYALezi5v5z9rgH41fGLJ
n2qEGLnxRoGRBu9hH9AvzqMbE9EYx/lQUMS3qX6gFS85sD7NufT1lfZnnutdYT344UkdF52uv4En
TO+0HVhkPhbt6qlSEs/AI2xUuFweYTiEZKMeBxNINEQGVaWMZJSMwQpMUsZ20Px07FUnCpDwGBzM
kzt+J/YQIOCe8khzl2zJ0YwtWnwg7mswXs+Vb3xDubpR4Nq2X9u2aTQeHQUnX7lWbbTk7pMdbHyi
2P7klkk9yiwzpok1SVs7EnK07mFGt0ho1dE5R2gMorWSrGbEHlgDgLmLY1gdn4VJSnv20pRCTKEh
+zZ2mII89fQ7mBqXR/EFJbKxdGwTx9EJmLyTOSxWMvrL2MaHv2NJlaBShQbGtVjd0FM3HCdMB2th
T6czEacijFD4IodI6Bj3fx4vjHemTzmmQDCIJ2tMjPXd05Erl2qIyUMHaEdhOXFyXtf6Mg4wFb7h
TR60mi6w7DcY0JDfwxfZhCJ/KyU/7TkoiJoG83qIZfAKm/qA/elnxGB0r/1oyDgiQTfz4LYwNnet
gCdsfRjkqrNjSm+q68HUkqKql/kiN/QaKYjryDjgBLeIcy9X7ULPhYssHHUhFfofALG65zp+U4vL
YT1vGTcyPHhGJZpRA3r/jlUhN4DtYOyecPfZbzTKjAvodlw4UiYJEc9miHFSKZRnyVz7HtikKvZv
5opx3X9n1E9ft94b0LkRab6oANUF6fZRpqZjNmRoFED+wFDNgEQMHbU9gBqfPaYIvS+O7otfhA7T
Pvh1uAUs87gJSU9Tz15JH6ThEyHleOfLsU7elkpPW5AdvgKUXzb12hRAAc9NnYcexqITxD0Oxo64
JlViJ7ytU4sOeqYn/hOTXj6guGCYr2Ctsy3jRPieZIcNZjr1Y8uwvGJNK7yI93jL8NmiUwG1YNik
havQSzz4dVh9Bw2CW+M0lpwfYiEhhepDlWAG+56+dpKOj7MvXR16UzKNIP8+WMsGg5Yd4KssgACx
5+QHmTCGueUm1R8IRujWpYc1xfrFeH8QnnQIQl7lp6NboncMmwfWNg5VbixhwTzDkui1zhp+/WsD
pl6l7WPB9gUU6Dd3dmkNZwERaYU8Ag/qqL5pL0T9vQv5nicjG4+nXwfhDEMp4I1V40sczP2mviyd
QzV7QQn61KR/4Z4SmdfEXZDSXlyByFAEDaoBT+9e39i8A5Nsq/kcjCYhXg/BOPOU2V95lpX1buDB
2tmvfXSwzwIU4oNE+wCbCzWnAJojeVGcWFGUzt42RGCB49Bp9ZD/EDBmduH4staPeXGF0/Wfc83M
Xma/nKD5yJFujoExIuF01pIgvn8Jbj6PSaHASDmPWGS/DpsHAUN3/IIrSbpAdX3yCRHSowgfSMt2
7onRJsJy1TMARDfXqnxWILVO2uQNEz7ErrD5oCSagV02kOUlHsDaCR7aBtbAySaeRTFCxUVImySf
WxdFet5IkEPhr3incujbjZiBKUVut/2M7CjKbDXX4QSm1fNTFXyGtrez1MWyvzV8LBwQFbLtbWe8
aZO8r9yRQCA0hDXIoVGA7Vy9/NCB4EqRFOaEhXbYULgRe7TFPT76RL9l/MXcsFibJrg7RYXgrLUE
iYMKmktX0oMw1ailFJRoOSRGB+1NG+T4QMJbPGyLUbaGAmtVDXzONKQ/VCO4Ps5k7HAH9rmLMxzU
/DFHULuTjoMHsyfkW3CyXqzEFIgd+1nT5OTUXa6CzsdPB74W7203lW3+i6An/Dkq0ERWLerFp9g/
TRPN7KgyXqTp8v+XDzA4FI0FagaMA27y81rs3hPJ8fX6SNtnrA0race73umQjkbPsJn8nUNJeMYk
VEXGRD3L8w37/AAZ4+1JrSNGgPeMZpWzO5/+WoHAv3Zfqt0CyOqWph5B7+le2wkxtOk7eIRSIW4Z
Sx/DCaTRvG1ZZ4R68eFuRBdaO+2IdL2GceVLjyBl1XDbL1A2jfUqSqCEbckC+BAGmWz9Mj87srtM
YCJOiazcS+enBaO2iy3emgpVNvkTX+WRliaBJLQ6wmNkcwiQ8OvUdu4r6e0fdD0bMDyxwd8bJgzX
C2blgymfYu4c5aeU8y2iQJ//Uwaxbr6CB1Lk+ogCM5uQj6dWoedAYqtxIkq5AMoG0cCj8SuioRz/
134E9ATFnRE7IeRr5ijEIkvij94hWxCwemQztByC0n1d6AjaaKaL2G3LzcnwugdatVvxtpk2lNWM
cHNPw+TQ5wc8pdnfaiKPJnaCpUNJrfqLtntxrWWV+cHCx+yEr/+YfwVKyJJi+uGzj0Mg2B6h+Qls
iAIdnjEy4Dn20R1YBr9SnsTjwHLIPu8Jp1ed8GlLxxH3fhLPEloN0B9XECyt+sAogISCtGrdE6d+
Jio02a8L8h8zhsEB+EQ8PYXBdBf9EBau30NnxDPcG+JGGWjFE6gH+i0E2lUuFo31xnSPqo0P648B
XKidnkS/RRGjNU4Q8B9TTBpDDyVhXjgz/hEEKzDuS7EeMjH7s4nPh5tta5fSRr0i4HjKtcGg26+G
iJTd5vIup1ZVX+OS1CU+whvk414TCylinmqypNKDpCF0HvfPfDSULZ+naARmojQB8Xyaf/Alffw/
G1QoDwBchFwwGTJrKiGE6dgL0WGQjdyHbse3GMMrdn2ytLmQulxE473/Dtg0Tk66gy3+HYL5snrl
Zv5CP/n9lEI5q1JsgVJCLMuuvvE7vLcOLu8Ov10/xEIBS77Fzs9Ib8+lFHwfiz+0Fdp/9sN+ZVYN
DtSQ3H5XK/Nd6j8SCMwc5QsOJ9o6PFH3J3Y7xGGsgDQCZO4Y3PouYozYWiUEdrrY4an53RgWSnpd
luN5PV5ALiQI9jRvTAsN2/G443uRfRoJXMbWmgvM6ihPkLZ6KzJKSDJbXBheQjr3B74G+x1ljeS4
4vBjoM/nure5ZgSHBPqdwlq7TRfFX8yCJqKYl9MYyfxjuDWHeBRfpparxjKGV5+UpmethpRBqMeS
QPIwOzgibAj1SHJGDIM4pd/Gtw3FcZ+FkMlzTm2Aaq/ZXbOGjZY6orJWK2N9VpRNSb/juN9s/ngS
78YT2EqEN+PcLqFOKfEPMVEZSxicHSFcJeAdcZWjI/RKJEek0Y+eJjJhO+/uEW523H4BkWiaGpvl
MIgsBz0E0CwsyC9veI7aBAyEjepMjA3bfPmA3acutgBW+uZTYspXHCM8O/nTSf38JuSmh6GUBnw/
Bq0oAkJ8DTmQPWMxH60NaFNuOR/1UqOUsz8wJBbl5wJ59tCgMpkbsVnw2FYD1ebDqHkl7ZP5cKua
+oeTMFeSo77qN/pzay3nsqZ4hmkv2EwlCZBRHMuqy6QUxEC5gc7jn9Wao0huHG/XB8LnBtpTj6GY
NnKRuTtBE1dtaEiYJGuNe0PWFP7NDQ7W0Zb8euYw0Db58UIaDeRu4193cPhF+gps7RkxN1MNijJH
/w/xGrT3HGup5KigQeg0qWBB6BuGqev+urkHz/wXs9AXVGGQY5WBAJOaJrDJiasQ7/j/FcR3FBkZ
/ww/sMXdGJ8tBnmcnCOtF6XY0z4MKV6UZUuU5dxipKQQZABDXwusUJPFNeanYCTw5hgmSUmM8/eB
IqrEYZ6M2+S5mqFAz5G8pl6O606aRk1LPLSZGBly8rOedCfle2NoIWebTxvbkjBDhkEoU5P9WHxL
P1P6Dco/Pb0RcFUsQHjc7ABHRE67X2iLjrxHErwE3Y1+r4d/r2KX+ueI5dV1+ULEZygoRClJS7Jw
ZsLQaivovqNkfQCiisqBUU38KLm/lZ+dUmWVUoms/x129Bu4D03gdlZimqAQvUDcu779PbgYEDR+
Cz0ZgDEO2a3GvEUUf4GRv6n9S7KStGxw+zUdXaG2G+Yg6J+YPRoKllayqBQze3jRN5Sd4wmCf1G6
Hd4peEfm3deS1nP4L9lGi9kecdcZbKrT0Is1vt0Ol0pCQXZ67vgWouEtvDQUsOhk9y5Eg4Vk7too
Dy+YNtWiMRVWlmnxpQyvphun63/RMha9vDvFLVEQwF7rML5ogzgU+bY0Dbb76biEiSDeeEabGcL1
OEhLaMAYaOzC9aMOt+vFasluJjH80CrmGFvNKHXiQJerF2Z0XW0JJG9rqWKR99mLHcDIOGC6EbEO
XksWiGLFgeiO1Jlhr2YuzZnnQttdP3cn+po2DsP29ZsrR9algKQ62SsdwSl1b4bv6gWkZpr49EGf
oZ0lhcJuDmc5Pw1xPQV1Td5TmeM9GWc6AwWTpe3mFNVLCdxJHzrChgonrmZDZj08UE6OLCTv7zGU
t7yLvhjaTMlf8wxINUp+6yFS2m2hoKIj/zab0MfUzzf817g64zZ8ln4YbW00/h70YRNRhIv0ndVe
FwyM2FiAsV6FyO0KJehgxOabPsF7F4lkkUq8TKK+kJI0rrrJH6BFQO4zsZ2mn7tMpaGcaP8o0TUb
ALkXy2o+LruwFOkw+dI7LVVAIiNA2IVxayZuPHqg3uYce0Q4FSRuo3WjYqE7KrcZZHAC4Rd1Fnnv
BpeoHYlDH2O1bgk5pc3WLFKo40MTOD9p865y14rCw3t0gH2JnxvexmFeBYI1a1HDv8vtuIOnle9b
KQuA9Tz4rQGRFZeVJ4PbuWYoNZC7TH10gvoKM3H8JKYLpnmY9Y58kM6L25BnpVk1xXvvAyelbphw
Thc8uvrtLGcIGiS5ONuGTBEkj42wiFvLqrDoVnmHKnPtIvW98U+CUrfFaEt6JjhwlUHmzBUI6DdC
mQaothXH0hdmjiIW3Yrt8Xm1pTy79un0Z7HQryZLA+bctO4CRXZiDud4rzZ31RosjdAELh6ioiQO
wDVJPE4kqzsh4kwAu/saLnb1Kp9yvwBr25glSTlE10y8J6klJSc+9g+ygsrbk2u/WB9MH0klSD/6
O+WsnWYblFDhvRKOxnmfsc2JJgVuFJgjNq/Trrl+CaSuYX9mj+cDPo2DZuZvrGj2IGX3DfEjXJCO
00PSbap0D+SgsyGw2NFMHt2CYaIzAY7b14+czqTEBkXOMuu3SGU4e8TnTzmE1hFfXr0ih9KPj32b
7F/jfrWmeNtj26v7vucfjTI7vLr1IETI2I3ymYCx0e9bzFTkDRFnvDUj605RJ6WS36Zt4G85Y7IW
4RVwP1FzkAc91sEne5cXYhldKsg6L7KldBYjPc16/1ii0dzFpvh5cJNkLISFXJMmauqOGYTKiBqP
xH0n5EbbyuU1ckbmNFNqKjB4RHl6y8qeaFKy1Te+EdHJGFJ438ljC16xkYeOOBgxbmr3vjjFHbaV
2Kv9eQ+KZKgeqquH9hbyww/VPgZ3mPNITrBPzes8nYVllM25l0QtTgm+CKK/9REJteUsIR7YGvX8
L+TS5LFYxHqQemVS5XVuNShfyseDNk6vOZQdNS5MWmrvywUyWEQoIsn+Jy9ecYZLDvKWBN2UasyV
smbL4zZoCgKFnF5/MCYeBDET/g3XGZmDbKLDNxfXy/trGcdxQH0eJ1AkcJ0SZ4ww4G4dV9RKsHbd
+Xi1RwDwdDK+2UQpfVXhfWXW/f+FYKw8MVpPH+duJfP2ZU4JzYPOTCuRfmwHiUmLnlLY6XKWp0dD
3wJbAMw3qu+V02Hd/p93BIOA1MyrciZEjUb0jZZaFOCtkxwQ9hRZ5bdyB7v9fr5WSrDTtbIHxCvf
en6pdyKDlKNAIg9go/A5T+b5I8ArngU3VAbaT1mZHI3v5S4A5cJwiCc7R+lHiw2ZnxO5QnE7Qw3Q
LaHS7AfR5aYkkXf6kpsCox6q8yKffRi17Oh/vHqsxN+mIf5JsOTtf5jESSD46jcm2TW1NsicaCQd
3grxDSIA96eXawbnBZweOOI1WnA8sKcfasiQUbGaqmfpUGbUOAMbbC88xF38cGBWN1rb9SFOTCOR
F+U4QvFVrl0HYwEYNgTkcHQGiQTY21AlizcuGrE11uNhSR7c2oD9/tDBp7uDg4g2IJltnpuq4ZCp
dveXh5kmJcL8Dwl92k/Lvw4ZG6fULtrr0cGJ+qf8EFG72mtySY4GALy2Ew5904psWAapPT7vixXX
LLbC8Upy5Mc1lgsKikIFfbdaxv6aj4p6eza3VtkYVA8H2SG3bueFakcyTsIAio70YGa/0rjUVMY5
1Tu64VfBLmJ1o8AEg7vuzsqK1aSEjSItYZ8ww5RVIicGSkP9yUsHMiG321qlVmDguuGTFk2t6NkU
SoUdeoe1SlTgtmnLcs2NRzWoqki6ROnEZ66C6cNPJ/5kA71rSjwlhb3N5I4sxWxHe2S3BOSNXl86
yLY5beMlt6aE1NNbGd635V5PT6DrOdpgEJ1s2FHA9v/cr9CDfa3qTNWu+ehgzexnjOSLWFFWuXRa
beOXmN2shynecxC89drLka4GUkBRtaBnRf7A1hpOZNIplydeo+lL8m0rO2p6oLA5z1bfv24X5+hc
fdrB33QzL3RWiDt7cl7H6RRtVuyYC8IypMSpYJHpShL7b97CIQzZ3A+SuyX98zRwxKMzCcg5MADM
ncArqkWa//XNP8CJpq3elwXPlY0epPeqsMI289uVH52P4DbtXP4Yc0yVQ1nzfXrl4cw+EXhlWuhU
hKc9+sbhHSkgQpsok9jKGEMSXFu1ghHHrFeHsf0SxiByFWkvBr5mbo5mt/dDpd/i/deXCoX7H5ox
i/t+3ekTxs+FSZeIHZ5tfC0nKDZl50R6Ow6Bge+ZMFXEfzq1oVutCF42Oeg8GYwNzfn4JzyaSdmY
Ppm5WIwGBMcSxCN6Kl3j+xCmLEGuHDlYdZlOuYnMSx6bOLCU1GFcGerBxC8rbg4DvEzOKqZzf+Hj
N4NRI0CwOpjgxQ9X0iWRr8diy0AjCFS5ZTLfDoRerf9Gs+0C9k87+YH9o6MPqOfOxhfIrUJI9MpN
X3bXTj4RaFSh4hryRUQsteIhNtY+ObJlfMCgrbiVKrPEnpMa8oq815JJAwpD3qAye/J475Rcvrrc
dJ+BRPVrOc/208lytF2KOSXa1DgC/9QqNkDV8qzZtFqEdRKUqqdIdxMFWpaKsSwXLXPZKleTzRym
suzXrZpF+TxCNrL8fGzJCaD2GYARLLpfuGXVqvl6TPzVX05KJo+QHMXdGZRszL6DuJkTBuxjTidQ
RMlZyIv3WNYpyG2xQo1XU7MScr3mbzIzjWEc8uqPtFVur36g4/S/kjQ4el1BLAfdc6U03s1queoU
81epkxpmNaMfVlmrVJsqH4D6+oyekPGHtV8dbjOYxPDkXkQH+AdhQXjyVxk9HjuPzjP9tvYOs/rY
tPqZoDHc2p13UOnM1w8erTpLJc8S7LK8J9YLgYFAZHo6Kgv8N54P3ONuB8vLy01j1KSc/O+3xqHn
2ul+tGJMgTfrhTUZkSsyy0GT7W/bGZtuSFjXeN/0PGF3rgv1/uudXjALUT3NjkNtZeKgEnDk3JFw
tcnz1UAYe/vL4wPfeFrBfoUSmLIRxxeyZTx1OcDqU7UvRZ0k+tmYUz6UktDNDq9EDXcjydrpneyi
giOnZx5NRM7FAiLVXQyaLpwz8tELjPJl22qy4gsdQyZlnTNy37b8j/R1m1v4xki9wir7zelDTJIh
WbBbCwMegb2hCagfiULFvn6j26iZrHiCn6BLlZWAZnfAwYmQQwRCrMaL+HzPUUjYWD7eZQ17JRpa
JZHz0IsLI3PNyd8jL2UvxBZZ4fZtqCxZhMuMFXKpyWJ163kbds20rmtoKZ6HfdH5aq4eJrUEvnBO
2wHmehpakBwJNJy0cTlsJZ8sH1FPucCHmzMG2MAUuNaWu9TwUSkec0wn0Z59XORZxNU9R3gDCLRi
SoBVKb8rP/2pZXcHEAErre5Qbs/EhkPU61Lnvp6J98mJ/qG8o+iKgzfz1lqoeQDdlpX5+SMhbaDZ
eEMW9zxRcFiU/rXFA9UNRO1qDvhG8v/PFE0z1U2RQk4PlsAHaMg/DtXNUZz/Z+7aUEtfXiLF7u6z
gczmMm0psmvVIZWleLlqooKSytMgvSuft1FOdtFzSpY3s6n1dmAzKu/R406A9x5D+R1H9PGnpjaD
mZzE9M3XCAhfosmMtTC8qWrQ7JLHQL9syzJCe9ryUztxcF/PdhiQDPZlfQpzZhbeA1w2v2LxtbUj
Jt+wZ+esww3PwAxgQ/wdh/8BVfPw9KWGA8iKJzdagysgtklJ1qtiiqHB2atfhaHWmJCqEOCSnB+Q
FIIUlL4cwV/xcgwMg7GMT+0cZFplggVeRKeKB1fNAVzsdH42OId9T3Eekj7BiOpl4Mg+36RQjRCW
K3a8RV/oyGd1DNp3U97L4Kjb5PiXs26eiCIUqqQHkylW7BVYceipfOLb0CrNpggbunU6UaaPpFnL
/rIXORXfPnaMaq7k/NQwIo6KuWylRJ9Ame4CoPl0FExvMhzy1fBEAlGu30X1CosRW6FLxhpuHQYx
XcY8wtTu3MiOva+OOjveuhbql+Vw8+WIb78pi6KRbPa3wP/LOhMRLLXM4qcbjfa8MjuJbdsVtflX
u8aaDqBi1lyqax0TZa+fCHutwE5zL1SGc3078zuF9HsyatNQVWgQT0dc9PxCQsXJWSNXXa0HW2s3
5UMCZpyAr+A7miZHMB9PZ/UNrGHOCqcyqLctLCOyIDWCd/RCb0LM8lyhKzvGmMR/VFJSratzTywY
yYOrQksKegDA+mPv2iUfnZBfjAWiuuNMTn8sFe/hIcUW1e1n+Ak97inMKh1lnUe8/smpXnSLbwCC
QHA1j6MoF2MuAG8eA/zl8w3wikehcsqfwOQgpH7iG/wft9oD2MQuyXVcPEM5DelOrY7umLfmC9Pg
Q7iXv3Te0uNUSmYnplSdyGS8M2bersv9f43von5gxNJRcqrIgu8Gte0OXq//P+QrE/MRX8QUW32I
xsrJd2lwkjU0RH5S1ZeFE3eI9EPIA/+YOKqx0MvbSuxqLFys1sU6Dr23YdiyFAhcfkp11UHlXcmk
9AB9Y/fpI7tUeeMWGKBtGCdX8VyV3p1Stw0na2fjEX/4pLun7zAkLRU8ApeSUDO2Fa7c1GnsZ3s2
6BDXwBt5xSM2mqzUt22BvNp1IBzLo99QC2d4T0BC9pciYurPWu8G/BbD+CNC6ML0/7duVJ+h/aCH
R6ijKT6hQjRwE/8o9c+Xqs/us95GBqZAnewDXemWVIyM7ci/qjcCYYPQASH96vLbsH2PhIm6j7OT
sseZ3jG70jIH68LBLLfiMz8SYro+kqcX29P3J3LWgxRTq9h76TOrjKs4OnDoIatuZ3faCjpT7xKv
nzNovQeD+yFQFqRrzWHK6pXJ732BUA2FOlz2WqzCuH92ciU7I+etrP+sfzNmCUzm7uydUi7T9ylj
SNnrfvMdrx1pCTfbvQ3zQLUhclZXKVV6wNBpelnZmlKaiwiQ4Hi3H9cKd/GBGjVzw0IG+nvodA8e
C2b20bvxsEEuS5wzfjLfB84T1Wf/FLIPdmqHODNA1xG7jCn9uoTxmFjEz4bhzaZNT4Msu3YTc7sI
H3o9q/qWrUQVLw3MkXtIoN227rGWjm05owYkiQ6HM/q5IjJFJserg0p2yFn73q9IIHr0LEok3J9c
rcTHnt6hw2MVZGBfCCaQIG+hcZ2m2bP0rNrvgPkZl/5EUbOP2MqX6Cbzeb1BUMRqxSyuhAPGVPXT
m4GILpNT2KLNCLZP9aWXEJlruMMMl83xwNKwR968fRlI2hO1UMoYE8s4Cp19wmSwwaIYAs8q8hId
nkG01vrMeNpjEcESSTKT3qI2FBnKPTIRXQXIY62G8Vbs6PmFmrkYaIo2JLjmYPalAmnORN0HiITi
PjvpY+JvzVzM+r+KJtQ1awDpe1zxGLXH3Bdl0s7hjq+Um+DVWFa1WY19SpWo3TMcr9V2mekTW8Gx
IyhO3x417zFmjAtzrpPfB48ZR7khea38y3oH4J09hAPckwEWTuuVwDX99kTuoNx4kMFghnNBWqC7
g7JZIvLNevJ5z/kTxe9SF8IwDnRVQN7b0ujod0tyBSTOdZVOV7xjFAWetsPlMK/PmBpr0le88UBO
SujnYFYoXxluLS/YkJwIOD9yyeskDcnuamxlXydBeyebwnuHl5lQUqtfe5Q9SlLqG42+6uiCEpKr
0BMkKxadXcmsr+GcDojXctOtO+yEPxJvqRqe8K6K81zrrYRfn3FWjOuEC8PhM6TpvcmZ+UYQCmZI
xFklvBvE/hQTR8/tRESMMoMnvBZFOM50NQw9XFxibuVSRd2vG9cIYfB1xKyYZQo69StCei2V/FN7
YgeIJHTDQkRftZz2uAAVAzE4dW8PBDvOF7DpgAQcdCqcF5PTVTkn6n0pwT+obFtn/di+PDJNCpiv
UZ2jDsX4NFQplNz+1g/yq1b/WVt1G09z89sgcKY/4hmruIUZozTRXdYueOC69LVCUZdAyodJQyMe
e/W5sc5OKoLdUovjRP9FAk96CPjc/hLUWCHksHpDyS3EZrIQZcucMOTIlrfduvsUTcbwQXYjGMEW
PiybCZ8l/8b4ZfN9gTwefUz0ZJ1skadnI4xNtmVeaeVoi7HaJn+PpcfQPETQn04UkRCnrCz9xzW7
4YIwlcEG2I7iS/rdNblCVgloc3ZXNBNMw5ND90huxNskrNHfRTWf2pMDSayRV3oXRXa1JLCPWHPu
dyF/Y+9mvfznWMU7lfWRAHJIocMCO/rlWHngr0dSJavEjTIstAPP/Zrh3fps70BKFwVMGy7qyf3d
HbiOC4wHj+kCK4mzqVrHDT/H6JlnKQX//UDjXcNaqX8HZLqMT/cI+rhdzT/f1chhoaNI0ih1kc4m
DOR5fWqhoVNZMFiZhJEOvt4/nd2K7RfOi9U7p7K025sKjJC1xiucUzggIKM31R9LPhIYDDxEy2sK
lh6GxzA7/DtLu2vgoCpBYwFYiZ/JzpxaAwY9Z5xgiDKNSsVnpaXKNxxna3P9m2LQD1m+h9yAhm4K
7xXiebacfMZY/hwIk5nMbAnpaL8E9CReN1BCofOd36eshs9fd92IHuUu1yvFuLwY1HSc/2LSgaCK
TNZ8DsIqGeAcl03VnQZOyIvvXysutVTQ1/V/6eA9/GXHkr/GO5U/HlwoEl91dp+Xa5OuYHaaGDig
aQn+WqPU0bacSliEzkEUAngvdkTpxl+GyTwZAK3W1qOVssngZy0uE71QATkGyXFf2OGriM7eZlKh
8aNe6BbUHvnCxdmGpdEX48SoXKlPYiV6GFz2eAutq5g5aMXK95u7+LBogn5aqjeveNRjLdMubgoZ
km/kfXLaixDxcO0ybzWsm0T8mt1McawcM76V91tAk/r2XG3x772zCmfjaUh2MuIE03StBYJpyIcL
HCOvsLmRE2qoxIImNjLiWDEiDCoyfeEbvinfs3cgMoj/6mcheUbWdSMIPdcGaupSGzqcWlC1ClgG
R339/mABno1AlfSzu0aUug8vWIR9W1/caaB2JPwqEtXspLMk8Re9aCGTMZ5Pp/ZbW2CYe4m1CyFd
E+3RYtLcElQAta0/o4hB4fz5MqsixhFZgCAHGJmjQgw9uRSTEzuQQ5RjkBoXTdMosauJXXggFx1Z
ATCNzyccPuUZIzUc9EW04qL2xbEvSEq8Da1FseECQFfhqBVd6UntGzcN+0s3hkZPsidRChWPFl1A
2F2CXVk2WvSL7PTVR81MtRwZUZY5+DwUjs/i+/GzEkxiJBDMh0stIm+IEUX654NiS70XqPzcuCkw
hOQeSNA/tHOEsSBX3GjInWbPA2dBNzpSKo8H6OoEak8td9NtwuBB0Bx+z9udXCLQlHOCNqjeax/l
oS6s/9vYS7DTPA5pqi8Okxr0oWwaRKttmkOs7nQeil5VyHaZT3t38JYmOLWrnss1TxyAw9lIp5pT
0QpsAAykc0uTZuJ5xXFojSA+RVonnDCjO46MD033+Mc4gRKhU4S1iVskZq5LVkkbwRsIp/Z3fiZy
YX0CPCtD71J9/AIm+Wp3g8JBddP+/2wKfFDlnYeO2uihFl+9BkYRHXlhphTpexj4UAm83obb0nAm
O1p4lP/6EtTTRG6C3Vw2gDZPpgJs3swseb+vhbPcPEpD+lZxNWkH1mj+Dzsry/a+Ms/ZQ1xzScYL
25nXKLhIHavIxSqPSIoAKOR3FQ3pjSyxDyxgPODXoCOkqXEYFIHYTG/uKo+0oNY/Eax8x4ZUgpYr
EPmsobdh8qx7nxqywiS0Q8qFC4lYlfJ4yhQcnP0YSLEYOfPayOjWyc+gmktTJkQpHeOVxfLD7zIT
01UVbtA1yZMnApJQAk9B33aCCYJ5FysG5iym1WZDCtfpjrHFrDQSmfoa8jhT9vxjXYdp/kuqSh04
utUIrNDGHqkjejST/jFQI9Z4JSQb/I4AlLzvl0dwZaYEl9Fq3wgwwsAqFLWuWCAEr0XOJVH3O9Wf
UWspv/yNblwEB6LhTZB+8xCkCKSF90SzpJ5OH6TvcARoOrCoKOximMtK0wNahGPsyPZWZStXuQ4i
QlL/cA7WsQT5nZm1UIvJ5YM2ZQunZ069GG8S0tvXLTY3NMZKoXuoAoPLdXyHsD5zqCHnQa/jNmQe
vo6MkENfyPNwBE/OgGes5wr3pgphZodDz7js1zybDUbctLF3D3vkvN4lw9zXKthKFtb2QUaov+u2
/QXDXQu0Z6jVOlmNCCesfkcejz7SkpBjdSQXYzP7LBQypCW1LcdL7BwDu5nPaRe2+I+LjFn4+onR
pFnhw27SFiZcB6ttw1AysJeyygBGeyEdkzjR3aWfsXh3Lf4SC/1BAb78FIUyEDMNW3BWXmWdvwJI
gKaWX4akxX2RjpopNEDYvSlm1P8XQLyN87f8DrHD19wfP2PVCgisKr7lITm5QPo64QvjO8Vdpa0k
LcVx7n8FYYPfxtlKHw1g1y5yFXTGGicsjvY6/N+BWR29PTLEBOHxOiTsbO2n3srINKk5gNF5VFPX
ZUnHjy4bFw8oaaYjaDkaYhiOJCBokwlZL488QCKhQJj3EAXLICrD9eIJFwgWGqDV1Vs+GxMwnw6j
13/K9JK9i6KVA1MxNJUuco3SSt0h05zo4lD4E2yfgMXHbgl/KitCI4CTFL9bc6so/n7GWmjDHayP
sWsz9o0jzTWzFAT5ziUJPefkbabUshyW0dWf9nSsVnv1a4JP7Zj8kg/6H39Ixde8P5eerfajAVKB
pQ/GQvuI+IdgBAmAzymtlL5kCf4zfsEu2rv/ivire0+/Mq3IatvhnoVBGHO/ahu0i1k375Z44CRC
nUVgurm0UGzExqq0dRrcuQNK1+WBtYES9g3vAbvnS+HAYa7BwikMilml1ShwivPd7bylBXOIAfqO
mSK1MpB5GhBOmJ+1Pm27z/vdS0Y3yr0VcOOvaO/uoPFll0rjW34Fobp0LeJ2uRg7k0lgYbmcb6Y9
zMPd4Khd1bIDorm/Hx/IZYphzjUJhhwe84gzXPf3UO0BZ+C7E/m2JEc6inIwvbN+Ylql8SGp/VL1
LVAgjGoYiTHUt7Uctz0nSYXvVSiZHX5AjtDUPAgyCc8uiRa4pILkDQtGY1o0LC0Deu8DoJkHAPOt
MqDc6oN0PHVU09jsqUYhPL+Yt6OhU0GxiDkoNbMqxS9+dOt4CFipqzbgiS++B2jNv3ro+spt0/gJ
qY2ON7YJSAk+PGsFMYQQjID2m92f8TcjO6LbbeOpEsFJ+pXb6aHtbRAPm6wjd0g/Fwwa5liECYUU
Nv6Ku+J8CDvp+mVQ4zkwurdE/o2k7tb5sh6H14lnI+jF/H5C61gvQXdSgh30BvlooqdFuN1qd+H0
lGjoPxfctIDvba0XyzkVJjP+y589Ey7Mg+jKMgqUR043DYqJWf5RUcaSmj89tRUfuArCsaJVglCW
aTtCBcqyVy4IzVJ55ZKdxva80cj/wbtH2ijYxJFEl109LxK7hIYHjw1uhd6Wd1o6/k6Aa7xEJmMf
MIVIxo7lBTcipx6yiyMFmK/DupBBFC4eGhg3wYFIUVsBFwhOPwmxOe+qcomT5GGH7cOkpYv//5iw
1fgJn1mFxNrcS6cDVun/zY0q3gv+Ss3kf3M/Lk7XtK3ZQ3NtZBMvtd31/QEbq7p85onMRNZCFvRa
18zb9bZ3UKuJ9FYaxjxIUqyYsI+F1P8XZCMi4TcHhj/TSylnZ67MnESKK9IPgB+mr1UM06+62NAw
87YKu4MFrH2ueyNGbcR64EExLhCZ/qUFntiKxIRVo9V0q7TrMSEB3miTez0KCaDUhnTWH/8HFE7V
olswClldJ0e7NoVj9taSPAybWf+REfoBv8ssqDc+Ljfw8QOmK0ZVa+MQc6i4UjalivQGnxRCbQNK
Qb7pTtGoFsiBAsuQR/c7Gr1kF8w3vfpOiPG3ybfEq0GAArBq+3IetVPPUH9CD0BH0a30yPfwGkYg
39UuQRwZFsd5vHCYP3e0wUxBZTJ8lsBd/ye74/lI+6YPf88UtW/U8Wcw21xglC5H7R9UfOlS0tQv
6HiN8eVK7+u2ANZURNaY2xcH1QbIUdfIZdKsi75clbW/MuyDNuB6fdLM/dgevyWO7OmUP2XSyAmX
ypuqBUePFri+5PIeO9G1RQtCSAVQQRpRjFXwCRo3w+DtFoOoG5KiKv0Epm9zcAWx76BuJpRR+f0T
/SQS0x8Wd9+TzKj8WXxh7VRlFDejHo6TR/Yq1+aJkqsdEzze+M51RSvQFwnvXV6QtZBFLEfiDbtQ
aOwk6hqENJ4UtiD2iBST5xxaJHFacZHWPPS0vmGQoqcWq8vy9Vd/QTP8PVQ/1Zq9QhIV2SR2q1k+
o3qleXeDJLN3pO/+yX2YMuJHyOjXgReurfLLQHGTgx85iG/cjj9UbuwV2rzKw3Y6Ql1o8CERhwhc
dvmTpieU52a6MwIG+A9uquI05PJSw95WleDRCwsTgllEF5pGl6GJtPnsrtQyQP27875lNYPEGDt/
CWbkoFdjBcfUbUZEeA0msO/0NoD633R+UQbyTk0FKI+36nMGovk9QZUXpR6z/dM0cNbd+3BKEII3
dZAXZya4zQXNbpvEFmRHwFVuXjx/hdjNOdbwpGWeH5itk58frama9C0S5QrB04t7MO9fqoObmjqA
DzwU01LeJR5d7u81SRkx2AC6SzRsTY6oOk9OcfpLh8mxs1W2ucEg2qvUlDBjMIHaARywNpIQAyQR
4i4OGhaQxlMwBt8JX1aZYMW3NLmzoI494BEKZaIJjgbdvtg1+nH8xdpQ+OTWPIfiOtBpL2/dChTi
yffb1vWWzDVmz+idsNwwq8H56jSFZ4SwKGOIadjx4KcP/7LRaMHEbbRC24RoH5HrDzlYxrLj9/LI
MOYxReAx5qSPaYiSPVkQSZ8aJhYC5ulo4YOd6cnq0pNN1ABr6Y/RfgHj/rhJHQAecm/vaDZgpVH6
NbQlbM0stunSkUNdZ9wExUO36NwqlohFQK0g+Yhpimmevs1AwxFnSOrxTZHSs5xQIOqSbYhUEJ6C
PG15Xtn8/g1DhIOk+VWnhEsIssPBiK2gJ77eVGssLkQ84gtWlh827FVkZ92oelJ/wm9IL7ER3rWK
QcaQKXylem61Mn4oE1/w5BlYiFKgHoF0KQ/T0bYgtUprmWJM7Bx780DbmPk9onxL3ukAddPJclnL
7C47PMew9AAK3ef2fdIty6Z5MlC/IgtRPg3qe/A1bDa0F2Ubhg15Zn0YCLFWhlTWq5VoweRwH8Om
xr0+r5e0UDpleKNJuboeUkFfC7vp22g5KIploqV3AH5hRcUCjgFpG37sm0NGxet+yw5lobTRV7bp
lvLOTQisKo7YcB7hKx1zXe6aV3iyQS07IWE297zGVA3Mk8srUiKP2+LlmvoJI5DhwTIA4CqHrZl5
XhmfLNMvX5GOBXDc3rYxVcfsXydRnMgaIEYRaRFaTXi778ReVEERGBDW5XgO9FhzxRBxnF7Oi8Jc
yXh9mu2QEJ7nSAlEZIrUodfP4YtlZ+SuAgNPp2b00kFI7X1r3tlQIMZeFIOJE1pcduDRCZfExmE9
mScUpHCl4xN6N0IVsewqm8/HDoptrPII3X4o6VHYk5n8nd91S3eT3UCMC/vFXotB8XHBATfh8stk
XU4MrHBOrD7MIKVwkmVEYHvdb9XzpoutanDWlekxIEm0+6ttB417Gr8sigOPa/qOSEgbLyuE5sRA
3sKOeR06tyhrWtNq7uaDLKZfn4BHvaBPQQmxXV5UGasty40FNkAB9l6rRvmEFayJ05w5kTWfdWqT
uUdcK/e0KypVZB3P5kAzxxMbhvdXf+4gIBEtQrWzgNXlK3D47Zf6vvEV+qHgfKo5yEeWgIEUZxyq
nQknfNupAg2PfHbZoSVyWqZ3DZmDAfSnFsg/5GxMkLutaDC4WJ3b/xg4InEjL45tCMHNjIgpzTHs
ry2uGZnyYnkeZQQV/NNoYWP1BB+py1b0CGlaOJ1vStCBvQBqgjxmt/itcWzr0O75F9mTDoSGALE3
9NiM7dsXN+yb2N1wWsVXPsshXZcMOif9dNk3ZYC/QXsdmHk94IN05qm1EBys+aTVGI1KQynYzu4d
eQ2JngrvPN2QnwANEtRtp8hFPEhfAd0UP1dkWQF3jOcSzz98EIyVQ3R/i8tU4Eb9KabiWts/vxKJ
IGLesG38my9RqcATW2pS7A7JqUfZ+tojTE3R0e84pn6I4bYw/MP/qIAy9amtmes7hMJ1As5XlrRe
hCv5zdF5M70irChkZSmER99T/aCvvJXGJtu8ktQ8aOinrMYOVMOtj1fo2YuNW9wOa1TslR9yXsE9
v1Oxq9+dHkKBxIBWnTd8pgOBDUyZyo+UixeeFGlJWmSPhE8422NuDTqK0+i4FxiF3fezf3GSOE4b
ou3Ktw6saTTnOPC4JSATI3RXvD6mlDxWAKQlBxbQa+Lc1PzmO+7T0Xu50/9WH0AtEkdC7h/8wnR7
w2H8r1jGhBux7tKQyY3DczpotIpLruPKf+zBIp0lC40U6FpY37t2Y5IIbPv1G1G0sWJyG9JMvkru
BrYyzgSjHwB0rdWzr9SJ4uPEuFa8Bl2oZ7ta8SIxOCEm8spzUxwXxjK7FIFmYzf9CEGV4wmaXEqb
rFiq6SjTiYpH+6psxX1cjeMh9CApMfAIT5zfeJV8l9kQMbyt0XB+htlwSCDEtIbp827OU3spCqhD
wtyuf45/pP9Ww/WDBiMQfI1fEu4pdVUOBraaGKI+KEPzY4ajawDHq84/uAJ7+eqmTo4PsV6OzdwD
KWyCrXBev4wWfLbSRgtRASfIMRP8kR74gkg3tWiFNWre+eGuX6VlZM4LAAdxhY3dlb6ld+3vsn8E
yOE6m5rfedSSYtbe3KNyT+0CgGlyVl/ByQSxetkL6eUfI2EdZocnfSrhLAXPetdwlM2gZOS+HfV+
UQaQdfxipbJZx8Z+UE9suIsPtyNqvS1BdircyGjD4Il4TpuYm8gWY4pjVtOSBlO+3nAPyEOT4AHi
gNCpoUG+0IaDlVHOnLxyL/0QAWZK8Dsx6cec1BslQPvD6VEzaC3rdASP89RBEbUZdHitxr/4lEHZ
5bk9TQXA2IF5MXFFtCn8FPaFjuZL5F1XKvkycjrw7A5ZjIvaWZJCmgtL2AcbNOzWoAJGHgB/va7+
MkqNYvO8iXUcbyvNl9UKV+qESdCt2axO4veDt9XbE4+SKej94Inc9Gzi8ULfrGJpyCXdFqkR7WLb
4+SMZ9M+D6855951jw80u2eMx5gy9zhUX+ggxxF84din5VjnPv0ZOuU43FMlFIYtipAXvMFeidWq
61QhUWa8P5cDy1BIUM2mM5oPxDm6nn2lCAYE5VNOJ1v6Lz4LxNhQbyUF6qRf12kTtUxZ+Z5LHQEe
weWIvn9OSYvfQFod6afMwFzocG0D2f4yPRhZRLSkMml7WztxVZhdbuErQLnKt+aOhqaJPEyFpY2/
EAtOxaoQjBDSTDFhecnx3L3IBuDe4SsI5fwM9zZj0XOnneierkuewZftYHhpb1vWJIjM5AiUoSKp
qp4WjVDR9SpJH8bmm0j0XXXirSBVIEzRyN0wB7x+EIhGIpqxnTqMNINu6RzsXGHkXTHX7QQ5vSSv
oBAhT/XCOxriVjQnI3ADVDi4gzrv8yzksq/GG5IhyVS3Z57EyZLOvxxHl8jMii3/la7pGCzBDjax
3rWVDtHw+Z8rDLBuYPjH1nPB22eA+Q8c0W9KsV47LTV5+cWeiQMZDnZ+mWfhQdXlwRCW9r3J04T0
bWdtSzntu5t8Ms3tnzn1UsKYbwGZc8gl9T92vEQnPprvzqxk4thdep7tiz/GHGhGU0s7GEmViudC
CwLV+WQKehqMaAgFb7+ekhDfXJ3AvIam83otMTbDDi2lamP7r6XPRpDdZ8twSRkbi24Eg0GUqJbV
+ogCUevove8m61usRV+WrCfVd1FoA+9JCQyZjR76F1ezCgkoGtJfkqqXUuWiLYvaeT4oK9h1eE5f
0P8TwJk7DoJCrg86/+MPKRfQP5qmqweWRnE6fMcXkN2Li48LtftTVbpN75ykcSF8X5IjTii4vJco
OcOPhsMshBAJc3YY5OfwfIpo+Ium3BX2TvhVFyjjfqny71n5SNW3h7/CDhOzixuSjX9m8KrCLfg5
IurgklaMPrLgWTSDaJSyfOpc82S1jDDaoi/uvD0XnyVLgxdUYwX4Um3+CMpLEl2pQvDC5sLy1KQz
1+L1ByESlDCq+2A+OKXbhG22RzmTIy2DGhHIJKsWR3LxrWrFoVsmdNmCYtokpaQj5u0Uxdv1PTvI
PKrmITFOmWzz9KoY3v5jUBwiVkiCUv/UhTiX5AU+1xaVHfAmwdZCxJwuUWqA6R1H7GfrPYZET9B9
Lwq/FC1u2N5v+ranS/Wub/q+BdZdHgYoozNp8T9cXjl5EHwsOvFgBz749qHUA+9PbGlMsWRkdQHN
K0Tpi4l8dATjwRoEPfNc9PkNbWEKPGXRRI9zi9Zj2hyrCCC0Y5DYaqLLhbj4fw8cWtNMOs1APRGh
+OMmrk2mwV3qdUtksrI+Ncrssyr/HJKdjG3H+Yur2n7d7mcsHY954w87sKW4wAs3RgyU/PD+Rlg+
E7xTyZeY2W/qKrUDttMKBpGI1jPgxW+1Q7aUj/rxw8YKd4UvYB+8JCnAoOtY0pUnod1Dnxm4sohL
E7jYhOfaDYwCUGiEOBNuJQo0p/tgzw4TUbfgb5caoVLUxZhln1GCDGdBJKyILLMva3tn1Tv5x4DX
UayGo8bn5a0RMyXYBewBkFxhe6KHsjk+X370uEnSAsz0WdYL4GuFDEE9dGpzi9/y2+RzWfFlgqfE
mwj3/9UsSf036aSKs6scjwgV4okmDZRs/Q4todjC19T719+yPN59rbxDqIircAYBHt16+NiJi1ce
Z49OTfDMdIapdP4oMbOBh0kaChHY8HlZ3BP9huXI+R/+HsENazN/vN1vK4JEQ5yKsfaKQGvopoY3
FTWc1tBZ1xWI+k3BDe/9bBsKyO7BmTafVqthJXPsCX9GTBeoIXYmT6fJpTyXn2laoTvglxFowYIX
2sqIF4inSWAgv6FIge9GTOjneEmH6wjfBLya+CzzaCKIoZIsl4dDhB5lO63xYLiKIfI2MoWSvDQq
p0gXRewxkR5PHv5DgBe4AZd73IHmiQTNq2KtlWxcmeZa9EJycUcttrCMloLB23flhUN1k9G/PWFD
5dXEpa3JJz+DKb3y3UfXYRksbx3wSwZWm/rou4MOqLYQpRCCAECR6I38ZiwAKxgyotvQfivWjxei
9LWxfLSNL6uHSMO2vV1nyP85VkUgWbsx6ycDw3XA5+sybiBbxSldlzByyH8xHVQAXiBXp96/DrUj
imw/eo10iffGoJzH4VtsEpp8eWDlmyYBrIHci7qeXbjrepiZRigX31yR9k6MCOXwY8AGZJRLJyht
cNrmypIepEBlpcnoS883rlzj6sXcn3DjWkpjbt+5/aWTdAx8N3tTupHcW62nV9z/r40+gFT1Nl5w
v8dldHMC6XQY4SeFu2J61qgEc7gBprfYEPHVxH/Me1IaTv01gEgFYOer6TqWjL6wwdY5wytk2Am+
RrQZXMIhvjNHMg8PhVzghRuIpm9MADSi0zluAwn8i7XHsBaq9hb5gq5NHSXdbMZ6wsC6L21D2xE+
ZLDy0sRceWgMQGA1pNLm9XbXdZ8rsgakuj1HPmEDiGTKxb4vNvSOBBGL4Ta4yG0Ok4CqsateX+dr
0jN3qOmDkFLLlfWGOfpKDYEflnzHh2IBiavSu33UGWIPVz3gbVifiAbMJA/lvn5ACz9k6tnNmhPP
6N9+NPTiK493vtaYPHHy7siVvX3JmjWkPKzHxzepfAy7fypG9BcpUQ6AmpUd7apkN/P4GDsZmvqU
/dARVm8U4K3vbZEoiGVnvObnDIwWUgVM2r/xM/QI6OjMYT+8pH8MPsV/tgJU+8OtXRFwqp9g6UqB
b2j5mHt/rnC3Cm+0ocO+HzCjXU4C4WuDERmyRE/2e92boATTKaCnMPDIVstKB+3cQjhaBSA8xFDu
gu9otBrcySJBd4g73kFWUoN13aHjueKRtxN5+DBtbImidKBLvdDxFLF/eH4r7A2+tTS7j2G2Z+sR
wcSwTbP/6QW4xey+OBKVy9W2vCXcddNU8OH/YGpYDX8TsDbxn6xg+JV8vJn/zvzlzELdt3NaK/sP
RuI7AhOy0zPGteB45CZEkDq/lBfoMr1H/TO/CPC6bEzhb9CROXDmTuKB/3k9A3MLH8smr8rBBkfg
ju6aZa+aY4o/y6T0pZYXXfO5bLazgwSR/HUuSDkAHBDpG6qICaAEuUCMcGpJIJdyd60jQVSwYkUA
daFWMwilruxqHQ1uK49GQmBVMJphY7fX+uqV68iiY7CMYUUF6/BcbcaztB+9OeEpL8kYLICEyV/2
PpmGxv2CK7cABjGWSnbDmjO0FpzdB0hfunPuWtzez/hMRJ1srXpiT8IXe+p+RwFTWp6/rtKhHL+U
LGCgtsETsFnI9kpH4MpffLk6NIKiplZI52ZClVTgtJbG9mnR+FRqZigjQ7HcIzdS5r3pfPOT5sRL
Utdc622ynnST/CcGVc3tZ2O25ej3tt31p1/QnSNHao8vr6tfxLgCb5i8MDR/fJlmmHcr6qe3hsqu
CWv4AqbharP2sLhdZQQcj1DDmi5h7Piila6rdm+k86V22QfUv6/Lc4e0PxS0+HHhzp2s0LyNompd
Fd7c+a9iDoOiNeAC12++2yFfrpOO7HctOH2ADDnTOLYbtCMqgYemYbdQuL88Am+h3XcbO6FR7aj3
YHIbeOy88JDt/+QzKqtriErPCkP8uzwFAuSexXwmYOoQw62E+0cbGceP0B1+Z2LMmkA7Ny2aAfsR
3FqaSFr2o6OR3qdEPWqJYn2iKftfaxYi03F6KdZ+j9a52Li1aPNKZ1GjD9+wR7ls1fp4WnAZYHOt
4++1zzd+82XCVpWI+4G2KERId2ojnuEMtCSR6HKJURD9blqa/COz5hhrV3cGYpkahPvIGPx5caqS
WLDQ4dinC+xZMlwHddkC1qKbzkf65qpY4xP60vkqLD05dFGSVB3/1oRsBu2aLxSopYd3sZJWv1nM
7UwsbDVZPW4Wbr5IMzeZFuk+Vbb/fO0qnlcHAmsxPsMGzzKWciy2ln9K2+ca+qJXVSh0ubAzzL1F
+NxYp3IhYH0Z5i8zhwcDeLJxFpB4GpOzuVvUtYyfKGzuf8PRaANTDt0g7Km6WjfjwfmhIk2XlCfa
4yPpbMCNsG7LAw/efEDkgaA6xZ4ErOEGQf8oXkBtIz8pvjqrA+ym8vLbYN+6uvG4U7NQnBxmlk/m
J1sHSEK9b5sSJ4OM/E1ytmbWEMzGioaCVJI0VO5yBZmpB6oHjnES3/bEIcXqislJ3vJPNWGEXIw+
o+1sh2Jc6q1dapk50fvfhAz5A6zze2yvY6OjqG8rqhgXjY5DZe9FqXotoqIzKPGhm+RcTNfd0dOj
OH2gae46VhPugl4CDb8k1JTjCSyGi55EyerHOg4FYGiWb+Oa06dqKJnZyYNqrmBf3bTJ9qv5QgtL
RuAHNNzr9LhC/EsZguInXDqIbOKMXtjVOASGaA9PzG+mSCxCRZ62g1itUUSmdQo+Tz7Ge1vvrfpt
Js3SdRN/7htMd9iQe9rENmLJuh/GnHoGHGZeLsSQjVGWg2qzAMF+XWBNhn3tpds5tvZdniJ+zr5R
FIriUtfrTzcSsSWtMwuCEzcjduP/TYV2dfLI1DC4NK8NENzBtmsLp8B23m0I+tyKT4Wg89Xzj5Xa
hrDjT3ZwYLs8m8nDn/fkyqYLOGj1kNWC1Doq5lIsICKke30jESHTUVPnbhHOr/IqoxI3QlyvFSZp
NxKdvGne35kM7l5AoGJFMIz3lx4aGXm+FEdgHrWmmJROSODIBKfyX1VdZUzNGoR6Sj8e59vvaYEU
hO49vAFvJxSoqtFumfod843BNbwMjrUxGKfOo228qz61e736XR2TsdveMcFEWi1jYcrlfsjmB/we
Aedz100X6CJOD6uhbOKVFuSjNIVv4xxc41j9ponvykB4zILQOWM3EHBE5M+9WSR+qdxGaoyYNW8X
Nt+ICpxNjMN/GxRJWUYlNTQgiU+f9KTXTFUvN/tFaIsx1bYV9WxcG/llNsLs+ET95y19YnIKRrjm
7ByZ+2OM9ii1ZJ/JqchTYNN5/Ig0SIKj8TegSyiiSFfnk7oswXaXXFnjl5LPEGfSJQrxSm7GT8Gl
io2DRHmlrI02VomWxAD1zgEsDWS8oFYFPRsM3k8E0kx3PnUzWXFNZjzLckYGiGXfijoTkUH25c4W
hACe3s/3AX5SBnYlSRbLAQeRtsyu2nEsHHcZfMwMqcuI0a5PNBAP+cZbhWzdPezgfWTtcVGBQi+Q
dTpNG5XrFryQStCtybsgbXXzi+zOxImXq27cTncCTi+5QI7Ee1JB4SoC8cOAjnmyprP+QEIf5SuZ
J0K13OJBVC4NNlNQpNJisRw3LOOSmSnIFuRTId210l0nZoDWTV/5B1cgu1uR3RO+qZmDTXyuMjed
fleqcsXBKyqLpQBYFIUTW1KzUTIQFTeeY1gLxK1EqDqxhH5sphHvaH1gcfkEn5gbu/tUwV8P5mg9
UejOM8891hNK3VnKKRuFcP6lLWUJowKFBqzu5hRdEf/FGX/LOoesGysTHhPEFpCLOfqWx7VdRZgx
lWakzPHLeTKM+bv6Lw1bp8HTXzzHoqVykf7hVIz76r8KilMxPeOx77f4OIQrkWWAdx453VBdii+X
+K2fISd0hEPBmP4xPzphIQC2K3Hu6HKko6axsR+5apWkwSIxEzDimuavHQa1V25WGVXMb/yNS+sf
oC1CTCul48jozIjr3KWnRNRUFjrA09deecRGO3q6kLWhvVB/km3TTsTe1l+uLjwKLHFSJfJDkrZx
Jofd2PDRKtr1DdxE1fw+tkYuqT2hH8QE5VTCiOPsWoxvdWNcCCr4fDqPX8Ix6roJgdQ9iHElvRqr
q6y3FcjyyZ2FyNopEiNY7ggOjPsz/l8evJJIdGDYl5QJZY7xqOanLhepcaW3evrgVagSwhpp6R6/
M6rsY1gCR1cfuxtvMJ3oWF1JGk9WeL0lHrJlt24pClzYhe4lZfNZT6leyfm37v00Hg5frYDCDrX1
CeanZX7VqQ85lVo8Fa+FmRS/pbFgvX3Sa5Omraq4PvYedrv7qrX+eaRwdYGei0xWRekKU+YMo0qK
uB8Cz6AvjgfUzHBoSoEnBUvIyPEHiTbqGeH6tdI8NFwNiQAowu9C8LDisC+B93tR6aZx0yhMsySz
dRezA0CacsSrQ+coxB05ui0kmp3tunc438Ny10uVhdjIKRkbQjxB18rM3GXO3A8n9bGBH7ooEA8P
wUJmGsm9ihipctL3koXlzF1Lcn0ypp/BkNWKJqCjXbEsV/vsiNFtD0m2k3g+Hnmk/yuBf9NIlDIm
Q5i6sSD/M7U5DKgZrPlUeOPoLYMGGfdkwVEZ+VqBC2k4XQnGJV23n2SGyuOhvnYTR0xnczErtOsd
R1dCGxVg6tObHk6/acbfaEzExvCCpmBU2ajHqtQu8xapo//nGC5EekmVGRkcGlMm5iCmp59qjG9x
7Hu3Fyy5IXyqVyOWApgh5lOXl4QIUpHw/qGhb/K57MY/LoFYAXQ730rV1n1miomOMBBC8YBq47X4
hNNiHTj33+Pqd8aLp/JucgtpPdkyFLkN03jn/zSgiPotCcRFGkV8PNVdMCK4HhWvy7nTUdtitMaV
lpNJ1Tao0u206r4cUYP+Bya+O4cWZcQHv4zd2DYHkE9CsGgUTo9s5HxxcEJ8+/CFDANH7fB/EfQI
BmsHO2jusdGi60GEnPmx3bkLpug715hXF3GUUBVZ/AFLWi5//qfOuCosTUfwqzUMVf5ZpDBNBe4a
vJAcGjiN+ejBVTtjPeERrH0iRmPbqv9ZuIMGPz0UQiMLgG+Q6AO/G8CIZBWpL/KY3nWI9QAixplw
UbKgLokIA8v/gcem6YvXuSFMuTuvpQhv4EiArXOzGOKFg/H9+i6qWM+qwm/JNdqGdURVgAV8EpBv
V+WvZpXeqSsCXookOcpqH1uaJFjd7lprKO1rSiDhEHOlvw++zuKuEMzM8l3973FA0GaIZFedfyMG
NXcFpmT98ZX37Vm/o5iEm0SpZWLdstds7vOrjIqdhvWu6aesroxCyBCHd8lQ+o2sPU846ysogeKb
epcGcpGDiDY8C4vTv33IVn91FuoRVrU4XV4G/eZJbCUJIztVHwNx2bnkOY58mX8QB4iRXruGumuX
kKWkZCYQD0jNrUwLb38oIbDd/gz14EEYzGPrOkeWcnVB0ApOpLBcWx8jGoVvIbkwqC8SV6k20usW
KXXEoWgVheNVwhRm4NAnNcnlbj8GwVjdFwpiRvYjjxh8MBPaefagcaVJRvPsFe+SkI4LHJYrcQGT
E4+UpJBYNilWNdF3BiUT0ylb7HVjWweHYFHLBhOfF8plS75GLfTWRm4wOjvgSwn4u1dVcnMch3fq
qV191qAYQv+lguppldH95JuSDmVAj/Si2C8cLMmv1mTEwZNfzZD/Mt3J4WMDen+0kTKYlYmsMMbU
M6/i4gWjSVTSODcP4uzT/v1D8/4oir7jCOMJ0h49KEOL558uKw1vI6F1m/6kG+YFR7v9g1tgaW48
kqiTd2cPh9k7gYhawkePKt8ERxm6BG9SjYbG2Ji+R7+nGS9w9PUqywzZ1eV03Zr++GDp3oi4DFJP
uAy1mWfkhqVXhvPqSUXyh8sTsPZAypJ/mrJG21JZjUxuMiOglKdrRig7h8lXicW+syjBF7EOFBkR
qn9FprZnQWnk2GT4hqcowYuoS+OU8O9ROhoTM8PhRgRsszmmXwABWSw7Neing782aIdhRDxB5SCz
vx/OwKT9WEiYv8bDDBLtN//ps2M88XwH4MMd/b7Yf90AGQnDSb1XLd3weyP04TgyQwQPDOeWIqxd
LXfvzmtdmpvU7TXwmycVyWNwkk0xk8UvIT1WcIkCFin1GsFcAu+El0trEmo8M8TBLNXYMbvRGmWp
7yfifOffiIMW5DMXy6Fw5xJWhQf5PpeGCdpBKUILooLyvrhcx0eA2BOBy8XFJcnb6HFpLxl53JZH
cdjUZHsDZlXCCBxErETgs7JuHi4GJK5eYgJh5rEBU6UTP6bsYI5PPrha7m6pxN7fzIsGKZe8VdKg
tMPhPidtLvNSnggQADDejpuZki92lpSnjz/AY26WUWjmr1cX9eljs3JFqqEg/ufdISOoNyMAQDlF
l4aVNYBy8elTUzVbltUc+zg5jwmiSscIOcp5dYZ+bkyzHZky4TttTKcSVfqHUu6bsUNRN4vh089i
Tr/IVYjxqUk8hWgbpiKkB5AbLg++1+TdhxQLSdwiYl55BW3rbeYDYxWTYZslTv+c5yQSiNCRlAd9
sva+2nYCkErHZvqQrPJ1VbTFx9AVMPxEpYnmOcfj+61bmMuqsSkHVRiymaIGPIl6jnejOVRrW8cT
BBUD4LJyKUcEM+cwNypdMhh7N+rQXWHEXkvRLP2XDwvQoBaKw5Vndf5chMPuG/YIbLVG87l4wUIL
i3Vgej0uKjquhsvDbUhd4vLeVVP1bJ1zHA5OjnlpjdYwrfbXTiC4p/EKEEDCl0jDzMYYJvnoyGmi
NTXJ2tklotnmWGbJpheW5zyuOjZcEKh0PR/HIB7652jiP0Hs3Q09HcBdd6LWx4sX6y2UqsNRi+Yl
mJYURXDZRlYqap2kbnlEI2qvoqzK1y5WIWmQpZSV4d7+C1Q5+u1VeoLNzFdynvztLLC9ZuRCVc9Y
YhCW3w1f55FugGpTJiF4U+UdJLpmbEmAYN1ebYZG3PndUpwgsAjb1oy1zBZJEkVYf2zqViqXhT3+
daROFBT6Vx/DYlkQSyJK51FsENUl9ic6Wpx5yzktQzYbj2wiil0TPIhDatK0c0VboyFzwxWhpQBr
kxpTuXo8TkNS7W6l+Hv7Jn0KgGlCViAyQ/U05H9qMgRMZEgmQA5U4YHM0Yav0crVrE60Qx5PlgKj
H3syI+fKMXM1DvXzTGR2L59lIAVHxxc+VxbHkSuQXXXfXlFERkKyQDRBQkAfAtT9MMtmAwUtTlA8
kigsVCkPzpCG7mD8CpMGsuw/vc/j/AbXVRrqmDNOtO2p24o75QN83vokZaYDx74KFqke/Evvkiz2
EHohl5hkedgh/2U6DH7rll0bchviPhy0tGbKFMd+jDrwof8q1gsiMUtay2pCp8ZOq2ple4eaNFgW
Pza1lzee1R9bRxZydYWKBtg82DWyVJt0VOX4dTnIFYGXQFciYEbxr1Xq4DOkbC+7Q/JF8h1QQnmr
OSEeVYXIfkk+NL9CwKt5zjTjWMR5B76xYav7FS7M3JC1UI1ts9+WInim8Mq36Qz8lmpgv9jEXECz
9RHE1VXbWbMtltbFLlrjo9bHwnDQTUvqZG01x3mqp7IGZd5CWpvmjGVnPTg09Gj3+w0zl8BH8Z9e
aFQhEVJ9F2tUIKnW20UIJQQcv6zBQUKUpAugecfArWvepr8bvlBDMkexJ96QMrIuUjarCowJkpv1
zF21Np6BWt4Yki4pJ13kqBhvr6tIGiWVCIf9hWQ234no48RU5j4u9IarPkZyscJK0yJcnS0hclGi
Euz8uUIE7Xd4mJUGZmF4irSTCvpw+Hty2iJRR/KZ5STzempil7zM6blp5/y6fJxCM2/AFS+yrpFf
UxOd9aN2VWBWxM6gceEwb/te/mksp80IWXLMrcKjOj5HlHe7oCg1fraRJpillcnth82UJBvowkVo
YYhH+1XQtxfOKNo0paOm2QV7GG25zgAspUWEDnPM3hPLuPynk/9kkM+p39pMtNnQ7vCSvs1VpqqC
jGh9+x/R0NCxhXR734TU962fvgDEmH+1ZKpu6xI5NuE3E5bnVjjj0h+WKjlg4/IKbqiHz6cObQND
ktIsfYpC3EeyeL3yMPpffJiU+ulruD9aos6aZxqrES9xLasS0KYrLemofFyB0G5vkF72jXerwfec
Nq4G9Fw5OafB5p2dgAQ4Y7+TnhmwprEzXi1xkKlxBjsudiOEW+G5gkkuwqUrBngeTvdLj5JkAP65
oAJxgRTZQCMiJ+jsz/lNWtsSNhzpRXMEHRXTGPo4iEMv6jejt5xCMAooUw839HQqzCO2XqPmLvJs
imyehFt6c/3ki+UdDpJLlw1wk7bEsip3KyHHPkCL8rpzWRPIiqymvY1aBKwaQrSUmGxwqyPUui8h
p/pO7/CM4lGrKuM2SLPwtx0ou5r5JCAtkYRmAm2QacajZRSf5fw+DD+SoQUxo+ciLNDHQMhFrKuI
b8bEzeHxX7uQwln7jWURnxWpLAMNfZuLBi1lnwfiuTuuH1cIj/7bIA/Cx2n7KsVA9i787r87ZqF5
z80lCBgYklDyU6GapSCDTP9sreAyS2w4E8kemASZwzl1xPOLaBHvkVTpSift8L1MorgKqFr1etN2
H9QZ+RLhSD7PmmTYmDHWPbzCmSJ7a0oDTJhdOjxjK7eARSR2Uu0vnX8wfwk9LSjC38G8RNdFyTG4
EYgc0sgJnPegpReb3ZUvF0qDTajzc6bbl31mNAK7NoYCoV28CEKTTXr3ChK2ASPvh3TgiKABSyu1
fvi72lYL3I8cFyon9sLTr9ozG21g08UZsvqIIttaRbMPKwbhm8zetTnfbWYvks5OdWkaA7NMx1CJ
0YwjTORb3TCnCfs9w+G+7CIlte7jYH6ccA4K1oC+mrPz8UVHeisKtGAYxL/AfS3tVGhvUKCmO6Ie
/rYIvr0AqDMaCiPLFoLWjqCrsqn7Sid7mkMG4a/9Gx0f9WMuZSgfEDMEtLssYX6KKKXV30Zf8hZz
DBBlvkuTooOikcI66YvL/iRAt2OQvVsQzG8V9AjKLirQRgY0easgQeshAn66a42bbmKZrgfaoC5J
pgMHldXavn2QQ6TbPx05h5HVNVBkZw1ACQOYPsJyiKsuzxGE2p9nJVK+4d+7mwcHoxHULmOw6GLm
Dlx4cvmdIDugcPq38jlJRSv4yEY/HIrXWx0VLChXZO+/n2rqkw/k3TsUOj7kjeM3N9FxuEuO2c/e
g3tiIr9YK57TY6pnAWNGkWQDbM+YdqA4SvH6iGaevZEfqW5ElZg+6scQ3A1f+9FIyvpisxaBIwNG
mdUMc+569P6kBTMXIMEarrVO0w6qwd/MK+NkwfezRHu8P+lI9c74kerPcV/9m4HcDZWECe72xCif
m4DojD9fFn6QFyfMXeP6agQQE+DFvVFyHwDXZFv9+2O64ShED27tklm3e97eypPKVPBedLlwIcAa
yVC7hE+5fwED1OZZKIPbaE371isrrLUreIh+XIwG0MF0oc0JnOtd+UNQPC8SUzI9qE3fESrppOHk
eiTaTAvG7S7SWoyubUhMSGqPROD/koeUKFmsurG49aiTArWubkeLfPivOKiKPn5XeOXOSf64UPuD
nkuOcLYlphGPWcxFeA1Mu3dqbChtDetvTTDI4Z6LQWEX0wfhq0BbmgIxpnlsQzABZ6gmQorGLRhG
fUnAFAoItjrWxRKlG8tZj85FvBcohFDfAdMj/vqd0e/9CByTISHavfBJpnMM1Cva4epSpGrvRWfo
pKBcj1WAYbCad+58LUCtTenZTJZ9zeMKvDgKJsEtWoqzFt0pv9C0iIIarap6MkUP+fG/Ln8ZAx+Z
ySG5bQqZ5wLKELV4IggLmXRlOdYVPpqsHV3EHFMuK6X2QhTzbI07dbZwEjHdTJjDh7y/Bh5DvZFB
rliFRlDwfulDVS/AsYUUQWTo9B0fqEjwzPY7K5fWufEWsxRji+JEV0OyBskhd0tlmvlSNwJLYgh2
TQ8hw2Yi/mGL7Dm6xyTo1hTyBi15k0Qa40CBrFymP4gCRqt1mJ/g8o1wdBMNPFphDpg1wCOvEMA2
GY0cgxeQ2mtVHTmvPYxS1Rk1z5IB3vP+uI9tanIdPyn3dTbo6z7hb0vZnyU45oHfSpsBX/UjwyO2
vm8F3/eL08IrMSzgC97rhGunM73cG4rM+nfKdCF3zxIQ5TcHdh6wlgFvzfWprVQqxLv2sQFKbo9E
2n+yOuDoQGCYIftKpgtfRW+lY4kbt3jqxy4XuUMSrKVYTS5kjFZZtvkRP0nGOwgp+F45tLJ+GvdM
tJA+ISV/SOLEaPuaKDVFp/RaZ8Pt2pXnLVDYHgNmhj1eC3nmFaSGvAYr7EPE/Wz8gYS1Yxky9QzM
QlB7NQy9sx3CraU5hkbrjnWf29gbc8eZVl4OAKV3x3P8bJz7ny6UZXJnpN7BEN/UR/nXAGk9azQq
1/Xb4COv4MaHRdhSudGCa/GuyIWHG5Rp2riLTWNUJv+dmogYCbSQ6B2GFFx9H1juBsUbpUp6xZVn
wRQpirb+r73P1KN+8v1wZhvDGL/H6MDKbI7UDjC3jBhHQJ+c8sBo9jof8nBEqrGNKz+WFoYyGv/4
jv4mdVmKnTJD3IxqKq8fDOzZ9H2ozMef5Z49m31jHcYkKlHwbdZSmtm9o5sxaMeqSCy6naWb16G7
T/yobL4WpmZfMrcNnFoJeuT0m95qxmss1PHYLAT3Tu8tPNq8oObIkYnsRaxiByfA6CzPLPa7YM7q
Br3XWD/wP395Kvf4lLvG+BawdphgFjpeiWdutREueYZ807G+ektyqcAxxkC/1t4I6RLk1PPNIPIR
fL5oX0r7F5doVirgaoWVY5zXSWiwgDz21CxeIeCc0Vz/NJeaqkgFwdsr5QVDgoNPb16fLkTLaaTf
bCAOTV7PYbhWKLNPad8gAF/kjKR7a8BS7iZnZDx2pUWikQpuF/Mltmbod/a0vRGk2nl563UbhfLz
D7VGFkmVLiX0SQLVQEWxaB0mjGzbKDVJYnfScGjCLKJxeWOHb28b9UjRYrEc7OxvP99xYne6h4J5
UGdr/ydMwyLkcKezjBV63j4+I9dJOEMzRTef3JOvdYTwqrz1Xf1QBuT9tLJvIToZIjMw0mKECWPK
JK7zWa/Soy7v8ipHcQHL/VsCZeNZTaxBbBK2HJPtMFvSVk854IqnKWMoDEpKcQGyJCtBIvtTsti8
4ubfuW37fRHlxqkHFQnbw1AoMcfKLiaumHWg2N+WzOGEM4MDezSejSKUYIHbimLHs6lxjFdgXdYj
4PcjzL1tPfWrit6Vc6ieImDHRtHe1oRwVvPDLYl4mxAkv5TGloSuUY0NoDT4iMl3yblrKOVTgEUP
iq/Qu20sNgb8h5GzKJ8dEFfoKaXT8MIxCJfs3VZ3/LvUYMvv28pIG5fpqA0/yhN+An7JvBSyzkFv
SqtO7nB9Unv3nLi9x7TeMMMCMqpbPsh8TqtGyZTLGs8PqF64e9A48jADaYDnsVkbxVW1EYWPFxQq
W84T/Ft+wmYuhJ+ZKv74XMZKrO8So2W6eb6WC6zaSLCQoW/7nmBx9KmDo4rvvdUDnaJhu0ytNskz
pBst1gau8M18Wq7eXv1I2NK6/GSSFEK/sVKx0UNPMhpjD3gmV+9kc8t9XiT9Fsl09KIzqovRYROt
uvupwQSTpCxQ6ETD24C8f1ujNWVCWyax/mZwNK0mN8SqWQBvgdibzAixR6kUwMQCc80SpgaQSAer
eH/3K6C6/0xCfp/lZiwdlHiVtSGldw2bjVb1p18EnmXW5phOeV0Plcoax/b/ihx/EFYkFppX7Uw7
NdvNYtmqsOY20aVVnjLxaNeGMwvQ4uymeVFRo+HdN8zdmpiuFnmR8qFn2JB3GGKyGKSDlHDFe/rM
9ctPhcImp/agGYUH2tAlQrQoHuxSNDHueeRr7hBtCDFMtsWJJS5p3rgrpkv0amE3t6KrkrSjtMSh
psw2ECbujs8UBoW5rybCXKV+cUSEJhhboA5QQm8ep4RdM0I/IIu8z0zwvK30YEmjc+BGVuGspAxx
aPMvmtZuv6M7kLp3w6kwzlLP0FgJCAD2BegsCKDltt8ACei3+G5pnPnjV2cP18chlGVvaS0mfg98
mzF8i2ruWT91uXo+2awOtWEIIDVGUEiu/Lq1rOGrr+sRayTLVcxw/R2ovNhWCN9KruH1vuFC6OgG
lFQpdRlCFkxt+js5eq4VDM+mrPNQwdirugl11dBqrn43dUl5Qb+gMBveorPn2P8nMjd0wwd/uE22
iZwH2Sb71YKFvNvQ1CdI/hfGI+ksSH/iVjE6OjDIAXAkhVIPXQT2UqU9zueuEVtq6hBaqDLG+j50
wEUY1/Tm17EZs6hh4dYHdm4RlWLp2tgG0l2/RV9ffFAnVUY8rppBcjvgJxob8UqTDW6Y9Z07hWgZ
5/Ad21NqjwSTxoEiu5jGdttctIynGTe31gO7FgBv0HHJ3QjHNwOtZ6CmxChJFkqeD5RxuF0VqVe2
m+5nhL1yJymwIvhnJvbAki1F8VtqPE13T1qjEfzGM0LtCL33XXUtdgXdRHDUQ3dh4sDFOFHpOgkU
4ZQtO3JNR/tvaCSzacfPdD1HWwEqBlPnLHBr/MxegTrW6I4A+Co0YWZXe4ZA4hYlyYpU7abxHp7e
FGAtBnj2yutkmF6ZW7hEOUYUU564hq+u9qWYtGnBQY3f255CHgMkpmTawhJ13UFCZ8UcgkAXCeJb
JOT1TSnAPTKotIZ2Z2joBGrXIB41GZwQEAYRagwGIPBV3BHqvwOitTgxeCp+usBdUkfVKLdHhvlX
58WTrxStwU2rZfjE+UOZlhfyCS64x/U703IPd3OCC+EZwor+v/RF7iICmjIUqH38kbrZCC/docXD
t0Wlvz/dXF/BIfP0qq8UUtwP+jrQX7IUCcxjefvJ4vKbF7/mTwgqj7qZ+tpE+SSFgpG3pXtSED/6
au0RIVy/ZCZuqbMiIMM9Q6Gw30hFqejOrYg7rg8jLBeMQ1fZ/w1IZvf8kzX9tov1wGKVeBjlWLhz
2IFuVRFOPx76S1Xh03bDcCDTn+qVkaWlQIDzxBDEmcBWaqFqERtGPlyPxrtL/0LCFwu7anAOLzjO
mVpo0Y4NaUacMJ696GldIxqMnyh6zhW9E/okE0gU7cOsmaX/mxPMXXqhliECh2SQsHHncGVfj3NH
9dEXA9nne1gtIgtFvx2luWC6FNfhadwmymm1Ku1NXNvD9DVYokKzXiEGWv9FP6psmOF4vqKUDgKa
eo+wQ45qqKMG2TBFDDzMKJAqS6ZTa1+OLCVkKTkRVd97kyz9HdBzzrFvv20V42ZzGQGdydKKwBmN
XBl5zx6hn9RE5FgZWbRZUWMrZEwG/DbEGSF38vfHDv63lCSR2qYDkxAHHSAARpdtHW0nqHv6aAnR
4izKI3LBw1G6uXz5qI34x2iv7gpKiBp5YodSCZCe5o37uF6pIejS/9KAODTbDOAubvsSp1RUtS5E
XJOYzC98CypVcqcoXIth7WrVHMhvembkv116jxnkNeJoHYu9KlbNWWAd1GKhrzzakuq2gJZ/ZfKy
yOVAknORW2xyPXgHS2wlC2xyI0G2eF7+6YijN38EmtzMQr0Vqo8WMeUc5+RHXnhKA51VeSY6od6h
chZHKSW6IrqJITn1Q/1iDxKh3wJXTOJQ/k292g7vsD4pBLE0sPXuoPdcQPJhUxsEu5t+fsPOp/ba
y3Sq3y8f5H45vBbOZVsxycvlofqYcN8/oUfco9bAAdzDxBJ+zqKI/B0rWAGHMMKxbHmHgDec2gGf
sK185bpYbZ6kGVVNDGsjZRpQy6brMBEVZVU0fp2CCeLglq+fQ1p8VtxYrcO3E+XeeKxe8ngBUSPv
75MqYEM9Goh82ZpuPQ+ySo762svIx70z/0NNqUkgUWITQxGDY66Qixyry9RpYvvaNWM899/JoC1L
jNvxeYQyyzHq4JRJKAbp71AUu6Cdne0ZNWhN3M16c9wzcD/2JlTkdmzKPAU6mDeLirmKVpwiNp8h
v4HE1wKeUzExCJjmHq9vuRW21sqmlDSWUykC7QRTM6GMbfvLxwLi5sZ5fM8u6EfkknRVrKImbmXk
/zU7DPcmSGp2MUrPmOgy9KJ1bA9jYZS1ioz427lsRQmb+AoUE3BgNy8OdqzsgTb4vQNozntxtKJY
XzYkUBjzOtSkMIo0ftouZLvyJXL9a2yzj65nn+2tc/1ZYjYGRqhRNGyYn6xP9UJd1WIDYAVtk2tE
tJMch0QR3ZGMwdmYDDYB1byOwidXS4+WYYxRr5tmpyrYqwGEi/A8qYf8O2bNKOkdXzT8ICiss2Vg
AztYkltgtVdUvnCxaRPC2+upRU364nxuVhn/dfrEklCol1y1Lq6wU2calv+ZSxFLhqJtv4sAcwEk
KuUdvnvlEU3JfLb+oRt7SEClFhzuELhr9IL7HneSKBvZ9dlEpi+zbpIP8L/z8KP55hvKVUpZ2otS
SS3KJSZqiN5qq8aLllSWF4BYA9ylV0JZSEDnr+vjXfJSnlmyhUGZL1apGILYeXMBTmH+aZYmgZTB
8tfq8QACTVX0BvrW0etX3sRc0v5OTAj1TWIBWxuq4DEc+15YpoCniylAKiHvzt6aW8/sQNJfhMmx
bl1J4FwXxsXUJXwUCZIuIVuRFFcOUYIVAPt6Gs9f5xYHITDc6SVpOv5jMGnScfz94vXeBNkJ8uG6
0pvbvn+5HTUzQkEgPeca/0UEIYOU/B3qfGywGPybDzBoXYZw4iU9BhTNW7skit5TQk/q2ZIUF6Q3
yRj1k+MW+opna1Wsj06vauxhoa9HMzi1iPvclFF/70K1rzCIRdg9Yu1X31O7yliEKNdEhoaIOU28
hlIR9KP/oJZO8OfkTfNZNZX5S8IyFVz8y0cpZwu1uct9h8QwzuLo3Yqaq6IlMAUs20+Lsj0QXhpk
3x7gZS4DU+6qpGINH8mtqF5I4RprF6FpBVDC9Grt0895FfKpeAEKaopjTmni55mX5n1RU4h32mN6
kYrwU0uyP8FiA331StzbRIMBkbisv2nILG5rzYbsXnA6EYVb5L/y21m/8I+kQeZHPE7bExWERRIQ
7+TayJ3zh399KR8EJoQ6Uh3q+hhHVEOy95IR8vycSP84voFgJUm7JfWV2RaYsfLLh+RweIeXYq+G
ehZcgsR8D8UiV7KopCxxD4gdCkuVfi0eYLm5vns1pJCsyg5SkMJd1z22Ry4yus63pk27+0Gv/okb
r2a1EoOJrsaaf8ZRgxyEJOFvmJFMbu6H32iQuY16jokEEHDhenEi5Oyafi8wKQLAZlRbEIjz9bhF
+pS+gUhYBvZ3FpFWIPDBR7JLzCkTL+qoTly8/p8HM/49AMRvnN19fkOEk9OuRTCjdcsgLCcZaUrt
ZftK5PcyesmCadpErSCR8r2zSMGkW9ADBJ5jNmqtHj7TM9QLWWVJiBye53BaMMeffaDiCXWw4Q8G
rdPkj8BdDVSJEcIYR8QotWKKTUDlb3Vymj1Di3z9DeOMZV2AM9t5ms8QeDXS9Ljt5PCWqaZP5whR
I5UQK0FelG3reTAmDDQldTul34QewXryIHQiwrKKO1PQb1ET3NZC2tVsnMfTsGlXmCaWyyzBfapI
RW+vtt1PvvrkrOikXo1TpASa9cRh1kYjbC2WuoUc8I4wfoxZ+WUeQ1Zhp4pJ/JpXrnkyjtAorf7n
82errHZeQpicFjmqH++Cn3J8U06RULhJqHzGVVr1y/VMXWAzIFGvFhR8quNtu8X5SMDGorfBndeF
oUxBPqSXUc0lWxzxkg94UHDW5pr2xHSbHeLECcEXCt0SA2NWU2aLBYZ/KQJSGq6P1yAIIolrp6R6
3fOru9OTC/XOvAs86vpChbSyLjs2H1lm3tFqzeCadt28hHPo/Ifq0HcrGmEUCGZ17bvHMBF3sfyO
07bRtQDcK7vCO9pl84bY3o+N9DmAao0sbcz0K7HAXo5EcOhXgn7cXI8X44ZT7uzbQdZDr5j5C33f
Hy65754n4THpdZW8D+2QATJjbGL0uzqlsGHJ5KhnGssjLspijtMHJPw266rN6k8YWB+T0O7+HPNu
ClL1xCpHQzbEdD/4SSS16JJrKTbpqMT/ErJ8nH1AUAesinK0BGloxGzywoqdO/O6mf+hvcA2nHzh
M3IcgokVROgipUEslNvPEL+jsIKQcF1CtU+rNcM9HuTP/o9x7VSBYx9Rua2dAavzfxgR9AT2Y+z3
cZyx7R8xxChNxcvnaE8PwFleRwwQYLP9wkUaPbWYbMr3xLW6Ux4hhq/S4IOYi/adn/ytuqD/LYse
2Gn+f9/Q+oNq/x8lvk68xKVwRWtJXyqA6hsyMW0/Q+2hIikJUuJWSrDyVh/rEPPw6Jk1uOyxDDum
zy2jweHNiPtXwxlSTztLU6z/oS+DDBy4e6HfZIs7aGNt7B3piV1p9NPj7ixNL1frVAuvFuW1FtpU
CjXBRLZkGe0Kh9nQSww1tVzrrTJgiCSnT4NZJZdj+Jhj5oL+89wb82iOTsJROE96kizjeH1lcEhD
d4JTeMtYh/zXai9KKRdrn8qe7sRrUihvxA9u8nuPQTGCsdnqQcCxX9OCTWNGI9sKzF1USjEoCaZe
qSQMC05BNcfqwXh3mmIwyQCIA2Ni5acmpQnMba90L5wOQG/7Pc09epBRmIrTHkMGAS8BLqs+9OdL
DrRKLyCmuOMnlczvSyDomOBIJcoyb9B0ZYgXgpP3C5sP+vse+Cg1/m6rb6UAQw8SEySR6CZ8cIGR
FMxkZByy65GO3iQqScVdgeG9Xz1puYc5p6kkKYosQ236hVgzP4H2mwf7kX/sMHBO48c8YdGx5Im6
OqSGk1ltN6+c3fFHxAc+U6IXGwXePbbiv3IbE0hq/IHJDlpmFeaWB5udjeE/77qhDzIluIudvsl4
GplkhXUHepY4ybt11wCo0PjOuZ1GQsbWl9W+NLi+AF8wi69b9r8kQYRhgnYVghfvcjyj4QnajNYA
Ng5vNbMWctzZMGFmhP2FJsadnaPO45CE2ETBxhKTHBW+lTh1gmgKMbDhHPrLjF8zj3wYoGWjNaZL
1eLYewtnoK9W/1c5YxjNX9JqDPfSNFcdKtKwQWk2J4f8BFOP3RnEBQjFSDWY+Ha9yXsGe+YByQvQ
uFzWWeTs1DMXhyVarKOUPPxAVgX1oSwZEKl9KMF7N+fgLGE1hXolP8Zx+sWThQOKXk6sKwA643tY
RfA1s7p9C3EnAkFk4nV7nI99jIzcEjaPfNUq//XB1OuLtOCdDA2ftb4V68/IsBE/RwluK11cEhTM
lrlPqzy5XxQT6ASKeiD08JWWo61bxvIhaPezRnlB5ZEOaf/uqp9B0QRUa4mzuaGRkDjjh97gxZLE
Adal6a8GzZUPNKDxuEwOZO/fJwOUYEKq9GkNOXK/9IjFxN9GoSyg+3aBVX4JdtbQ9qbBGOS9tTaV
CeKhohh2oUV649aW4pIM4/C5jLLPBwHgQ10M5oYXqlgmYbmJOtRehVGOkYvg2NjFNMX/1tKgKMHI
cbo+mOOHgRsDH4tugkJIJFzMytM9B6ocC2cdSIomMZZKptRyfGsD8c1LXaXP2DvTBnSBUjplqlUF
yaZXuQUvwbGu2Cu+AfJ8rQGC5AtXmIWo8/eyTTKrels3icXLBBrmHYUQFccodrApuDVqU2PbDni9
XJZayUI2fR4xzZJbW7dxh4muOINmvEC3foA4cCvTxFPQMxSfFMKcGUNFz9iIRD5f/MUU87Z4ycJQ
K+/wa+WfZ7+CNWpo1l55Li4Jptg3FQs6WT+t/BkPre5XeJdV3QN4VsjJ45Fh/JuedsJO3JRFhq0r
fTyhF+qRitnqAMAm4NTjqd8eah1CFROTsFXEgpPs48lGRspN7y6rISHdhyPb6l9z6DPMrvEt8Ncd
HrinPrxwIHvHQwJmgnPFZouX+2CEafi1hxVY9hwbyxiio4P1EPP4ey2LvQE444y3Yl1idhWjYjMh
m9aVapQaaBgneMYMBiK/Q0pVL9FdDwV3ogmCLiqsG1UBOltsLV/HmZn6FVdUT8uFHLCQkwxJOwbG
XF+5Qch5P3V0ayUuLFKGbwRdtmoKDkniSXHMWtpip29SfSmWmUqdMWbesizYpS+oshDvNpI3a7tB
igT4qLfVi3ctygwa9ERyyrQma3XcVaEOWQcCsf+8CcEYdThTzSWYUTJK9A1rPWIE2Id9EtCahJxh
sk8n5rGW3W2YZsUSHqqqWeiwZoRSoN6q2MVk0Qr8Efy1nPXakrlePVGgCsv/f+mdhwFkPHW42JvG
nSV5mjK2I6gUn5V2GxginGbdFXh8e+kdXMUcsfiuq4NEytlb9FTgTOMg6NBY73vei1JvSVBzV10A
G55AC3qzfikBZwQKg/IT8PDU+nMAc18t6hOVSUhkQApH8yVddS0EVeDSLySEvqjLUe/Zg8t9X+8q
6UhFCRLR/lbkl43yex3himcJSvoQIFeFmk/jT744tAvwMXObsKCKImbVRWMs1EECXPEyDfVyY5oS
Hn1YdqGIIuHv2ducl+tqS6CFCYDEmEDfqzDsLrfKfSVBuFFv7T1W0rotZinaFemjqn/mVaGbsG1W
hYpzwGLaqPdNZTDwQD0Nke9B53d1iFRL54vJiiwPXXhZzf0C+OL+023se/DDtaSSY55KSrW/rOFB
vbROOnKDCv1hDfl7yU4rd7CysLmwCAiLV1wOlw+ZXpUlKa5YT4A13Oq1fra51yIB+5TRhFOWcAKP
EnrVdY37yPmxM3pBroa4GinBtVjbErOSmvKm0Hd+POgZYr9qaX+6azA74mDlXGbwY0IAsyJ8AwH+
AnVb5olDsX3JBLJRkzOwm4jRyQLpX+kk5oXYH1hw8X7Xm16z0Nm/CRAT6IRNpdRF7758cqPpVdf6
GUthZUTfsQOpRqI6k3bYmwBiZ+dcyBMo3qC7dnVCw7hcWkaSUH2Sc6vxTsBNkasaxkPg/LkkTspD
oi55lFTmdZaSrPTckboCV0u0F6tB88zJH+EYESD1TMQfHvEJUgsRRU9MPfAei+77sPhqyF45sZxn
VYeyKyNb+hIZiV6Ttq7j2+UAElVwicJAjqATWeaeo+otrStNlTdMbUuUOZOQQz8ngf34Jabxbi+s
RFAgn4yZfSrdBQJu3a3qFkuv3UY3ldGU5iADflXm9NMmXyKZNmKceaMin274tyquL18lrW4MLdED
DtCqcFplS7pQ0SgdVSVgNIQg26cBft91N7DVoBNJ75RtTLxCPpBb2G7snElv136KM5x3gPVHxiCY
FxTs/mCZcNLeyE8+LBkEcKEv2M11k14iCiHbFZbR6kfN2KSPN9UsIioO3ue+fD5q/BSgugvYLtj+
1kDPON38nVOqckwqrY2rd/wkZJlXh0rx49Tw/Q74iZTEUEU+nFQM2fpWjr+Z9ROg9GFhdtjAhcYk
TvoZ3pCPOplKkOGG2g4r1XdmzVFAZLBtlgm0dDfZt6/2XcY4PVMp5HxXnop1f6ML3WCRLbEemPlm
OsBe039VAENGGn4eS1oegKvClsY9zjBszIVvb/t6T3PusvJbAmqQB/t0NtwXYL280IybQWbb19No
kAnUVemsKrPBQjoqAywZzOi3ygH7STM+RGVUlyQW73OO18W7Nupr4g5DI/iGZ72bfF3/JpfuPuAi
nUqZNktKvIJHwTiJ2NYhB1B8Sm4jMZgiuXd1HRf9d6re/CcGGdOKmWkkW6l15vOcgjYivctULFgW
8FqF0DdABv3imiXz9eiyK3DZtqTXKmN9yaeNbdBlqKJa2UntOLCX8s6xLzltzhG5RVGATHITR1Ii
/zs+c6eA5VEQKNB+0SquZUyGAcHRZBWk4xXFDZkBhpkfTjJ7wkg9hRcC9or0AfjbHhM32Csdjwga
YLdXwrv9jpG8e4aGIQZYmZ6gaRLgSOHTTfJ6NKlbANgAquUVswsw1WRwHNsJlKwNmfhMAx4Gm7wL
gB/fIBy3tFD3ehInc7XIrDydqFFzecRc/u5LOE74iu3c0j1CbWZxQ/LlFeexDAV985EFwSWxaFBb
MJH/jB6G8j1xXV1Lxq3BAXs5sfe3ZMlwicuKL+ruJzT3tovHUfwtfkWyk4vn8PMKa/hvfj8wPHif
3BFnxoaOSABXrZHczJmcQoyZQ+REf7nWqr/hhdQQJ5KtzVcdVBNnx5SC1DlfUVPMPQROlXrmTvq1
uyI7NgIWR47DxJIJTDCvgylVbuaCacfZc1mhL9MD3/Lr0IcxkMuVPV9Opcto2wRL4IGcN3QQ6Hyc
pXR0SQjfhkbLYoIns9f/1q6FnJS6g9kRebCmBHRP4ZkQfQfYocMmeG/gU2G/c9f3RhAyZs+IlaeY
456VVaSw2MHhAiI3voSxj3Ezfh40CjQIIMPF0hmBh4vRYMNlEVUyLNVaV+I1EuGiL9sMFOeKuWYg
8e3iuLHOCFR9CqbZAOatep5BiImiqJAx7n4gE6psKpIY63kwNXnjPZGdE7V/iJdz8Ia/0b4+pJIv
6PEVV7bEWHehK1kQfpxP8Kw3ySj1t//z/lBNjysEAm2w8pWmRoMwy1aCowACspW15fQcjqTDso63
EMqOclu0x4qRLcv23tUbg5U09RoM7ocV+FhhpB9PQCLEslo8YU1WykTobyddR+psJ8o/9xrccHhU
/gqyufrwhKRXlxoWKU75qJloLtbV/AbV7GWtz6Bz8nHj57qlrESPU0V5ZbOQVaEn5nZC3AZhMKes
jgP8a3BSeapu5T60m5rqMOICFI3wtwtoEenJ0S98HJWjKimAXo3nrx78/WCqrev87LIACYXQKs22
o4UEuCPRL3HWGAgBacpIsezV0bomZxPUge/rfFQpeVYWFTeGvoV0fnJf5VkFZ7UDgN6hWdgIdZHS
ep6wQ5YfAm5acxLqv+fCDd52C0tZejx/ctlHiHhElBJuFbr1YAe10nl2DxTy4+cbnPqPq6S3Eo5r
LbiWJX5ohqWFSH2FKYVYrHKVKCA9gj2WEEThOHcBHJsToOlj43w+mabdDButlWix7x+2koefKKSF
OcRnNAP3wpFatv/9qL1SAeJ7NUtyHH3zKQpANB16271PxjUXxe7lAwPE4QP6qMxaUVvAguFbH575
ZNkPR4SAAKsQymhhs1W5DW8TsIO6AmLnMnR634tsCxoIwOloO1Ih5E5FdTy1lDEar/KoWCvVEQZQ
bniHN1bsXuF6L/Z+IuGpySIEot1+RRIhiNzhu3nUPn+WQ5gkYsqebRDy5bxBZ9dJgikQ6XTeggI2
R1MO5NqF0k8PEYdKSpL90fafkFop0/2jrhkzo4m2gqRdSVpjIXuh07sjXtfQMCQg/iWP2X3OYZPk
Qm7XNMB9OuEBkYty0Mp8JAUDiWqmio/p3+eVDndeSKziLHMiDBlSn0P/4XbDP1bmEmivZXhoGR3N
t5MWeC6KV/JT/yhzsggVQVuzh52ETpWqx18S2RoFivumPthBsvQYmNbQlP1T9iW3vS1HrKkX+RXx
+cRPSnX2AofsTnNijpKW6l59yzSXcHuWrx98zLCcrbqAK5b9tIIUKKpi4C1ofbf0W4iSUYnCEQ1f
HFdEqUwZSgY218/cclmNHKpDfS32By8mf6OeR2UZ1duLNzDYPGi6b5J48+xPlbkYhWzDkACWPr4i
rwAfWAnXxCKiYwwdemUqjI4vAPnXTsHfgvmp/7KozKgCIthLIrurWywGa5/EUMGt/L5Cuqu1fpFn
9874PdJPvo8FokqwYgNnqarpqE6HVk0HP5ZeBNb/VkDrzOpWD0Llxf9E0SLW0IeNGicoyNPCptwN
kdQgx9gtSRsswiZNErJk+agGSSYwSDy91Nt3/7U3NXQyWvV2G34DrvznbmDm4iolR9BydAGpXMg8
g7RbSIUK8mU1vmGL11Cuda7J4rslblULn1V41hZAPhMZiQfnxcLzF/y6qOyX49E5VWvjf92fEpot
FZmi24YTtxXrvWPcNMiQE+sWJsc0lIybiFt+i5dCQGcxXcV1YnBT6WRko4A0qGQ+cotA+jDuoQBG
Dzv5fz7vmCtbQoe7UcF4T3ohmLYcdr1cFP6zeDdXaISsYKp55SoMDy2vo50u18w8puvpMiqRzFIu
UuMOrSgWetgPm4B7pGbEaGpD1eARb/bok+R5/gemcBgi7sfPxA+o6/UDIQM2Tq5iX8g3e36R5toB
7UY/kKtuAkuKyVASoxSMscqTqBihwUaEkuw3rGYfaJPAuZtIqQH6Orw1bgvjb0SJ1SOvAsO2C6s5
wCTkY5ZKYExxPi79L93JmBabAK1BaUotZdRM04759JRFUDMDVLSAlbFpijV1o0rricJrT9DPA6Qz
7k7xyFZ0l54+XeZhcFrfOkt5NizroJM1/UNye8eptq7DNxIVtgoAZwQwG82OeW6sZ6foebh4v1Fg
kwrvPBK4Ib2mYyDEyUf0S4wzusXcXGssjHYpPkiJPxy4W7npK+YhqCnbc9dVmxb1IRvzqkyRGsID
QJhhfpUnZysUXSW3dJmdHX7X+Xx7yPCOdYsI39XyWe10WCc3afYpYwZxlTEzqgG93SUFJ9ge5MwC
Sz+srhROQypcUwUmmR3U8pxpfJh6Ds7p1nFYJ/7X+39tnEI2RrIbaEAVkcLYL6GfHczom1+WnJGl
OaL26Gu/YXhXxBq4NLCixxEOfbDVs2HHQzBd9vkzcKW/VQxc1fOKt2u0iHh1hGqYRX+gf6eSM4ho
rIqG2rMLccfq+LCEF0Ayr4UO29liMiuxU6WCVR5qa41+qJXRfw2Im8saCuP26l9yTLVCztBmHkZG
vRpnDDMESEAXLllb8BV0CRA5ykr10FBf9KC0DQ/RmQ4YNC5ZLAMuYE5lV7Kyb+eakMPps8JnKl7Y
P5m1bBXkQxCABZn9aR4lmhhw1YMgHgo5jXLLd23jai8Mh4cTo8LvFgyxNZlLDAKD8wbTb+b451d1
VRcwiYL5xtzFPmXTdE9olGUrnkcOjAUAksJgra28yeFP/1HLptj7St7zCPsN7bRbKKAyl6UFBOph
txzs2ZjJYMFB98LoX1T6qKJbSEy7Hz7zwcljpydM5EJHLlC1N8WQEtS2IvoBMP/qDuOwia32vyGz
5FwQ16lBLdbj/3AgFfE40jFeL01YV0OwZ8XqDUUvcVAGe5Q97AWl5rRriD5Nf5j6Faw3Khl8BUsZ
Tb/yDj+aUJwApn0ov0ozhPvnElb211loWi8rLskXKETE0CMhoMhkhOGlEQDZQwP6a7vcrcB6OKDx
+YNqZhNFdq7U820A9JMTZmWeJQDScdG7UarlygJSK6DVOZreiSiB4IxvNnQ1gUO7O+VAV1xiUkqH
Ov5EwyrkfesXm04Rk6OcfZV691fnY0qHRWnAcay4Ojl5nKzHTMkA/lNM0VRTjbM9g04m0CyQb0k4
r0XFpZ9uc+m+PUnWqrydY6YeL8pqS+oKdAsvoa7V6BHXO/nndgkfa7peNhlzMVSdDbCoTs32o+cK
Kj2th79derFYkW16kNEHGsRgrih94CA/hiDfMjAgOH+X9dZFXl+EBLBalmcQwaoo+EZFlnrBbf1a
OnuRzQy+IXyS8ShkTkIhC/6RkhTodUUZHvpHQcXCf+HAbzpsU4+r/MsVq/tM2Ff3q1mja9gx3vZt
2uRMbZq9vcj3XdH2p5C6eecSGjw40w/gcJNoRkO8UzT1DNBUfLrKZzQ7Tn8TzZsGKUeheqUiPF/B
Mv20ttro50zYl+M3XAaqGSlCJzzJcCP/HyRRAQKPKHs8ViLduReHkml+ZVLI9+Z3IioryT0cVv5f
ICCBrj1I6x+3B1Yrsqr5JxKCRVL6Wq28M8rdysF2s6Z6NByq2l09hp9Hx277dGjcTD/u0hsmZ14o
pZH8mGru80wiPtJYFbuPmVqW4CXpdoeLXJG9rZf1goLhLrFGKOJHrvjcySG7ytWJAPpqMuDYq2ZH
ZwQ5L6GvA7qs6G8yRdWPJRgeMHCy5/4FXFSljz9PICTlDORbY6KV0LZBpRJ+XfhEry2whkT88lIr
njxOxwmnTGatQ494AB0I3zh6DmJxabYebVrggw20K5E9ae/lxkIRfAw1n4N8klwv+QzbWvZBXCy5
pOXoP8vDTSEE0So5IsnrI6QkgYEej1i8qZedh6LVBebYpKMvbEfOFLInKegSEZRtJ43LkQJZ3gj3
wSXY93lhd4RMj7DzmiXIsduTZ3zW4XApBjR2r4jcYNk/o8IfZH6TTFamuDXfpO04e45b+oYwn+cZ
k8GWYyG2Ad6kvNH8IIPSzYqd8ldoj9s4F7PsBM1KSk8hpvqkYp1JqNYZPdXwFmg0cuxujfIj8eDS
3Y4G3nMzx+XYbt36mFGfz6DD7JdMT+TIv2Q3oTK0/yZ7znf8LDSbysB8fCLF352a7bmyZ/RMjYnu
rrZjSGZfuWN+NAba9qjqODy1KPk9KaUKuJx3uYvgtRlAT6MtCk4Y3n2LRUBGJK4HCSoCIM+hhI3y
CB//FiYQMHEEJfpnJY/0RPClrSbz5PGnHYS6hROSAdApAtO2mrf8ew1w1lP8Pk3kgNNIT32jZ4mv
ZTet4MVlRXtn5U3BQDo1xs9ZZLLuXhBgtZJSLSck69XogsGFrLkdf1kzsLpxTv7OjI2v3aC4DuuJ
CcVTOEc8yU3mKidHDy/a1nwGY+8xZcHXgp7DB06kEuW44PY2giK6Yb52Ct2DplaYKj4SEBqskE1w
txIOn0IkWeiUj/lmyWE4su2aM8KLOvP5PYUmlVNow9+D5nN6MalxGDi78USsW/t+DYHp8xCTkfIk
gVXLdy8kN5ODeJ0VeQ4fEy00yiJT1rdShToaSCwi2aZryJ+7g+Y8UfX83JjYmejhhjbZozunSBOR
/2wK81DBd9Y90tvK4HsXh+K8fiowdG/y+rbqFyc1vce+zPa1YVoVWW6s1pS1dagr2KAr8e3ll7F2
64VxTHGVG2gbg99i7dLium7iXFIJaTuM7wKFafZ/F+LOdtJ1n5FhiUIeFaeW0x2My/QW2l5ZulBx
CJQSqcSI5VRjGogR8YuO8qYk3X+ezvmAHRt2CI/CdcC+v/hEYhkybvcKweZoFvNEVbgcV/Ab2XF7
T7xTHrd8hpX24wtoqJF+YIwSVtm1kuAreaGux5S4HNXbqJShDmH32Qqtqehz/6JHosNLRjfwLG2Y
4l7YIEop+5Xwwz3QPgcs9/0ve1Kh9eFSeG1U8J4LAHc8R2XAgDtcVMogFkzU0GAtbCL9XY8fa48x
FxjyjZNUjwGH5UJwKjc7pezOY+DO9v/AnUfd5j3U+zCKkdprjhoL8j1kQa9zoEYG8dRWKrdSFTt/
xrPHuE9q5yo3W3pabR29hp0zNmuxx/mjAnCByMSOzc/hHLe6H2Xyzp8ZhzGBgm6F15afPPqYWnQI
ci5zhszHmky2pulxx7W+SmpdIMMx0Ci1bIsw/P1IL+07bWC69EyepPxvhq3RNTsCcijWXvod3Kpl
mOOSMYXYij1RSB4jRIHNCl97YQidjKP3jzQgRCIi+fr2Ei8Z/U+OnZ/U14lpOTIRjdB11VAefa6C
KK+9+MmMrxxqsWljIRdhgboTYvcfZ1NJ6ats6UtvArMSx5f65m7Fq6dINj+yxyVsCilEuQDHsZPM
cUJlunCqDgVPSwuZM8MCLvheGGzrKU2M4FrR40FEaE9zVKPkvxkXJHgLW/9Sc1yGjb+HP1LRWmrf
nau9H6agC+nK8w+imVZJ84qtCR8qVxEH/2CrlakxztsSf/PxkzPPz3RvZR1CjC84TyafWhEc5zL5
i77v8cnFY7+6wxYnwS2ga0CXON8Ht3yet3OY42zSG5abw+L4IGy/GmYoY4Y6hW9KXYxD0Ar2cRzO
piJu1nUbXqyg2ItFwxjbRbL4wTZrPDPWrBLKL00WuK/2ruP1KgkIbYP1DEfyyYy9uLSQRkjr0/43
1C6CSXZE6cKx/d4mPasziUzdmNE9WnHASlxpPhmGSusnfIIz08m1s64lvT1XPRR5TJG+5FSekf0r
NXQlrVo8AQReDrx0sy3PcYEmpIVfaFFktsN4Whqhvfv1WSPZzDu5YcfnaSZbRmB95+FkPuHUvKjL
+UNqPHljD59xPZQAV6IYHsBRe9m/F+fa1AApIh50XQn3mdm2VAPYqtSHm77CsdsxDjGezEV4DA3g
Lik6bZxJAMyVPjBesX2FUXlelKIsPRq3bMm6ulGpgb4eh4LpteMMZa6IhV+dbtl802RKgORLJ17g
5AwNpBE/iGHjK9FaowEJNu+GAO0Rc5Z7mp0GMbngK2tA8/qiNFxyYQOWd27M2PPI3I6Ow+dHshsN
mc1LkA4izHwb43tpu64/Z1bVRCwtNT94w9xvCO60RvSaIaszT78OF+H7gDZUUjtZxBOdmpGsjB2V
j72g7vSfdIkVsZAMJ3qbA8aswIWDrol6iLk88Cyuq9/m84NLElDj+BS3hN1B7yk4xSUDcChQm0UI
CvvEzwHv7LPjXA9kfE764+om1T1ujRr+PLC5TzdAVb1QLp+AuYW4BibP2YWm/sXLJQrGhFyCigOg
+cY/WX/rkt/AawUKyiRYqzVz+3dAxpnAKKn0ACgNUH5NXuj28MqvtE1Z1psMviYBnRfhi+NvmQ21
5ACSVnECBgEC4qEyvpxJG4b34y9sUx4chKeqvRrFXS85M12kZ9MBeHhp2XsX1knhCnnDX+xmyguo
C1GWI/4Zw2um3yjhC2oUPBJDAXpHq+U1QfoHpMBqUNYW/beyks+tbLxHJqxKIuK5Q2c3NiiBTGGL
EzilkRS62cevznDCYVFEDY3WHwRiRn6BWK/P3mjEOj684A29BXO7noOKaPVbCQkywfi7/kNLUFJv
jOS6PyON1sxPQxD9Zmkdfvb2airxSx9pR1gxkVqeH7DIctD4ppZlEiqCRRp+AtfEiBLN4oJuu3iL
S0yDd83mwdnNrNAQv2WWWbyDP4v6CxSs0MagumfljRgjMkkFE7bZtzOsKF45LtCBtCd4aSP/cxnz
hPvG/E/UyNFT9amCSeC3kny1Am6yZY4hQLBeCk3zmp8ebWxBMyAQtZIH5f6XERK1qW+sLRLO+Oir
ib5iokeuA8YSXOF7BIFKbKUkUGFmxVlgwgOtWzy5dnhBLPS0peAaPE84chANSiydujJlKJaKcyZi
hwKp2kiTp/zsmYCIxHfzrAQh88YIjnVQ7Tkcag/pen67UfzoLCykchEjdULv671r1ApYNJcbiEjY
ArcDJi6oiT+ntX1elCG4pB3VMsCY+XiJtUjFH120aYlmRtOKaZiPcy3ViIzgq3uWCFBLRhfwCsD8
gm72/cY/aPJsTrmgHdQLbwN+OCrIuCIhFHrP4heHed7g9CynLRQ1uCLQtS0hwGspcc+RLchvz3eA
/7JylHeRzoOnUrnF/guiCBZ1ymBHnYx+eFIRC8Op7kuIre5CZQaaaRya2UQvQDHjD4CZytI4ixex
pfqTf5og2QCHkRCckVAmXNAw24xTlY+MNB5JTiiFG7lOhGgwQzD74PSurlI87iwOcyZhuP4eO1no
FUE64p079Xzy/+kaQ9yw0s7XBc7xRzXA0oswyjK2VJtEKvBdg2ldfAa855ui7Xj1oklSpXKPoweU
C5ASIg5+fGBYGYtInCDk45Byp4CAvR/F2gJOWcI2nSgqZLIamZyfAJlVLj9jyfclbnhgYcbxBglo
DZUH6tsmyEzr5M1Ty91stf8MT7uNhweSQNpSZk5h4JHwHVdrZwN+2bX6wogIPKQOzWaLk9xuZYpB
Nk+pIHlhS0KlWW5G5vhxL6OzxO1prvewH+4g2r0Ex/qdTxhKpbS1X5E+VevZfJZTp8RLgIbfnrlX
s9N9pBRs5JsupGsU9RjBcIw9g72HS2fHyvwiONqN18P+hGg/c8Kr6/c8USKw1Zu6aeb6CO+qhnzk
VWyRZCZs4V2txRF6KLrWrZZqhzuUHp7e0THuXqnpuLzTaALP/2W6R8GJIP/Vl3bSgxIXDB/ZiaM0
FcCC/phGPT/eo4MFxh/cCf1P9ZEXc8KpCuRGMuCJLusAVPuh5IfISd7DhXoJgYm6VNHSQSA5L57g
i+vbndJv9LHW4datZctZwtCb8Z0f+FDsfifZT4cwEBvTDgjBPLi2lZZTVLgZJBak3ch8V0uqvGbg
iIM82nKHDy8Ei81CJauqbtssTYAJ/9c9Ki9HK72Ljl6Pp0HmzcGFbY2jelRSf21BmsKy//SoUa5A
g1zPdc2Cor68az0Nm0VPe3XN1vPp8WBqgrNX5+EIvAWsl6fXVd3/Ji7GX9g9ccnw1qcONiWs0Ry/
bnydhyVe/OC2AD8D7vSYr3cxw2yZGjHCqGl6dF1r29yeFMua6hY8TV93Wj4gg6OJpzEGo/gZgGSN
mTFYZQ85saGefbjRpvyvY8QnNkQ+EDBcTnGgaMB23jRK+7VuJTU88MrBf7wZMaBoyfbQFfmbauWV
VyBGFlyM2RGP4WdKzz3cicx7G01KJkREw7cPHAd+LrrlJfnRkisbWbKfc2PA9RUbjet+uYpOLyLh
t4UyhbDt6E1HCY+6+Dtck8SavAFA7K+tG+IbU5PBTyCbGJbthTzQ9zVeG4/Q95lxJKmpDRMMPJBc
4qBs0/KiQuCQCLlFgJwrDgtv/AYn5RF3i4D5FyUHMXYWVLafbKnSlYputRFt/aqCp8gK2uOab6l/
s40RJ2I4Ged7V5i/5Y8k/b1Dm4gdaVf7Uqs8D9vrclKVjrhbyNmYqK5n/JHX0QxCFlYYSEfx6v6l
uwmy56P6Hi/YxJhlQxOj5Q0Q5SSxNwIbS2nH02JKYMYaduTvYZNTTuzo6y38YUD5zpc98RYs60aW
JnHc9wcqD+mS1umUysAmrPWk5N87K0JH67a17eYcm9HE892ZtDDPKQhzApfManASsQkCJTzT3yNi
llimgh1VGCRqIHUdcfDYvCj2Xwpp5Atf7gwR0M2r3nv8bj3iZ8l9uwhfzmQ2+0JxPxfI3nLGjBpP
JsyJJraVdluD6RpIiocZ/cOCw+eoAlqsin2ThUPNiNeD3VDswxJrrKkGox1UTUjBfKU3h9Km698p
Q5VkJb2EYrjSX+StNABrOvn0UoJT9PIhVyS/VPbG2wXIdP3S6GLETEzE3//sl6sOnT6wPmArxBLZ
tZ3pweIUbMART7mAdFCES28K6/xYEe2IUKySDGe20FoxlvrSKj6Boi0Mt84eLBpU0TGMaGl7x7Bo
zODQhOmXtWbarBP2gLNFUKKeTxPNZSlEf0xcV+Pg/9/1AQHg95Eq2n9Jyt95F2axbxn9Y6Orgiz7
XVhYY5TvmS9wef1B+AhEdxaCOktBdN/t0AqrwMdIITqYcaMo/cGKvDcxnzkwHSnxiQsnxWaIXvgz
Y3BYrhtQpTqPC98/GRHGwGsreAoc5OjoI6cMI40rSmluKnCljhyDsaZjkUD6rLX08CvVs6jQ0ztA
eSDcco7isv18aKoqQdiQ7a3MTYghPW0bMiiKH5wcsTZSKZxOg6qJccTwpS54dc78S6YvQHNSUjs+
/442tR6wiisQaj/7OklXsLYA7Rx1cDCpxpXruTx8/ADuqh2Yc2yvktDb6i3rkrsoPYHUvPkBcxqx
W2Jl5OAcmy0Ujhwy088gAGmRz6QILSUOPrUN6+D5hBs+Gk+YXgli2+ELEokOR1w7HO2XuwweXkiy
+Ezky0OCbn44B42S38WJBcBJ3CAL5wqTza3kh2dPPiF1S1s/fSaPYD7aE2S3ARLMhuMAVtROoYI4
wXyjY6I6NOM5aCEbe6+X1Qeq0TZs2vGmGA2Nku3olOwYioUeDscVeUdQx2qUAeSxcoXCI0dYsBzA
e6reasTfyr1x4KSftR6837cWTM/+qGFsheluzAtfRFS/kT+dLoo+pDr7wNEcRRmOPAtOwydXjlLh
rJhUYCaMdm5aBgox5c8kfOsOUkYTgJyAxoQ4pfohdfuxag1O5X2VJttTWPxJUyPl9Pv39T/bl+T4
XwVx+Uxo5pYchxIiyP1jmPE7hMVVoSNlm6s6y3oQotppJ2+ToV0jXdZ0rcrEV3UKqgQVZUtSiqCB
/KYrDrNXqUEsyOSMHocXkMHwi15UairDLZCxuktEQh+An9nZCvl4xCNQUpKJcuwhv4+t6lotRP4l
FGQvI7JJg6yiX2ikNVEv7xtnSnyoFRR2Wk9cprETLprCzr5aXp5WaTId+k7zF2wRMCfZ+h4jU/Qw
OgKPMX5MWZjWdyQQuZCIkCqu9MhPZldanl3pI9X/r/Vt1EzumIIpAZ03GSjZcBro1QqxB7xrCyHk
xLLe6yoTAuREklNK5AwHe30UlCb5ZKOkd9WlnZr3hyEUfn0hlCLZgZCK0vFUbsUBjiA0zalBScSo
OVGwdhe9mUNsqi0OW7WLkcQrITEPEyIaEzA1wdG7u8AfI85kKXAn4e18tPI1wBVwZKt2Dr2OQbdT
HSTRZ+92LPfUqZ1uc549l2PXugphCuZCfRJeOL760beBrNqGEjeDTq+cw3ohE5Bao/1WOg4E7Ly8
lobMs9hp7vg7snwDsCxcCXyH/sePIRNk+ML+HM/q89fTMu64I3STXDhr0jfeih0ESMVZ5LeH3voZ
3NpICqBi2Wg6EMoIddjD2AtbkeoqykkW/g/6eiC9xEOku6SEtiBSuMVWDWXhTzKYRGGF7dVtweWP
2CYZrZ2aSks6oYQYCW3XxHsDTjO6R8qKMJvKCjSRxgKf/rFmWdH0uZnj96TG1na2M7xM/km2iygS
9RCpRmoa9dmc6zeoeyRTQNnB6ajLgMojtOff/TWPpCcg0kc7mq9Hdu2RwLSzsyO7Zob21kXe7dOV
7nD4Xnl+ZhtrIR1UPf47YIlxP3kJaYp78cdx7W7r8uQHF2m7C1zb5gnI2Nri7AY0pnf6fO9ov8ua
XouIl7hSMcF+igs2iC1F9+x0o1Tp0icp7hKRLH/+WfxUsKY1ylBMmvr2vfUXsAvLwU/1q799a2WE
RWnNlmPPyxWAqn401QWnnNFKsYa8UbEN+A0yZ9k8zvJFmJwJjWnB4cnCIh4RawWuF6AWMEt4mNdD
e/85yO3lJcjMACuukorgORqpxRt/IKe8c2zaCXSeHt9gd5JoNZ+Ui7B1hb9qpsrtrrnb4kb15pda
khbzGIEVUen9hbNf2CqSzM7WRXMHNzjHPpoFVRgJNBAnSfombkQ5r5+3LfVVEokokDChdf5zBPqO
JnXPcAaOKTMnLuCGePLdAgR7M8gRl7zBLnYzRM8FB7jwRyQU9XBt1L7znyOCCBsIO07CHcgoa2mT
uVy+WmlcWhsuWN4RfMaT3UIyFegRctfRhHyypvUMq0HsVuw4pbE+KN2KOnP812+R9yXlPAQVr7Ff
RL++aGs8aDN5J1abDNVQcFMwvuggByVog7IV6KqpD+u3SKvUIF2qk/ti2mBtgInbYfNtQFnCcLi+
5fddz7kca3/FMhtptCnfCKwkINchtceTwEeKf4kNhR+FJowrepl1iBMa0gAPeGUT2ktNp0j3B048
JYLs82/Lw0mNnz6EGEmTP1IekAtjEq3PWh4667UiyNKIHl+WZ+SVtKiyIHWdKbMCotlezsSkrf7f
I9tsOmqfarIqouq61q+Rj6aai5dI6OGCOWQFlZSLsTRjJrrJ7kkUswgdEX/iBan6KWhOFuApUOtJ
NwV9cbLIWbvqDuhz3hh4naDKzcierUwSCZqVN+fzbYEuL9m25sgehueMTLBZoLu3DlCFBptOfpxa
+laFrdtJRkAVYjWjOPWsDRsdCtfGAjESswyjzzuJ573B8QCWVMKeySUV40nNEPAVCQ43xOzisXkZ
OI+BvGSgeq6c1NX5dEX8hVyU7uYAucZvhmNDn2ylAx/HnSKEL/zZ9yZ3QLTHJjAJOamLYCkKpfpe
Q7K/EFiZKOgoG2IPF7kvHShzfz3yKShBxGLLRfKG0ep1oUboyOZsl9D4gkp+ii2EMHHkD77TwVVh
oL8ORDIkZiskIYenGVJL32mf+Ohb3Vh8NcttqmoAF/gpHKJkNK7MAIB3bWwJLQqboVJKqIbuXsZS
oeQqGZEF9I4MuPwy5Hx0aLpDVcjtLMUrGafHb4b3Q3g0jJ3Z1Fv0baP3+XuTbVkbZTju7R1yNE2q
rGXPORHfHc+et+yH1Yome0oHuUp3+UWQOfDCY4b51/+cMrw9Liy1XeYs0KasDeiMTfgaHfHsXmeL
eO1vSUVYK7oisx+6JL5rwtM5DgG/BuuYS0XT2yfwmSdCNj0pDb35edsN4u382BvVccrH+mIDcfZw
v8b3xMuPxrOchNVG/Lbh7tT5FH2gKdVNhSTt+qyuovV7j8uNOf0gx0VfzrRRV98p9CU3N28zKDvK
gFYZ+zcEOK1XkFUhWGXAgcNlrN+soes/IAdY2eo1ikXOSRAalOG67YKvo/M+2M5uUw5J5CoNkAR5
yfZKlZQYrvRCkXjZgAIiD4yeuJMWSY2egEAnFmcZb/Jt+DLDlEuhJDzEjSKL42estI4WomNWYeIn
e+5zYxNGtqFV2mErjkTJNDUVd3Zwrb6UZJI49tS+17J1I1ib0ba/yC7bjkyK2jdz3kmPJsAnqFRv
m5CcAzRkpSyYgqN2c3UwoW1aO5nv1bDC1W2u5g3vbaPOo1LEtcf5ImNY4E1KNVnWI4wPv3Zolp4j
JJCTB0gV6RlUwQ+X+wVA31Q7Z3pfRohtQQd6Ur4eL7QLNRgiZ3fGTA6h3OcOBLVnebFmkMhdYLHw
u7vcGyc6RTvypKo7y5N5eOmSuxQDDrPiWBpK399C7biNWut+YIzc+CMl77ozkGOm8wsLmOL8kh+Y
N1FoTavPnU161IgpABajaQwNBQA6GQz39u+sj8sOZMeM69giEDsL0n/Adgq39doAYWxsqqy6Nc6m
TESSAnzTTayCvA/tpqK5HGQjLtuxl2744ROyDHK9YjQH5osiki/VI5bIMEgXVhnjYA6qQHdo0or3
CTZHPz3/JlTKkRvVgIW5GzwudEXG5oJGLG7HLivx71wYiVyXLB1HzdOQz3dX4zbUxEk5R6CqFolT
CGRs8j3IaFXNNEySrfhrgC1jIRIl21J1RcGCJzjqxx29+x1PEqM57ioHMNNXoGri3JFqOILOiPUs
q74gk718PJBKXtZkpVpiQ3ALjSVmynfzWzqD43useTMvCDTb98A1AzeAsLLBaqlZlbdWrAv/YNor
VXc0bR9VSU0WoxQJYB/DMX5st2JQmKNizkanG1eFbYtstze5M998dK7fEA3XT9U+azWp03k8miL/
0DFvSH3fU8GZZ33F6J4+1Dhk4BGDcMU85ybu8dJBPqPJ6Zj+HEV8iLy9hlfy2Fnvr51VL+F7IDFO
UY0Qvfp4BdbYphQvvGHb/1y333G+ksTYGqqaS49vOI4DpB0E81CXJxbb67FATDkNes3s3l+3yzFU
Xyllus8f6JvsSuymg2jYNaubk7iioO+aDPnjH13YlySS64NppGBtZBazvxjkQ6O6gSprJjUi7277
xeGw04ZxKdGbawxb39DxrXOmMRYc30MxLQfOIBNo87p+JyjYMsCLiRJ2QAnFCbbwvoJm6ysHDsam
g+sS2hYeRlYRIyCo6zXNdXbho2g0pV5wNgNDRWqJuFOYl1+fWo/lB6An6XWpMZX6cv5VJ60Ayk0+
C+HIxZmbFpHyXzVYB7tX/E4RHOy6JQfpxVNhQ0JgMvNWY71OOh/4Loih6+F90IEKpobETlpk/jL7
WQ6/Fjhgl9KKATo2aPiRBnDWYQH2aXVD3cZrlYUBGSBk574SkbHUr5iKvRu3dWV49HqLX8oXSL1T
GcojWIApaUIkG5nC+Kuma/EJVGOuEMy2UOV8X/yKWE3e1AKWU+a+YTBZzsgnTqGqicU7Ng+ckw0y
IVy4gffGo0t8YEuZeUhRTJVRpj2poVIWe76+kO+96nZXBz+bML7X7+Rb6oBVTsB8GxIbwZa8/Ph2
CRvf6M9sCHxen81hO5jg9ijIl6q8t8kT3y+xH9V2hPjjDe3elI5XvsLjhUzPvlQGdaziX2/iN32E
eRvvVK/lKKpImupAOmhX5zb5qF9Ilj0gjDzNbB3oq11wWMbdv9FUMBSE4lZj29Nm4PwYWXARhWpK
iy502O14WG+ITRPtKiPIxZIl86V3EfccjS++Z/vw3xbw8vxsML3Esow/zFdRZSB7ABZyxox2O1Uo
ycG8eHwNS/nKa31kvD87F0UpeFWM87ue0cPD1YrnW90G3Uy4lnXJIml6CxB5ORytXO4Kw3kJRniI
NlLg+egSo+0IX9LtaxMPWakzVAvRpmhFyJfXIQxq0Z1+UMcwABJcH4fGf5OqqH9Qk5PWLYrTjJga
qwKU+w+gMnIr3iIB6uFOTFu3hqFPOqjzHwR2BRqLK7sM7oHqVRLUVN0VFH4xM0tcG+Mt9pnhphVU
5XnhYtNeyEwP7gFJ8BA27yqT6on4B06x3Vj1GcTnh8i1Q0GUZ+u/c5hz42hHRZcdq+D90dOgeO+e
uCx0yNqdqFg3bXXG6mD6Asov2cdKTpPAyGqNF1GLSJ5wWIciOypyJOpH2NZrq8x6LA7t/dUuiK5Q
GqoXMjOwRDLrIzIFYhfZpgnOmBdqpdsEyCxx3UqxarzwA3Z+daYTJw8mjmAxLRq6x78noeS43/R+
2q2zHOCX/+QpsWmIMNQ6mojZk2Q25lDxFsX07+L1/m+YdJVk0mvaxEJGGlq6n9vxsaDtWzBHXgaC
oAYfq/fSeI/MWdLKrRq+2lpBP6YA9O1JbqV0YxQkhN0NrzmFiS1ZHCcmcqeDOzn95qUxe228DsNE
0OkxDodyr3e3IOjM8R3NTRq9FYStngj5B9cz8DLQ4GmWL6EXugowaVBqu9Ejp8PhOEkXqEWpIXIH
i3LJdTnjGjaxx/0H3pl9xjJ+UgPvp14u4xdV5vsqcrZMBtHXEjYe1rbiJj6q6WPOGj7+qt8SnnCj
ahvDj9Xm5IIJ0KVus295X09Ul7FG+Jm7H1ZpNEJjPTC4rQ2C5MRcg4zzmdwEpqLfmzqfEH3ms86f
K5pIKLge1odtCptpgoZe0YUy9aiiQVurMS5XSYCLlo4RcfECNszPHzQ/pK8NOcBw+72efcv1fd0k
k8sfJhd7pLAXG59OtTb0Ovmo8ukd3nnbbde0UL8d6ch8w1QeX1SqurH7PyW1Nhnd0zguS/45HUhZ
5nLRV2u7ZL32voD9RYOGVP0GTomfoB1U0B7QtRdpDt3k5eYxB4/g/bTmQ9tbH2cBtbvGtT8yc1tU
xVcvQuQiFVjURmY86YEMwfGxrdYzZvP9ypdXnVtrUcQ7x2U1TeMQLFeTw6aLWFTDmq+Df/fFM/Yu
WL8zTDNcuQlxh10Vf2iPZzxtAmQn+0omMRVyz/ise/lMXCrgDstDb/LOCHbwFqJ93OhUWiuAOyJh
H85Nv4V/C+Vq3X3p79aONs+YriP/QHmLGxGeNih0LPzmBrhboSOgtjgf7lpVrRoxZ6golPrXeVh/
5T7ynsXV7ee5Hxr9sDs66l5YcGLp5T+R7kYbT4f4LqhlE026CkgNZnhgV6lC5qa341Uw3BL8g0Cp
r+MXVOn7DWCt+ei/+JLfKajYSaU+wO9j05UyQYe902GlDSaEqnunhl9icNZpHSm8hbFJoxthG+8L
QFVFHXWx5hMg615AdP4Lxqb6pDFojzdZ9lgYP19X+5hChVMTEkmTU31DlFuGyc2KbwrSv9yMCBmo
V91XAIC3AL6GXo1r4wyiu0Nspw8hy3tMFiFSD8yaVNkdpcEb+Ku6K3WOkgaDqh6gUQ9hjKiDZYuv
4VQebx9cGtrMXGBFlzrrrzK2rdM8G2F57SLLQEuO2T36GtTJ5Gcp0ACVWf0J8XxdRBJdRH+p9Gbf
ZIdDNoenTL2XVF23UW5c0VxmCWTJP753yz1U12C+NhWGAhbKh/rfKQF9yxAf4CSJ2voI0PqARcF9
Lx2ITaJFbGQKLu++YkKbnP+vdnIHodB+X7BMXl9Z11kQCfvpzPDpSP2+5nB84ttYGQ+00Q3PDdLc
VCPK1SwT370LlzTbkboueaZmH3CXjmDahLidgOq5tCcM/x0pHDBIFvPQ/RyEAU1n4S2Q/WXd2d7v
xPzNXSZsW7RGUelM5YhXpQuSywSQ6JyJmbZG6dkVI6hQ7k1uSGqIluyVXKfcIomUwpdE4ZJXkuGG
ak/SJlRbktTWlF6wo6FBXR72ftHCSmD6ZCnJculnez+Jb90g9pZcGSe0yw0rB6WECAYp9IDclqZk
kLKyACU31PhZ/vQ5eLTRAFzbXuOc6t7Pym/7C8RZPQeApl9YuzEMc0IYW6/F53bet1TWWWNnVJ0c
hwkiI8fitcU+akTxqRFZdPQ96v4c7n+iWxzuhpCoglACS9xe9Lzcxx4MYVlYLvNwi6p++qASnMz6
Gp4cpfeK5dNrW/lOtlyzgneWTUnjzkGyuTmjQzEHRSUj3SnNZT7onQ6WMLoLHrwbqVtiyOobKoEq
tSqGvtaFBoownOXzMpcmmVi1fJuPcXJRaTfda+xscefH/Qh1IepgeCE78ZVi2b7bgLBjrsyEDWYI
meyDOqmISAr1p0UFoNdMUDjjtOn4+qFqCBIGXo8UTEhs/66gqnbSk5mpYCqh2/1nfd+HxRK6kAwf
aDwoyvng5QOMGE2JE0B7CUfHX2Vmc/iU1lVVRt1B1GqBZsqoYhMRBCyD6yebRl4/pUZ08qDblO8E
u4E9cPigF/kD0edIOSz7keI3eSwl8ai4v+8OVWvJTT1CxwhEgh17uVCW0Dq/2Nv61x9Ht8Md8J2k
9RDf9dqsC5Wm3nDf8rmYvkjDyBCGpy8YK1DaAPdyoWi58/xjuOJHvDtv06tLyo9xDp4y9VUmMqVb
vQ4UvsVeM9CZV7V03MXRGSaDAkeIAnHyjLa8bH5J+1lffBWCQp6+lgOH5H0ebbdpg958B65C6ylb
HmRKMFUijiAu6nqLDdF+fw8rv4EbZGZKgSUov1njgx8HQag1IlMgYfVo/KrjbSCABTqJAyH2lWW3
/O3/xE5QJqT9fvGLRewt2BS9JeCQ1vaHRP3VkfGnfjje8GzfwPesXsh6kf54YUuKQDXbJ3B5Ndi1
iOdqj1GustIptXrx/EdRvy7fWrEGWvzJKH4gZ1f8KXrJVkNXEUQ7Emu914NQr1DmorlsG5DfSwyT
PoxBkXCP9ZNJihAVVzT9nOSItRb7H8K5X+sEd1DNxHdDtzVkhxfyse1zRe32g29thgDoCO1pUQLC
7ttIHNNKoZYmo4XMM0Jls+STmV+dy/zlqFrOm6HZ8znfLx0MQCBkZw2y9J0pVrVUpi0/X2Gyfm7B
8l1Dzk/cHkdDK/pmmQ8pGQvtHP42dAFHfFOhc+SxzDczxuPVUKTYIsWx7HFCKCqYYcCorQpDrL4g
BGKhjmqr2dmoMZU8xQHBlV1pez0eC8U06hEyxDAI5Zq8p/1KmQ1iV0opAn1VynMbjY9QBgOFydP/
yO/DMDymSfcj8MGergJ6A+eipS/NE48gfZ/0xzgBzjX6wWrLNbxm3ag9IyASx8MsOkf6Q1yPrIky
e8ZZ5ncIGk20g0LCeJLZBfgZNHIx54cHirHl0DeUQ95QGq65Z5x8gzpWZEiJtrAvgqdmFsv9Qe+t
t9lxD7fJMOZz+SM/Tshs8ScBE2yC2ijlGR7bfIonEJajPgpwZG+7BVBM8DFOayNOdPrYno923byh
qJ+4HrGKy79yb/WGncX5x3jZCFltcYMAoF563TaxOi8mxP6JThfvBT602eDO3+z46XVsUox1EuBh
WVIgLzs3NXPfOs/gztMYpN3bQBpxi8bgQQXYBmnNWF6mgwqtjI46SbKQQ6WwJhp/XtjqjjW/gA+5
uSm1iIZLVlck9x9J2I1q6XaA7kQmQUvY2KkBGt+D7o871/TF7jw2o+c7314748zfUft2R5qSSfyX
GwZBYoH02FUsI/kbYa7q2yw7FVeNVENnGGNP6Z1rierFm5OpqAnhwR9752xizLYn9OxvnO4/0zz8
/PCLXSD7/egZTItXOD1IGKflkXdxqdA75ouDm9AcvLxGvYADuQBv8W8bQv4+fZlFSy9mEpj+a5NV
hVTnKUVKBxOwZYFaRYfwnoFQ/epX9lPrgHAnSk3QWJmFDmYNunK0VcUPKAblZWMKK/7GdYqfZm+J
dsieQSJC2iTJlZbiIYrd6S7hI60ObDZ5JV4ZhTjf9NNkpP4KtPcUeKwL6scUkj3K5L+/g1tMyq6G
Rtw6z4cpAgZHF02ezSm3aSnVwYeOU4hscM1F8wbxKtIXVgTKIwXg03GEWXyy6rprqIYRj6mNAhoS
ELJ+csdRYZlV3TZPVndBQ6+aBokPzaRUaUT2DMpevGQQneh0LtFjxjpWnoa01iMljOAyC/XiLvOQ
83pRcPwLCW0S9GF72pE0s/Mhc6GCpx7Tw3aGShDd3T8a2JyIgVr30BctanEr8ZSAER+29Wk91xSh
U18FONiLc7C9WzIP1GPXO3yVi+G+Kvq2PxqSD9Qdu9MFsIUW6DBdwnhVMwEI6NAHyVDX1shhQYB1
02fQ1Z6TcZBDWIZhKS6QvCaZ0Oj5lW9KEqslDijxw/sfKTmcr/FDX8lSiPXc1xiOi3ABpgpwtG+T
Dmga7iKHFXsZ3i6L1Zlul9fOz/hQccRlDDkBzjbVZV0rr/m4fLow1Vk3LsTsrkM3QrOKcuscJeIU
GkyZUnm80JYH33SK5eQz9TQDtDyA/PBPLQUUQBGgVhKV88yT0nvhf9RH686fUepGbJpf0A/LqP1M
rM5FV+MVYYcU2CuhC280tfx/Auf7WgU34ruaprC/zZWDrYSGmMOlNvYEn3+umz2J+ZBDd6WyhwYd
87dZ5waH3Zk47N35wVtHcT55o9LstLAcBZ/ytF8TFpAkt7lKBqgVDf+SygALwZr6Hb8z9pukZq7P
KJnTQ7f0tiAyABhnmRhN3yzOp610CgsOZsN9pdINreq2lerEP3n1quUn3cLBXlb61KqsS+pF4Q4t
Ahtfc3Exu4J1sr9W6G5X3BRuBA0LoTIC5W8ddrsnwTK67NBEX0WOiKoCj777ypl/lmdctHxXtkLz
SWWOH4Sgw6xK/6x/vHJRmEIwqG/QKVfAvAj6fkqI8ZY9B16t3BxlPDUtHrnJhiDGUB26KcvHy3b+
10RWuLUsTzhC1ppOWuUbGdQiD+DwGUU6SH60B5P6JS3y+huvSCOViv8VBSuzfDKDyzTs7TMvZNcf
p1nWf6SoueD5Q3k47eFwObpwxMvDurWl/P2iFKwrKkjvP7CH58C6T5pBWl6lRl7rJ/DT0Q2nZi7v
yJ/X6lCi/NiDYtNHp/InroyouC/Ff/oplz/k5evFJ4y3pilXDcPU0c02AW89RDsAfOLKtnR3TeAy
t56t4zCPlMTQQZbnUqnKegzPk61tW0EzARGOGy72RG7hFoqTl9k3nZZa33+K4LPQwmwb3c9dF9JK
yBGmZpAz2kcLuazNRlYpyDoXowUWlpGoLsrxLg4o+/7b1ELY2QjFH6g/VWeoeFuDycD7rQqaKV+v
ryGVeM3QXIFcOytJuIEn8u1c6qjAFTqWbJYDfI+QLNgm/FK7qCKuiViknU6L0usr1Utl283FzKcd
W36975HpF6MYBrt76W/zna2BBSkd/Sg/PVjHE1m/PP1/ggJNqvixsYzvLY4e/ZhJJUjUXAgXSbEs
B2w8CNk2QO2k/Dr4Kzq2RUMDwHFBa4VhG+mQ2qw1DrBpDh5YVBstJpE6V74b1eIIvOz2h+dfB7K4
xma6QSfO1/SCqAomm2bG3b1VqeF/L9qwB29fEpY07P0lmF3A9YDjJp3i3moUPHTXZI9Rk6PAz5Zh
RTbT48U89Trb35K4uk1Ca+dP+Cf5kdPTT+EaCR4ssR/uCZVMAMkoiuzIKO7hU8wc9Gm8Fx3zInQ6
/8hmIFzUjNU0CVcRmLTDdo3eWqUUR7t7AQg4dgiIYa7TZf7AKfMVMSqlfXRNIxhkfuvpTvt/6SEG
Uk2FrVWaopZoGUceSYiPJMSIq0ahAroTfEhOi7TPDHcmWMnfAPnny6jb4YPDb+IcD0xzudMZK0Yl
2UAeXHB83g4qgXcuSbmojglQYBp0e4xAtM0PEdnlCFs61nZJ/Jo2ZCXSqF23C6KPJTkd34aZlH3Z
NdICOEGqxnQK65C3EjezGH4G1j8uwUGTtBHZD9DuUVIaUeYCBBUK4U2yc1a73Om64zC6DfHKdYZh
cqVhw6s+qM6GHIkx/9o1Zy2NSekWxL96FDhDqzg0RW4ie2yWWuoc0o//IfE4mfN11eEnYZss7/Hw
kkPRiCvVQm2ldQN+4Xx3XH6gx9W+MOZJ8uXBhLO9MW7MClt67UHOkLnSfHNm/sdO710nZDwkPRSO
2qy5NjYvAgt9GWfRAs7cOoTTqnYxxsSyGbD+5T1XaTIgU7o+m6CeLkLZYc1L/+xzZdyV5ijbXoa/
OO08tdEVGuTem5IJ+YWW73re15P7j3ffUnTqtvodDQsbDTFTwBycWRqi25xb9h3OpMXDPjQCiUGd
l/DlwDiwf8XZI78YzG00fy9AVqsUhA0/bBrDn6cAqz4ii+urj9gMbP//SoL5YPWxot1Uf5BRjKRu
q/prvjsnrrn4CbOL4IHgqLkentFPH8QF+xlCCXAlhkV2VQ71S06I1aILeslf35C7L8suA/x9X9Eh
tmtdJGLa6LnyBIRXo6K1CZRF0r8FQYoqiKgDUkUNcXkLGgLN7Td7sxgqRN2P0k948mHySqQ7TSC3
noQfQZDO0IyjTzaW+kadfz6k69eplEo1VjMv5oRtGGyc2zj00SJ4as3o9AtdzMO4q57oOLMr6m+i
/jW+ljQhCpzKXHghYvfE177o5WmFlNjic2bkyzH/bha5vBWGZQ1XqVYRXvYMYEP4lil8ExbpuZQd
CsBKQvnRe5x2qTgYlk9lvSquDksDo1H0zMz+xSxcx8fJPN6ooePp9I+5P3LJK3yWMqvoWYUMk1wY
fUQpkrASUWU8S9SVhPZW3GLrYEmTyX+Dp2mdXpmjdIWsQpiWTFucGuQnITLp1dYL6h3Bm1AcX/gV
3HluWs2MAgcx/NfWtgtFi8gyW96o05/Ru7y7THh9D0c7a4Le3fAhsunYPYGPHUDZmtMCIE2OmsAv
ZV+9unkbviBAMJCqlIXvAhgQeOu+iDSOcRBDPIxOOj/51ubJHuW9Fo7zygyPhDO4qFdMP7M8vOiK
haXd7G/axQWkoenZCCe8gYQpHL9zn5/kztIPMg0sbAPnzCZjZOQonfH/Wnd5XQ/jy95JpzTAINn8
HzYt2VxlYGcc037ME9eySDS0qc34GNx5tdy5Y+NxvEgg7EIplnnr7TvO9yB8ujRHMWJeQ+ET0GRz
zKrL43ztIAJB74BSGwRDyeZw7xUqU6OGxPSrxgXtPu15qJ7Zdvq7rFletC5nYymr5PRK96i//tMf
csVXOmPzkDp5qG5Wk+zxYVW2RkQZhOoXxhkHhvXtxqfh2ls5eywcC6AYDE/yr6am3A4xKcCmG00m
QzlrWvQ+UvyPZRpGzkQRZKxCPFethVWf8u2KZPMaxf1kze+oaKHfzokHUQDIjXGwGmInIBGYcsxg
De8+CV6SJnAmu8Jg8AQU8jAMcesKmj8tl4DuvOs47q8GGbahAUZ75LcNkkCnfvDWRFxOP0Vs8unS
f9aeRlph8fTnwMMWgE080lZY9W/VIdLGMqjEZC+CkZEjXiNLVOdE3lTGEMhGi2/gMbMLs5anLdA3
vJzKOrehjm1J/9lWWomh1aLukzG7ZK+OGCog0kJV+xRVUgGnkukYHMdB9zd7A0bc8NETixX1xr62
sWEmCZpb4XbGBJasLlNQLpWY80yAed+RXym1OwrVaqfnvYERMz9z8gXr6BmSqVh6FLAuHgU2dDXQ
Uw98dOohWZ3r9FgEYDvp/R+Mc7iyL5lLulxk6V+jQ+cM4QZjpFUUKe2UIFaKUGaQq/RyseL6UMz7
hLAdoxhNCx3g+IirnCQcrhpfGCruhxUGrdfXMovTC1TmtybjhFA5/OsmPGOwvhTQUHZYW3CycqkN
D+dbZaIjEKCVTiwK/LxeQKBJveD6CjBEJf44IXrUAgjEUc7t3JKsYb3MAWtOIgQ79KKKUXo4IYDa
0SrSivPamaYgYC0M4fHx3fShCpeRQY5spfTdJ7tb0hhgShCYnc8uLWqQxdpEfVL5NszOAQEWtKSB
a+cZk/ansKv/AwURtj+Hpka8yc4OQkLvXORA7BlEFB1YfY3TA/kqRkPZxweyFK8O2K1csM06Xy2p
uf1lxe0E/gEG+skO5f7r8eG3EG0XoGaT4O9hsQL7AxqTY4QKjOP7AEHobpbdEMKOvc4xJaa8Nxnv
PsjlAFKC6tG2vmRlnurkrqB5PnQZ9jz8oq4Zw60y7lsa3mjhG1ybp0ABBejVkXtDEy/ZrLBLUea7
AAsgaPpEffcx0+/CWWZQ/HQRYrUHTjOzt4un8QAQXN+kGxdKZKMRD5+EgzrYau9X+SGg+4UVPQlo
Gxa95nOapVtpvgpM+lrRvb5xm4WEa3WmZGENbCc+1O4fiRXRvEAALikuEVSMH+7yp6e0Za0sFaNV
PiduuPch9vzg1B1ijjNvMObFAsE2hB7uYuIrdbiehXmcE0JGFLhKYhuKNeIZ1f9+RPt3hR2wiJ5E
mcS0FSFqHR1uPuHuLWd6WQoB97InPyxgzF8JyN/jIBQTVi1bIBuUictUqP6l6j9u2HM185Jj0m8G
E7INqLtIzO1+/dtIZNmD91dozIRHtquq5+RwXYi4zZUdlEulUZw1TjdYTInic3lSn6A+i+EGJsFz
gTsCGTdJFWUIcyVg4oDAFjyCOIKqQPQhVSiMjQKPcKB/tVcb/eeS8u8LOAZFI1fYaYZqXzz4HA4U
mlQ6F9pM7fRHUSIfVTflvFNhi9E/JJjEnWyCNaK1okSKX+N8B26X6AfdtLS1+hK5yeqqPgOAVayU
S72kregeTBlgicefJDi00Z+FjzWsjpit649sn1uhrswO3aitce66+gUlDC1bdtkGAlzmo/bJNO1J
c36hPpRpP5n1p21xi7vGJIGEqsXwOb9BiyISA1aB/LzUjwcP+7IJ2TYYKpk8LMw7H10zPwyRE018
a5WcbCQOQTppPqdQhM+qcVfp0IFhihsA7DgPISRXLPobnx0y1EYLJr2wJd4M6FgBkK8F54dpFx9s
Q4DN6ZaNn8/XucTh7Of607Ycm6Nzqw0azcyAoU66oiIa2rGROxKZMkoPnYoSuQ7v1o9EiKaCZ3p0
G3eMMKtu9r9Lff0UuPjJHSF59kNmYr60IyikOix2glUVc+OPgTDo7c8EMzptLowxLVlX0neuwpyB
D6PAGIsF+mh+XADk8drgJtNYjd80AxfAWLipZvYt3T0+1AiWZtElDh+X6KciwwBnpQOacUqiyyyU
sNxoVEF/7O+JnndPWNQZ2CoOzhi4++AvfqCJMJzCT7EOVH7Xp/jhMSnrX5xH83FuDF44IGxE8krP
oLxeWBKxOSG+ljADlyj61Gge+NkOspy3lR0SzNaGoyljTI9YokEy1dW5HWMOCUptwQWbYAQOBUsl
ib7MMGbMSUZkZ3JvWAU3tT/r79ULzt16F39xkf0V5OlG62Nmfn8zTBpvm7aHj0X10KdibXE7oZ64
A5Db8R228+QdTeS1YamCfeym9pHPGSrJNUyH9ZGR9T30m/l/H6KlDly1Iac/h+vIhS2OSW9DihFu
QCzyz5+tJnr1Oy7l+N0wQIkEgy9N6+zq5+ZD1UcTPGa1OkU83/8qbUJuTP0iyu1gXF7G0Aza90tB
73OBSqq+KvQMt4PaJZg+iut9jC6f2QV/3NlwU32EJlHRna/Ez8btr71Lgn78g1P5cHnW15Hiu4hx
57k7c8l4mDC+ZoKZ0/bjDCt2Wx7ER9C60MjpHLNRI98+a/lfOKGiTuOX+tRKEUDVYP22iBivDX/Z
Tkvu5AIB9ga8A/8iz1v9IwpPkWbS6dHzJqLg7uTdv0f1hNRLt/buzfM7dsOImee+Y7zlIvI1z6W8
SCSXgAH7DeZkjSYuLsf2xTUru4AcR+GRizB9J+2claj/c1JfyDhK+uXr5o+ggbHkivhz/27bN720
VqK5z1aELAbroMJs3F3VgA1E9Hu6F04pNc3mD8bBHAk2BRrFlYtzPNnzSgesOFeWpQG0u9t3HN/j
iSCfbCv05CiuNU50XO/6jPCma2QGUIGCU+o3e0Tce4+Y+nrRBqnvAHmSd+jRZSirQushPruj1tRs
4uUjHJbN5UvNk4BpT1qfJgVzHSDW7lh3drqkVvITF5jbTvctZdGmQrRYYXVbgx/nYe1PfqwRQu2q
gNeJ6kCAmdO2bGKytEl+mnd7hEXqBkqhdFrh9o0WyjvYg8wCEJEOwiP1Vwz5kRKtQVThUV1WP2BZ
YE2NGsaKGbXu4EFRiwaZgLoX/gbiCHt6/xD9AmFz43s4m87zbn9U2doiaPoOB7oJ8keqolLe/DcP
gBYiIX0TVVlimMeLPQ3Bi6OnxdKeCJo3gKdjTqdcTUehmP/CYFP7WmohyukqAU5ccLkmc2D+0wcO
EgAJvYKxek9o6ym0Uro/0p6F3XCobdkVtyYTiJb7vMJqTSXUeImf5OaHKu6EOKAjEOHrxQciYghL
7tLFekihy0KCmrMHaltT8AqMU8/aRoQ0/RWhP6MLh7OF878TWgiKjnPLpHdTY3Z7jKx9AA0DrJ1o
gdZ5tPI4bt8GPkU9yJLVIanvwXKXaPQ8WdmdnuP79aWLY0FsEv+0EYDCZO0JN3xn3ilFxiBKlWNT
H4TCC/5Oj136YCGwvNP17NVrcsN4zUw/zkL9Abp5olJtamm4+DyEKsd7xFuglpzVeNMEbZRU0l+z
NpduMznQsRiQH9xvm5O7MKY9D8WvLUyuY+PyiHM8AEpZ9YoKqMz1gmBxpWmDBZoEXpIWjV9wigzn
cKhT47101mKDAwR6cKmggu9sY1K7ktDsMGRH9z8/NChevjJNqHiR8duIFFTCSR02cQuN9zMYdVsP
vGzhYsxV5mwVLVEfnESzrmflX6VajD9iUFxuKo8Qp+Xzv+fF1sfE1Tw8+im47y5PcDdVm52P52VJ
p0tlGUIbSWIHHmagA2qE2F+iLNnxr0SeLlkacrifh5vcdF20m/B5WZ2irET6qn3NX2KZ6FrtsnJv
P0NYa7ro8Tcix0B31FfzInLMySZmu6uh6C7xGSbPmjCSqm9IOtPaFN0SmHzjKBZrPhuwBFOFW+RQ
fHJ8BC32BvnugDRbbUEw1LvscjMmiFM98/qhiQbtMq2VO1UOz3RnjL7TJC9cKVwZBze7E2j57vKw
hUxP1rgXCQtxaJSrAGNUdfID7tNzhwqGi4vurtO9h4xzRQFVYZhnLIY9Tq+URuZ1ktFReks04uS8
w/64eGJLgpE72wRv/XillQGwb2cFoarRU9vB+HhfMZDHMbN88woUcb/IVBO/KVgruT50ZMg4fqXT
709tMSd4Whiqlmndh0WGAidXnx6u5T97Dv8wh5UDThtO/M01cAm3hSXQZFXGv5CTTjanICLo8/lW
g/BypTO76g60xhIMMVqUaxrxHVah1KuVF1kcIJS3VDOVtXMNqKnIWk03OqcZNIYfcayTQAEwNpmj
GkTtRoLYM0TGSYt3I1VWwCxHLO0Yhqq8M+vMSAajk3H3s1DTjki+QVsUO4hWCtro+cS2LMZ7l22P
Bo+YZ6PoMKPk5njB5K/5CHU30TGu8g6KD0trmMv8hIDmscWaH6iCleeTYdakW1z4uix/b4Mb1FOS
o65h1jrXo6uBhWOA4jBpkVhV2lkhfHM50IDIKgbN65evq+aI5+ohUkMOaZNhKY1ZkEzbKJvJqv0K
eNXknpkFxSChIwUQat60Rp178D9dfJuH9S7OfEYtjyC7TuF4N6SY5JY5QFJE7Iz50yWNNbOvFgZf
PsfkY1XkMs4aqPjuqNzBLBkD35uJDdDyfYWSENKGRydLHrucKy8vjImLKo1qr0RtAlFxdf0LSmCy
3bIZprWAj26VFSsrNBmdKvj+2cSW3zdKJH5YL9BsPj6QprY8CoBhVQ5Yefq+lusIxKVj8Q7VW3YB
8/hypoQm8pAPyKQW4ncM53HknP8fBLPiDkXHECCZeXcEMmMktgRZlT27rjriaIjtgsTY3cfdX+UJ
QIk+8ATPSI+sIRbr4ZhB7yJqgGYb/h/SF9v32d8jOEPVZQkvsC4nA40Qdh/0oG9+SdMUacqc68TO
w/IO6xB1oI5dYUDJDYpN7dRl/NtOpTa8Allq4gOs/5yqjfQAeoQGsEosFHYezclSKldORrqPzRNy
RSwGjG889Tag9sIXMugXrwcRxPF5pgHp97SRREaZjM/M7clOn/BqUqRR5zvsuDrmWxzmppaLtLFj
tPUO/I3kU8pYuSfjGxGH9E/LgWGLDeEM8KClR8TEEvJ8QZVrRLc2IR2GBQdZ7dRRrNJN2iwH7Tnr
Oufeb31uUcZuslr7WKgkn7CQFJfo6GyPirAgR4d27WlqSfomzq5cQ/5m08DjQG975VHS4hnp2GTA
bdNOMgDG0RpFhb55iqnnvD7SK1uHn8JYO+UADHMfc4rjlpvRt5ICOqVfk5tbQwQ1JURrp4v9qvXx
Zkm7c7sbmmtSYcKYbBHPDTR4F/gAYX9VpFQAjVxW1+1w75atHt6QNxUNz515zoWRb/zMnMicQwQl
3aymDO4jz3FD97ak37OQc5cUEeQV6rB+8nNDJ+sm5rTeyd8MhIdWs8VduQDNP9Y0EhcFO4kPbkLP
D67DAJ7kBwbniMKEQRTciQi59gcen/x60liURnxy1hwQ1FGd9YL+4C5kl04Dnt17nVxaZA4R8Q+3
HNt8fMLP+fAY7d7u5L7/fW/t0MjDl57c6QoY1fZu9dhcXBQ7rTTHCgm11vGVoqVUW2tqKSMNdD0q
w8y8dbetvsT942VYRKamZSQfRsSIx7baboWob2alchDWfX/+ZsGNUeJufpI8rcwRMwrh2J/4LIsL
j/O8gvuoIZFIxqCbPcCtVUfvg97yti3uWWOvKq3NTAOSbW+l69nFGfm+yo3oEyjk19Rt9SvgD6b6
Yfu7pD1Y927ypGIzfKzlBGj2/aiblAGwVAXpdvBQVtxrQypSlfCWZvRrx1dV0lZXmoL/4HeO8KBg
gH7r9iU7PyjPciAGF4d6CwS/3FdOhruU2p0r6j737UuayRYYSMVP1HFWz7aNuAoFoFMbSFDuzQVG
XeQN6oKxG/7C4Aq1huat/Yb0azfs4rDn5a6CRJsY1Tuysi7QLDg3dIpTptHKyFHklF07NHYMG69s
oui0enPaWD1aPQsfU20B/1HHdBHyNsB+G79r1nFeGl956Wt+XH+uzUcnSaDOM30RIINYS0IOuM+o
bUsinyAqaHsv4Pm4jZn1ELlEMtDliB1G5ucw864gKNj6YOKU0KZWAhRtylAkZrmGIjIQGAEV/fco
ti1YfUhOuYG6c+WoV76dojDX1nt0eKf/mTfDkCaLUx8wH9OSkyDjitSueURp64jkdtjqFzFUBjxG
yqbHMtLi27QthITutgEk4sUhupZ8IHiLY7p8yXWsjJ2grhmRVM4uaLNQIP9gocKPd8g/xC6FgN68
cyMez2uqAB/7EkB7WjB9s4leGXgVqmssPsKXnnqD71BpxM03ZbkxoBjCSXRxQUXcP3TarR4cPU0u
R5eFNYmcK20wjXCWAW6frTRXz4bpeFhyfweM0mAkcjN4urmG1nv7iOcuWFxE1QQk554tBxYyru9n
34lmrm/GbJTwP/ed6O+Jln/UYuY/KwBZ9HK92r/M21ZQfPtS8f5qKJ8GnTM4UKTIDOelc7529hu4
QeiMc+YXIHDQ0zpfj6oZstniAfWCQuKVR1mQG5xDaude8NQtXouWR1y+Pm8+UW4/HT2Y2MFabr2B
7Kq5kBk/fgzgYXsS/pAoXVTxwDE8Rg9XA7+2ph5sSQegUx90EqbiIfG4E5ODdRO3hXCkoW/mcsQY
ZAPDdv9EO55tnmaXQKanScJGS4G4pLbe6bVLdY4jMul8cozeak7cee913iRbPMBWlJJVnjr/wrR2
w2UN/ZF4b6BEw9OOW3Qmn1Qj2/IK1ex/CtpxIxhJM+jDvN9ynRpUXmcW6bSqlHNqt+l3g7qI3K8t
MYafm5MmzUnVhdAPI/0u1rekrVO/yxiVcGfH6ePsLPWfg6Y+GdSZytHqf8+h67yUigJpDSrEQpIV
5UcXDUPZxPoUAVy4+CKAiPgyU4Few4hT/v+JxQYj+W+V5ljQJjhX0+d+JRifoWd/5o0st9ykHUR2
cFImozxAHjb5cUaX5ZilEQ5vteLJEMFav4TcPqY9Q5htHUmx2Gd3k70DIAgFtUGmdHp4AFfpEE9r
z44qCZANTYMTIxC8EQYDtIxEYD96muvKBCjJXHqZuqmrnm2qQkE4Fcxf6LeZHRU29ZrE+Oh/Y4Lb
PN+QpDjYJ/p500oDI409yE4ZVOu1Hqogh877y1XF9uP98BWSGbmJOqoWVOvSOBWalMOTMcnzVuOl
f1x5oAe2yfF0n8FagGwPUtZ5GmQMishHlunVFM3MPQH7it/7xvnCMggnPhDoXLBu/nMGEb5V/BOc
caVHvqcMtbIt9baX1g0NTfWs/FwOxggACz1lQ1fnPQ1jF82ADACNv6omtxpFA8jRnKIHDSuphAM1
EMpbpjUJZLtzy8j4WCT34EM8F8eeaw68mHTeUQpwGzKdOcqWTf+ROu51C9V532j6Vv1yO1qd5nmf
sv/Glm+3ICzbOMW+//xEh3Gr+FlK05xcbKKHRE1lhRLIkmoC/GRVkOEPTi+wKxOVwFwEPL39b/zb
8igx2PEnV8tETf8AsV59vNomWosmhG2q3pmyk1HYAIyYl6EhaSNT32m3bPpX1LnFrNTKeVPYSqRU
oqGkZ4cwF21T20vaNJqwzYwbzoYTAxDMUsKq4xa8IvbWCW4nwmEjcrfjJWl3uX117kWU77iFtA1H
GwYeQ0Ef0ocAgZUO/YKHfhlnsQ9Qll2/3in1nBwCG/nF/OHAw9W4lFxXYp5vkbQjjQVOLvdCkVNS
wYDv1jtsV6Dtzf7uhKSXzIa9POuamFmkEq9gtvq6tXfZT2vzcoGLhK1+9h5DCSAB0mdzpfZsiPRd
Enjku6GnWM5KY/9JHgHJOyVWhHCHiqOX8xdXS6OmxjSmbj4Bfikn3z4+0vzcNmQQSfuWvmyRi/e4
SW8uIAvbKPPnO8uXolzwOETAgWuZK5n3GIbiAN+p6Xdk9N92GYnwKGN3qsayBL983OBO3XEn/zvS
wM/FWnVZtEyocEOBv6Af7mCI5UkQUrjmB4syUHFRO9HCY+Dx8K73tM0PZrB3QDDNDFBOd7qPBCoC
Dy1nDRA3B2rLqnewrnFKOFjMBu+HNNCZWjaV5G8hTbhbR1FVXSiABZJi2LfMuZoWdoorYG9K7Nq1
79RcAPosBzSaywj5tBK7Jemj2cTdxT9WjC0X1R5nUGcig1Xo2PLA1aWUtK/cjGx5sUYBLtzt5rQ3
M7klOPyXS5wgvyUOn5l9EoZ81sdn5DetTF7OWLdcqmODZtI4KMvmYcLeOiF+MfehvO5LJ20PoKaY
2kkQiRxqJwg8JkSPGvOIbPCWHuHDj0cOrDxr23TBO5wLeJXsR4qMf2DpzcpNUXAx17qpFoeCzRug
Swe7CkN4unUTcEbUOJ703pUNSzrrIAMqb4+YX5zHQ0Vgx0/GQeJxW78XFKmY3wLo34XBdO1jD1Rn
gUmRJqpLa7CRHZiiJJ3dlAeLDaQGGb6dCNmW6JZSOIf+d8JPulKPVgiMG6AnkeLbYcsPhbWIrDyj
2Z3QJ94lLEth0RRDLVOq8AWG8yYQ+k8QPjduQBSHfrSaO5HoLLendEd5NjORQMMpRkZz4ybPaKFB
SST86uYPDLEmw/7GxYM/SSN1aHC3TfWg2Z9Gxa5qtxfghKokVN7wLOVYt6KxC7hvInK4k1XN0io/
aV4Nrl+kFx3PHRE2k0r5rHRQkVvlju3hiCxCtJapzcab+AzAdDEkFZsTl5+7mbBbU4O8dyOq+rFH
1vvxOtQCc8LLRuQPVI2OS1x0W4entT0AUZxWwnV5Ycbon9Vz9vjdyaTvUJYQlzf8AoSj0raaaB5J
DAIA+t0aHOLhTE5OGHJLabXJY+2dPrbwcFpCbrWlJ/7NsfQA3YQpwAgeCVTQo+MZlOE1akvkTXgf
eA6b9AsVXfEMmmhxYjn4+Vj4hmmwd7hNibom3ySvYJZdWkFzyh2MkZQZRxFv/jp6/5B/2pHksVBe
CgXMGZTya18XatH/7zf0LVW0UfNZ2dBcO6KtVoJq/zOoU3ijE42D6M+txAozZfhmUXtn6jCuJ1wc
+XiYKhCsLobm2sOXSoU2yx6B85Hep3I66aVDxuNEoOom4Oqorpi3uxQJx717RqgY/l171HMj7SiD
deig1hpbA8ca17eH4nFhnV3flez7seP/AOHKaQvrkchKkroKI81f7e5sSnmR65DfpVWnfPJiKyCq
JRQrg0SIXLtCQFKwWmgopijfI5CU4IAWNnuvBIIQO/qkrAXcYjZ5fYa82ni3vTPxSs3fto4oxFHF
7yymdNMih2BPYNZxO8q2mkxCWM+2uTmvmI63/oYhTJXogqv5n7RxqZ1aUIqs8KFJCpZSJUsA0XAy
zF/TFD/oIk7Z6pQITHf5hu0wKJW9gZtfmjuFG4A+Vdkt4vTkkzt5fbPIPV8ZSUxDicMDPW6ETdLw
H5wV+L3/h06Lq0xsbmgu1miJ9F3Z+0rz0f59+ssE8FWvyf4x/r56xuxByVekHrCISsXmh9P1HCMO
Ax0/S7VuN5FCIajVimnkXYUAVI0kIadGrtJsG8RZE2xcdqc0aaDvVL3BXEn8eP7l7NPibrMRkIJj
mSxcZrVWoX3Cmk6wSflg7yCZx4bzyws44FQKvxXVda5dPfDUzB44aZwI1fKjTxzzFZbFoB7dIohk
Pqp0vNvHEdJUx9/0Oo0RuPSoKf75z90L4I2Dg5kiuRUQYbh/lx1AKeCfiCZRPoz2GRUK+JiHzZsS
bAe/O3OYGNgF60FnHW0RN0ZAzOcrVLqKkPRxM50REC23CEQJNT5dlnJfQ/oG91mD7VDIpTgNa1oY
Q8pA4T8p7pxeWGR7IWTSfFGPEMxIfjMRwgJfXF/sZpsBPGUm0B2H3SdElIxWj/1ZlcBm8J2jqECx
CzhmygiR2KVIKuyf2EA1GMKEfn06CxjS9lAzOXSyYOfAbhhZQTchHp4lRywe9e9Z2oLVQNPvVarr
Tu3E45gk7hK+mB2W7EbZnLG4sM1n/MTwIG6WOSX8/hfEk3NA9wgNWi3qBcZqw7kHeI9npU+N38ae
fJj14JYzdrcoaq7ZMlCHUjDWss5D24I1zT3tbJB8Kt0uqhXhU4+5l9T/MlLAJx1bF6LFJygel9VU
Xenb9UCLXQ1JLGiK8ub1BdKjySLNqE+V9ZecR+bQ7CYqcTIJVHA2Esq46cmkd70WOvOwYmJeAPQc
CJDeWqzs2JC3h42LY1a0Lhrh/y/2kRkR7doqTrLPMpWYyyvNluOpeJJHu/N9n10VeNkymLvscqsw
I1aE4YejY89+VhlVgwzcedWNxa30Sb3nT+0Na/FvUkV+qXHYXpRbDM/9tX36IAy1+//GyLfslaxe
jUtmnscAi+Aoj3GvvWIa4nx9DXnyec3tbrJuhGpZU+N8CepoZk5fFsSEsS6s9nHd+IehmqRAkgL/
ccweqvTaWeR6xVgcglQVz4Kma7GVQSyZ3QkxaPAWMnlv8zIRgUibTxJAMAP/F9QsQvyL9TaVwc4i
cW9Rd2fCHaTGEE9BotDEYVX//n10NUz7r+5j7r2+M1v1i/ZUNlADTu4g6DWqOxj/r7jkC14saGVg
aKhWzsdqwSDFibKHGNBkIDR47WJA/o7e3jUeOhCZzW13FubiyL+D3x30KRN4eJEShMs7ZY1XUg5q
nKNV4rdAL3mt/Mexk8ryiHuk6V5ONpQJjPfHEpEH2GIcnxvgI5M0tNE5f8kzRLaB7di7Tu0/SqbG
k/Gg847D5WNqIRKhZHegE2mQYFyUryMddyY4xbLMcsM0G4wdGUf8j3sUSYyzK5pwK9JlzCtlbGG9
36ZJh4pow81b/7smBG9JGtlRiEABCXVxgTgc3YKy4yPy9epkhFwACOpzLY4LDVZsVwtjxhH65gkY
65nDnp0G0sDYdYeb9Q6dtd1p40qD4hNCM563ZRqXKqPcUduZGFdhMA8x6QkbC8zyBmKPDndST330
551NfXYM7U3be8tTub3fAETe7GdWhoDvdm9gzC9EhvuZ7DqTw6FJ87rmQLC6v9Bmq1lRqDYtjhvU
RBRny2HSD9ea/wSVMy63VLrUdsnEmCmM4f13KinTjSNj0VSdCsEmqt6V/2iRE0AvwvSxMPWGFDy4
uHECuOczr5F+gPdrFjO9T81sQLA3Q/SJwkR1b/DGZ/79CrPO3zipffgnh8phLaQUkkhLNyedcIa1
ZZYZL4NoECXNDcOx7JSd/vrRZKaceKYiz1d+J1yl7hQzVeLpL14GWpnO+QVOuPZ3lurQjv4o5CEa
ZzAIokf9Q4Sn/9HBdwAU26Kr/AQBv9YkY0ubrVCOvXs++qOHRCO64+etTVlRXZ8JAWQsfI8jZaNw
lDnKp14o1XNb88NKHF4wc481ZuMEy67/kISVJNCnpbPiwWv+TjPQf02nj8V/7+enb7+qf+fiCbl+
mfDD6p88Ld1f/V7/0ROdLj6SGC6PBwe3N8ACDBP238LFg5d+DEhpv53qvLe0vdLxKllSHdtcVlSL
9EyaOhD3de7cbLQphm7qiugoNaIOyx/O54zhntMsJe+YXjc0t/DGe1+Kyh7dH+/13t0gEG7sqjoz
szQ48Y8WDshy9f5gF7fIi3RwvT16SFHyFIrnJqRMmQ7oZpX9CsVI40CmoTkdGKl1DrVI1P2fMqcp
uUMdUP3moIF6TIZCoQxTj697SLQ8CNnk7q1KkDpHwVgwNgz+KExEzn0wnF637+zaD2F1h2TV9lYb
n8NhimNwGIuRspgKfruibk5tqj0WjjXs3inO6jZ/P/Mr5XHABHLXqpyJQTUcxzflYRpq7bTIjK9Q
EUfAaX/5SZKfFp7RwGjUnJvyx5tewGgTmFSjY/dyxvxn9D4zgIVE7g4bR6emdzfEUEVUTKrwcX+R
oH3FJ3wSuy7stlxdwLJilfff1adV7GXN9Gzk/NU2UwBRjfnTx3bwkBm9RGefqFsDyqMdqKcQ6Zub
+5zr9+ZvhWi4yvrcGBM+nwLGa7qGw8pMYNfJGBN+O/Vs68EWek7Ae9LcFJUyfotTtCWBnuPpuUFx
tzV8spM3PlaMg2OrxFeeaW4RFFm1+eT/FHronbMoXqfqZowpsFyDmIFm8EHn7YZQvaZezN4mSDNR
n1KWmI8a4JRt4tVP9dDYJ24YNLfns0zvN6h1L0TqU5cmfH6/jhAyuvhVZwD8F+1/REbkGLuhhlpR
QKzIGiKFD6ssN3dxkc9fliZoArEfLVLGAPMOrfGlKoewJCyz8TJaDQCS3DJzskR3NWCCKmQ1Y/OL
3VkfRDMOy6Vl5xlfS+r9UoRqa042YDhJYzkc9BBYT34VI1GWm31HmMSkx8viFx/8Z70m0aw+TQ4l
gRmolH6hW0oKfb3/JqcaJYkQzuheMmZAfdMRuVlsmcwq8HQAGzsLJHQGadyM+8Fi+DCKF89v6FiY
ZnATeKSZyywpUJIYdXwkxiLz7FSPP62xo0/o1UvAWkRqfmjFHiLxGKy3CzPo+UFBi/so9z8sVOCH
GllTNt6l6sbR3D9+3hyAmHS5t5ajrIOVkHbH4CSvE7mycnjcJk+d48doDCmZhRZtE4SvFLZ9JHSX
4/1SyTGlzq/O5R+PWolxekRl3NLkuY7a2CwvCCHx0kK2q8fgqPU+YyxzkxtA4CSWll1AdTvA9G2+
hcvB7gDchicAKOmavLVuuI+Tuf+LdBwMtW8fZcogGAKJLcvjEenq/iVs3wY4Ifer+NpzuOeAYro9
F/7C1XrlH2eUFP/TWijZOXFOOdmrRS1cuZkfbDVaSThCIRlUnanGEcH0BSChL1czeWrzS0N2UbDY
z9fguUCCPZqjsIvVi9YQXUfxAqWtrVUAjCS9qb9bR+MDgybqgrMuXOc42EGguOywdM5OgoqHVvTg
VVqSalrKahXVaY8btpVM5QFXuYSUvFkeetEhQNaoIE05nM5rB6XxeLA6TMvV6QYkXTnBPDDmAkdd
bBDgSpBvQFd7wRP30dS5D9JeRWzSbVfZgJ7yes90EoA8496wGQYTlA+DdgzyFubQpOJSunXorAnP
ND3VTPz5lamEnJLa6cCnprPUirmDVroKdrH0JLVZwbM7mFEKaMLX25l68PuH+W+LcENl/osp0gOu
dKb9TfG1loFlcvBp8ws242K2jrVC+THgWeoA+2o1pR2lYjrgWFH6m9rf89GqXc/N0xM4nwCFAb2o
5rfPTmouXox33wzEOBvt0wcXzFHMqaM2qCyNr1lCy5zPKUkCOuJMsqJN0Jy6bIvL675P3n5mu34E
JzWhhD9J3FWllEUlXIreAOb2Uv4jhfBSFEe+vcIFxYjHvXWwhuA8KZRQ9ZGkR9mCtoVFPzuK6RGL
WtU/BWhVUW2TF5FkigNJwFLq+cosf3jycBXqLNfRb+zHO+JOHCzXDT8xDLa4pfa5q7ogxstvYKQm
gcc53bILf9s7ZmaXJloxA1VjBlAWakVSxVTo/K1eZ589Bka0O1O6MNQK+uzQjqM8UsER3Q3djX03
d2AAoqlgJn4JNbNKJkTAjmoVT8JIeRDEtOFumKZbJWr4pVDtlcJ/7fDDEvOXYGUOebxbjJAAPekv
GHeh0CXn2NdssKW6EmM1JFqqkgSxnqXgh+PvnQ6rvYnuJq2Svoxekapid144b//Lw9APtKqZlUkk
bCyq0tRipinkjigRRHXB+AXKakJbcrUXQqxt6wFWwPgTEGeMkRbsrXK+7pjD488j2EhVfM8PeFMc
U0B/UfhcF5qQLX9mUX9g5/Y4G6fpY2k7xk4r/fbV0PK8XwO+IzQOaFURO68ODncvLfwYIzaBwUrC
PDA0A1b5rY8KIeqilnr8555G+XgrVGItHTjBQmX5CeOawigN2IqCjd42vu7pykNFJSfYjoWEU4+e
+N4okx67y/6JFRManr9WDDLe5MCIxSH2VTK0Mbd1U8ea5Hxxtn8zkg+IBYimgF28bNjWYrAOn5ms
hktoFanjuE2Af4HyVEW8NUVeMz4TRAjLr6DNYSCKCptHBvRj7vvOfnrtDbHJY+kMAR2MIDU6w1oW
C73Kxi7JQ5COcSS15OYZwnHDwqIk7LdVhWSg/YTte6rkJTrrgUAHFBzyxLSwM9snD82v4wkfZxKv
rBrW7Hm1XLYupW2+4ceNRrBc4lYJ2T1iOaW2iBfRdu9i7n1xXxQu/2p5NintPbL5HwbNPdeLVgBI
fozn8FD7amHahjrqfMO0x74/OfbmXsYzlfO6OvEayyqMdgw2fdbt0uBY3UY+nvOgPG8rwRVj0DZE
zBbcNGVfZIZdKiLaZ/VVWLtn2F2mZM+T/Y3gq9RHHL1magnsJGZafg8hw9BfeGmH+WDqHJmceHpf
yW4KfFU54n6zL1c4imbfB/o1k1gLitQDbcHadhVxMxAAx1lemeM7H3uvmB3G8wq+TYzEUNcpq75E
5b/vCDyLpepfpr9jfox2gMWXejuOTohZ91Xt1GeHU/Y2eT83Cs5rNjjyjuPcYQa5n2yrjYJEkcKn
xWU3XdbPsfRK9UYVTy3Dtppic5wbTFB+hLVagyS1FNd/WPheJVZdGnWxeC6gigncRtw/nAfcaDuz
tkYGhgPSiKiUXSmPxqXSclnfitugPoIDWOyTKutG7fLzdc68KzTGZDt8Zkv9F8WctyTgIuiwg+aF
NgocjZnADGZnTNB4wk2SyVcJMJXJnCKISv0nqLD4q8W08U8ATRe/D1sjq+qb5B2VHmx8CIluEeBI
wx/G8d3b4eIbE0/Yxb4yl2yhQkEFz5PhkYqR3hJnOuA9ZzLBlR8kdLYMtwy/WZSk/Bf8O6hZl5Ag
KpLfD4KcxT2m2+yLMmZDFf3DB8BJRXKeF5JrW+mDGscMaDW0f+Fho9l0GyA1U5PlZNHa/9932PYW
Ut2n0evKhNzTHlBL91AWeLTKZrPqkArxzXcgnc8JbaEnlQ7HzgA2DOag7yP+TdFM11xI7ojlvkLh
08RLpfBGJLzKGSnx84UCo5V8pZpHGWP5yumX6hZ3qQ4sXQSqN/LqgA8jN5UOr596loz8/xK9OcaF
wthdoflnigCVbq0gDgWSbf5yoI7yON1V6pLpjF0FH0uRDqHP8TxddvZPkdT5fuuz+oeiy3OfgKjR
59LrfqaNjgYRgc6fW9sUpOs4FUH9AognRuzQZtV7Im/cJVidv6NEk1GmiYuXIFSOh7ZR7ZS9Q84H
FmYlh2Z7xOgeNFyOkH3hxBYP1O5vJqD4ubc5ypDjgTeXafxNhA6fsmTCziA3gCkW724IaxBt+bxT
4moMUQ6YrZGk6IF+lMOPE17jlEWSN4amNlENvaGWRkBhQC6vX8WVd5J+81I4JFUPFz9Q1eIjJSa7
mZ/2V1Lo/7HH4wPKF6IsY8dOr81dTK82KkR3hsCNHfR10qRmWdvKNxIWvfZGl/belHR+bZR0tmvs
DQDTafGSp6ZBYAioKEaGDxeX2D7quc/OEAJKytuXTIJmyt8OLQymVT771hboKJ25SP/+0EHjkd4I
ROkvlcv4VJw2zrHsBpa/T27Wz18nALDB00PYw34WQSy4VLUbwA2poONGKqIa9bbNlJYlm9CCUhDU
dPafHCfLEsy/nFRwE+sGd906jzHlEpliK7w0jrjTgeQL6hBMlh7N7lxX1tSBjxSy3xbHa0HnCJp+
EEP/vXr3/K5w3vxg34UdBeo9HClNoVkmjqbJlnX/nDoSHxCdqYIFAP42EqsmasijXx5YXFjfjV9a
leiI96O9v/8QaOaSRRghUVNm7lUPopIaO0RVKRDZ91yqZUPwhL167wpsxcH6C2lwonCzIEokpEGS
TPY3SZ9JAm7KtJV29IRt//drdmHi9Z5VNap3bQEP7j3VAjSx/JotcCJrqyHzMdsP5j+PpKNSV/4q
Jdl4Qi7Vc0Z71X+KZdOzohhEQQNqy3QWNL0gZBMmE7f9MuZ842xMV+7s1Pzrk6+QxF728GuZaOuA
QN2FMLUjyorIlxVuhr4FtxIqdPJ/GlD1nIjLYXQupZ6kYBUWIvsl8g7I01yXsshC+QQRPwsAqfvZ
seQNOAkdyrdHyYgQPqUTe/UY9gy+8WZdtUAusQ+Tp2Kq6eCwMHoJOMUkPUDQ1cPwae+AW4+ZNKIw
HEgg5mItRj6pODQdrOfWwcbZ1e6xF/nbYER4qsKNWpwjt9sGikD0AQhAbOGWDjnbdwaF9Gki0zDX
TV4qHJpw1/esUFiSfSKtiILOzqpUx3Orv3qnsKlEE1N/NayvIGa165+B/pJEjSU0NdAZUYOhuwi2
T/cdpdmyFKvhNNpFUOcp516m2w1UmKSfB7wd0QzJrZSfiCgPXLrRD60Ks1H+g98JB05AEm+nAoEv
08jHJG8Rla63cTzE53bxe7jBCViuIfxmQ9gbuGOhqQcLrbBaBSErjhw8PHCalor71JjXtzARzVj5
xkSLJlcmj722HjwUNqNpBJ3W2SjD1LhUe7UF6w2s3Ql467lp1QS9+7QTPh7/u9XGCo5AoNRenhl2
A9HGFltV8EHUjSjMKOAOKAqU8zIhekCIBbwt/29VrPwuBO2VqYdzvWzeIIWQL2Sj3wnk6vvTfC/c
NUKNTZHBYmNIvpX/yg+4FRWE/DCwkicH8cCCDZ7oPie59KQVUV+7iIRVisShOVSMHLv3dChD7qVB
jCkZjS5lYM+WTMxBxnPUzM90XbVp1Aiq2sn1I1LL/IpY2NOHoOcsT7cecYrYIy8Cm5P8ZmrPfI6l
GFFlWi1qnxD82PV85UddSzjc15fNXnU+L4/whPVjrggD7D5XZ8f7nYoajhfHR3ux5F0gSjS7u2xZ
Ac2ekGuWMNmapohe8gn7WHKR/eNWiLEdG7sujZn5Kz/u7ojTTCHOdn7b+mnjDCBHSXY++gm/OGYr
7ni3dZwSxyT022/9y54M6KM5LCzVIGS1yEVmFpw2pD3bUoXPv/0ZP4OIi8ovdq1kgquX6XEv7W2K
4OTYL20EnNfosX1WtpYMhwAaSbF2euOkMBQtS5WCK2guxWkfKoXGwI52lN5aqr4JrmjudeRNszgB
bqoJweucSFxGFpM8TYae20qtXcW0wDF3mQAcLAu684ZdmL9/m3rbyvPZDw3G78nx4f87TZf98fzt
HwxjdXgWtOtvTdLtx8PXe/t2g9CDu6tF6TGc69o0FzFc2OpqFIsJxCkodzWGN3hkljA1SM0VGk8N
GwV/eY56qgDoNFjqARjm47mAKz9xOsaq6DggSeUd+EvKqm2FexuOzl66EtNsQx4p8unJhLXTe1d0
WmGctYrAC8Y3Z4AEGnLJdB9xNRr8wcrPRD51799JZjWizT0WfCTsxh6hYDHupSWSQ3kb/1EN7BSL
1rCxQrW+67ehenABAz+rjncpMzG7Wr0JLn3yKKbrWMGLY80F2KSeVcl4ZBtj2tPJnG4yKxHVwOwd
XdzAko+LIX1KnCAQR/naHttZjVhfS9dnv3BLnG0G6ytRsOXL0yJNQHsS3Oyy4KSLiQeFT/2MyuJz
CbeeXlNCiP84ADO4YuZcCXdLkSFc/OBdPVEM4YIULaSQjayiYs4Im3zdoTQ3oWZ6+C8Izlm8z0g6
/t2e6mU+ism79MHfEvsus81zbDd+n5uJ/60BTMw7tyxIbxc8i3rrwWOC2zvWX8jI0K9IB2XmufbK
TeZS16/RDgHwW+6FsSS1ykxi9vOMAJR1LJLHCn5OSevzkfnKWMWLzsqLAc8g4++bQ/fi6x7KVZNo
rLig42OulnNCmhl3pOFM0WGfGjPrwv6K5iVTl/2B/g6LUPSsWBtECl51NWQw77kyAMPlWpTISe1k
88EVk7wGatwvCfsUfHe1z1ejQfLOFcrcXsHJOm9ky12mqH4lP3XNOAe/f9piCiMcSLJlW2uBsS1g
b+1u8q63B4wDahYpJ1K69kV657cjIyPVMudl0281rdgBHEopPCrC497cuMfP0bvYiEBKKmphzsBR
jJzz9ycR2mvf/lmcqlRuX1qsQFa4q+PCpAA9JBdDq8XcCnB0Zsl9eXSqVk9LUOtzMd4B8qCvo2/6
HWEwVLJhQ8vNj0rnZFbca7GoBEtacKO+ZcF4eNU/n6yaDfauxhHBzjizHqHkexssOVIwNp0gaEd3
8Fxl1soGgOBp24Po3TbZIE2T30MsxdCt1ka5TtEFiRWsS1vKvmAU0eiDUsJYYuFw4eBAQJ1FuTi/
JGK6j8K23udZqCbalyBplJNNXIglF1mt8zkGxbncchfzLV4yyf7fQi8OQ1dAICpfOWz1ykv+o7j/
FoKQt5VJick6DlScBhA4yPfxAEGxk2DXAC0My89xg1aDpYtJQwsMr/SHSf9JXesYJ+Ep/fTrUlAa
jnLuzbukMgXUoHYTeznr35ULJ7stwccKm6Fr3vCOZqbIFBTARdPKO1oxQlgBezcwdDMUcbt7k7Dn
H3ZIHEgbG/JkO/G1qCjeO4SNeJuTYs84lZmNee2/ZyKW+4BGkFZG89xTgHwBduhfk9v6RKNtdFfN
zVu9XbcW0Ura9iF3Ko2D+5KaX4hT2KzHkT//kxRoKxPlmppufeD97nl0zXlakLcOvTBZx/7hHDd5
l6BtycdepYSSnCwhaX+6TPvOLXCEEHp0VBVG3DOAF2X65Sh8qQ7G8Gtsr8Mlvc7NvKcDBuAc2ici
pMXW4J+zw2jKR52w4+hOPb2/yR1JUM1D0QHRG7cxkVPt8GfcY7lpVMz9I+dXWdZkHOWVQ9KdZ7PT
zt96QS5PxHCz7EMO/EOvxLngxgC1x3QSSvlklyTsu4OvLn1SeVNrwbvz/VVXGZ5W5PKW85dwPKVR
vU4eMgyDh/hacARyiyR/vZcUUeY19i0TRJ8NrmQ+RZNI9I3Ez47SXsKTVTjZAqWeLbcstfr9edJ4
mj8d8HGT+56nZn/LDPpb2ug9ZbkWfXznmryg+sfc9Oekt46yBg/m9K88vsCrSzBPtVj/DXVDXHMV
hLQCW51tLGDGiS77tdaGK/+65KC0LVGSZrDww9HW9UaiQ9WUp+AGfX1pApzHvwW2np2tcAa70ypF
AB0zF5+pUFI6skWngcMjG6NwD9dAYyjxzKTWGx01edhGvdzjwzX4Z8Q1cj9YB1wZuEwOAi9xSTnu
z6oqoVBzCO8YbWcF4SXofO8fxSFlbKoJBD3hc8YTsdbI3mQUVTISq52eF36HCEPdS2uS6xmmpb14
mGBFvLD9exhO8dh1JnNBCKR8GkeLMrIjunZl7DnRBWCKNOFsTaVrvT1qRVgrMwbm/nj86nKwO5SF
wqV3Do4tGwEQcWtakzsikextG7vYRn7ydFayDG4DzLx81JYiEmpaVQyCIsz14BrdjB0U1nY6IyXJ
OznX+SEDCm00WrMz5JX8NClCa7quRoLlI50X8H0Ljq55cZfMGYu/fLRloxFu6GUTyzPEB1FxpOaE
W6YhQRKFHKMlorhxfiQmoSmfoN0G7ttl/5v/i2Dn1EnfEe1f8cfDNR0IXxCNA4DO9kgZFXjv5kYc
HHHNUvFUoWX8bJIwCShPomot4CL+Ijq4clXTwVaDqKe3FgHuBchjYsZ0s9vl4bSRJbABniQo28kR
ewJZgwBgMYDvA0LeX5Nt0DkqcKd7agC/zSuQ+MhkDYsoywz2D8Zf96jdxq3iZMDPYqwK40g/qbuE
r+3BCWBNJ1LPTtlFdm07/mb3FJym/AAzq0nlkvwBoDt74/T0FGAoVjEmLCluW+DIeoWZN8YoKVeQ
yQ+BG5fQHLXgRKDHMb58sdoi1jXCei4xnpvv6nxI9wJq+vq67W29A5IrNo2SpAhxqlB8i/2waDPN
tOIS+gqhJPcQNZE3wEyRoi3ku3Fruw5r9bh7ulBrWaeMB3e/KpsTHLIdPbEJBCFcspomluZjDsKj
k/hgs6YeNy8MmnH8Ch2at2o4L7rgM/1RME/I+mzw1yzavc4bAJM8o+kQdTWjCi5CLZQMFcNgDrig
wr0ojgwUrTo6zisiBy46WII/OHmiQffeUDCzDOKInGO1NmlOC8pj9jRLmlwFu1v064qwphw/kdnq
CXD2fDAGBCswytg2qn9CzI704X1uf61euc3Hkq2oDuTmYe28uzok8SkjBawbhj/fwKM/L0YRmR1z
fnu+EpGk7xTJ08MUsxWV4+Buvc72QmVrxK/DsYOUDjUqjQOHnMCvbNix0OR+haPWmbOtMAVGGfi4
5XQdm0fIczwPmFRC0UZA4qdpLvRn3FaNod1De5l2UMHNsxMoozxOanV2vY0SzSVykg5BYOat6WJO
RPv0A4+5TL1vWYNe14L71DXo70z0GkeX42YmG/yy38UcDgo72PlagtfNIwIu5+l0zabSIrU2bi4j
hZosd6+BOde+MrpyZupiB5hm8F+UbF4oWtlXrdQMRfom1dQpei2uFg2YcQsYV0AgNZeaOmxkm3ga
qI8C6xYwRpnV6CSxhGfFho7o6hhCbsXRPN0iJHYGjvMOyPDBFkjI4DqL/b2OIRUXrW+zn+Y84feM
pepiqZqqdsqpJgE6S/3v6K3btjJ1dDmE3a2O41ZAf/2BjDihzdtXe75PYTnHFV+eCP7lrORWoVE2
ExdD4JHFSIm6zhaLj0wp7jx2Ic1I9vC997HMUPZBngbOCi7rElclwYTaDlfnzDrhJuU9asdKA3PM
fQBDSO/rIoJPLLlGj3s3y9euJu1H5nzK1jezbjphrtQXDzqqwWuwwksoub/qYQO5tgt9sPOhHr8E
xMe2BSHogOLAp/uprCzPpU9yR+33gP1TybHzApGpEY9a4xU4r56yjGIRvxn9ckfwut85WbYI1Sie
U/ui0ROGWAnh/uMmhLJGxatJEZ121K9Cf6RnunChiOy0DawaEyyqPAekXxqHdq0nChoywuNOUzVj
mmKlJESyQVgBYl5Yz3QfxvSfkGFMNKkdP+8wAZJh5bkshYeYffrZ9tENJG0JAtIPrXTzfW5ZkzwS
SQnsXQDlxtecUGrr8rmD3Pw88cY3F2v3i7miX9DmmQi4HZJzR/DGiPuSABhapGko9hqmw3Zje01J
y2gdMLintSAtbfzJP4GDHKvHMa4XauHdmvKZk38L4wSiFsuLqhyrQFxrhyJFN9VRBNHyELnBBQA7
ktjf0nZiytV89STD/hyXMPqfG1WrFqF05jywzqTemzDbGlC8aRydipCXmJoepGkorb3LsfW7TKz0
xPNJNDXP+7bwJccSBihGDZfK3jE7B+DLQBMhJfIIhC1g4aOQG5y+dP99OqZtjbBjuLEmXe7FWRJ3
cWglPHwfE6eJZyJFBxTyvG4vW8eJMXTB21a0kYevtcNjzucq1TinsHKb1/iWdHq20gxsrvJVT80U
JDZfI0HIE3SzvzjoTKWTFp2tgLtgd6u37oxp1ENQrzBQ0BrhItDVJzg9b2ZgImSf/YIBTqkB8iMU
Pq+jR4XOomdV/0taphAx4bFgMO61S/I+1HVk4leFQzuCFO4iFK0FkxeXhpz4Q+hLtekq0tcaV7m7
qe4XBpGblHxbPASTGhzEmhXDI8T2qKF7Mqey87dUgrqlkWlXM4TsMzRV7gKaUjghB9/OLhs8Llfh
B/5qb5Vgn37jVQg5XmHpym7WKr3vcJHWMce1EYpEtzivEzuyR8P/o2wk46XiSJDV5WalsEyRouQP
sSqJQGHRUCG6Xac+LMS60rc1N83pkKMe7XXto+8xx66xo/9VAVIlu8Nk9pzyTRmXZRt1tlvEdOwW
a6H8Wmd+7N4UugNVhdJoYMbC3vR96HZqz+ysxM1JS4hWkR3hkO+r+2UGHqr+d0n8YBNpX4+d1zdL
qfqEB14dXlgwRdgVarBp63yZUgA/ZtLXK2QLKHVqw34AWTqda/9a7YM//t+HEqKBLhl5l6o92rLB
nMyaHVz2sr9axKhmgDxMQ1YaNJfqPrk6jR5Qp46faCst+f3adfMv77L877uYVefsoP+GSHJ72s3d
eTl0jB0LEIE7YyXY30M6jSTy4ZZdapnmanLRi1p04TOsbgAr9laNMGbscFRusRjpage/o1X7A4tN
jDD607dPQt0VIiwf91eGV5c3x+5GijYQ51ERUTx7B/rpY9hlSfeLygdXw/VyZ9akl3VaTbGtmbzI
hA3hooROf/GXvX0ZZhlxghsY4B36k2T5JRd+GTPaa5DMuZ00Yv+NBXdlgG5nH3SVxfYgXsEpBGW2
hZWMfQWFqD/0iaE/2eQLqQ/oXMVSLL3RRs9pqCmFwtOGwI4+J+XccG+UCkeHNlosp3htYD8S7cjJ
iBD57DfFzZMoyBZKKqP0RtBLmTRRNeTyMMuzPbicKgch9kokQE+pEHU9wybsmrNzRvefdOqLSaci
ShsIHuMjmiNmRh9WmEwExn6o8G8Met0YS7xmnlBEy/R6tSpubc7VfphFHLz1ojfG2rIzfjQFb3lf
h3fd6HKwKDTSDW2Pr4LunmkNMhpraX8rrTreIaEoNEaR2IA6MDxDHdZvj9YKIxvK2TT4RE/ppS4L
VrmESJuIH+KxlrJ6PCD8G02cXonbjLSCxuqm1jPUY0SblSMEwmTb9+TOROoToYjFW+GTDh1mjXfI
C6DatgPmftbQcyJxdEAkD4T8BnYK6TM+6rFhtUQct9z8ZltP3wfA+qWmGB1oFspyHwhT7vJ1KJ27
FffymtvodfIjnmCqfo6cgDJ6ko4JvXo+0KXr5xGbKBRFVVTyZcuwq16jcEs/F4YhL6plhTaZjBdp
AHQ/kabACMG2BgUJwlKnQKspnCxSQRTHNjTloUTcg9neqjQ4VIjpF2os3kP23Y+Wf7rUtcz7nT9l
Jv1oZN6XznB3BBPhKZyp4FyjMSCHMtT9k71E/qgWyK24G9dL3oAF/W5WYViNqJ1EBzzn3MOc3zJA
8C4j3u+/Oscen73Myw7bkwIwys1Ic+/GZ00nfdMd8S28e8VwFpLg4gNW/WqDYDfAlgPQKNhb73VV
MLA0v0lTXVfEwyp+hUiDMk5cetNI9Pc7lqcz2/RSNh7ZBsx0GnVfAAVKk+wLfQTobxCfyLAdbiFo
RAp4Rl28i6qXVXomPqZ6uxHzUk49kgWkWDMxesvRetBfU/+78dNWA5jYDRc7msZtSLi2A0hKKknW
PP7XwjkUVg2j5EdO8Hjb0ztHHFN8u9t+K6o1k8Ju+vixdUnBuay2yykQLDdoP8Qrpb/JNd/RvA2y
1nX0dhsorA5/3jlHwnhBsl2SgYWZYxxxW0FlR7pVAxOTyqHZRyqKOmOHnFwzE4G5NOJsUpVqbM9D
MKa1dLaN6OVys51dFC2aqumExpMpoBOI+zTBhFE3wj96KL5ak/KRUNn9cRYRJwSYhX27RTnhWgru
L1Mcy6Zd583YYbh/Vwfhitu0b4ym6S80UxF0EmmnHbjW3DnGOcPEiu1oB3UZPzVEeOGqJxBP/5UY
gXCrCcCKGcDFwgAvGO3FNDpbibGOAIQKiMylpPKRDKQeC0dkU2ZR/XDVkWhsHY4JcErdrP1Efwjx
x251C2mZXvsqKFAkELrczkko7rPZ6/++LXsUBezNOuPazAL7h6vgzTwzxmzXcvT1gEFcRwHuUrKV
thYHiMGiNKm/IcrvC3HKkugWMe1uEcDRrI/zeS1O0jG9dsuLuP1gOFq7iqBmpYkcUQMHGDn2PNDv
odiWbNUOL/bBtKiPifyID6Cwv7xJkbOpRGZBpgl0r+4smtpb+TkUxHy7HKzz93ISEn93TQ08cb3j
Ae/Vo4JQI9rHy4nIEkJ/zsTSVZj2v6qxR77mZmRmJvrrqXAi4KKrFwTlZPCXPngb5dDUxu4ugtLp
qNIAtbbmOe9vlmfHQyQ6S/cJeomC2lqOxfkZiK3RHI6PBdtx1Tmk+o8O/9FaXs3U4ZX05G9B+COK
eqDu9ygS0WWqEAMx2Rm372mDjnnm1UkzpkBMIipJVTv4KbE9I0lYn2Wd4ZyvSV21TUsjCwTxvZxp
uCavcTXDTdwxoD2DmVRuCQIodLvx8eLynD/umX47kOvQ/RoFsIQxbKLgb9oxu9PMubuI/DQ+4GRC
cQbDC9HcUqO9xYN5Ci01WLVBRKnQM+9Sq9vD22DIzaXJNaYf5d9u8X9C6y7Ch9fN7LQ5xt7I7OnG
WXul1S/z+Iuax8OfURwIgkk2k6nmB+WvT6TXu+SrH+KcTiqTmz4V9pVnNEoWV8NDKi5akuGQoji7
06W7tYT85hCR8XSKRi1jBvtyHkeWoVedW/Nt1lLXbPwgz05NXVXYmKbRqF20PXHj3wxvHXnKzFZu
8nPcNXwz+FHD2hkymteWp1a7apym1Yx7M/CS+jA3v8gbD7SCFLrfOSeWl16mvCjrRWBRhIXbPPtj
gcJ+BCQPllJlJ1XvJ2O5DSa5dhH4ViWdMIO7woB47IKJRLMgbRvedP1VRn9PyQmH4s5NKL6/6adc
2P/5QtBX3ptV1ax6Jd2TmiR9VCtuEkhepx1iXHmtbxb5970kcV+t1tbtJ0pDWTBO+hQZ8EbVDkR5
MINuCUQutY5QEfDmzkWbBjA3HMC8IptBBr5uFmQnhQabsyqc/oJ/1qaaYZCTncYCE3XySSfNSYq6
3o7Ehzz5sV3OYJO4MykYT8JDM4/8ryRME4QiQ0454CPo89zkig0sdZh+8VKti4R7HW0UirCX1VTT
lRQX/7sYZLp7NALLfCi+srReYyEVkPcnDjB1jbDC4TwLO82d2gJS7f6+9dOGmfY2jlD7tsKbbOpz
qddUVcKkAkaup5ALPUKOB0xm5kVuyUQ+nkLpXg5dZi3X+Q16t+X35lLlKC1Cg5P3+YKP4FpfxUri
251/I86HdDzImDsQY9FIcdoo7GUekGvZP6xZy+JasFbvfj/UlAFjg3xw8WEZzlI5OmiFpSh+LtC8
oNN2yTz7H01cyuYHQvAkE7tdrG4gfRTLYWSeJk60Tk4ivrYU2cB/CedGEqQibefKrzSAULBqRyny
jsBlc4SCyyO02BRc0UgMpNtsOhSSUUs9WGOH9FrK5zyyjaKuKo8kj8p9lwBFIceTv8fi0S8EB/yK
JmyjrY8UyZWQSHKluqq+c14kfKYgSgh41erZQ8t8MwYnvS7nMAfKd0wmq/DQOcMy+IHgdUHQS4/V
0GJZMOxvBH+pD4HWYi1C4QG9lcIjM+ZQhy3aCPJrnLCGASpM88TsuOG311eFKPsN3D+eMKeTd1E5
8E9qv+Gh6/57fhtTf18ENm5e5QAR34+Pa+IYgEr+u8F90LjRGK2jrq7DeU4EodmNzwlbaVqRmeky
0XJkWK3vH3b9vvpuJZUDl/O9m/0nGRaySlCSUU4djQkyo8RKh4JpbC/PAZ1tg1WtbU2E1mwH/D9P
RkcU2E8A5+Gayd31IcBKBKQHfLdMQHRU712zn0XeQFBoGfA3UXkaSXCJbu/xhIV5I3ER+NjdfXqu
KzUm+XxtjgT5ltdWcm0THTFCvt8+QgeoYMjWv7Lb/vTO+VoHIWwLTKsh7fPYRbKeL0D5VmEsZuSy
AZ1luayU3cqgPn2vYOHQDrdNjml/jDAhBVmbmkvIDunW7+AAv+OYvWNzxoiPSIkTlys36zMBQ8SO
tN4y+l82UMljD3YqDuIH7etuIMw7hZkHaoMe8475dZb4itwY/c9EeCme/O8IBHLKRyVmzbnTXX6u
CD/Zx137Ny3Fu8MDDU8a/n2Ff24g5N+EVOks8HPlJiTbMjtfHr1H6urvXulSmqa8qwJlJrgoFCIU
yEtpFKxYEqr0zkDirjavulocBJgfuHwmhXVGwDgVlZ2XGrFZYj6ZqqYHNJ+hRb7hmzHBd8PwJtUt
CaCd8UNRMW7xomgiZFSOXdTlBh/mXwhLYfWkylmjuA5avT7UL5qIbWi45fGABnjWa4UlCRVIVqjx
Qptey+pR48Imt8gyswVcgCScjXEqJBamC4evBxWcwZyW2xpBWUHvkyr9JGlj9M/m8FNIBkqgIJSQ
XBFBBQ1lXX0kHFeKsSG4gbL/A4jQfERc4SvkS3k4DCTMTVRs57weoSRi+PFhr3kLaqsoWVUFXQpQ
wPJnpY2jvaREoS/oU9r9Pbo8UcE/KV9KjmY3Cwz7Bc0nJiY4jE5soCTutuTSxxLq66utQYuVgnIn
UpQfxxVj6G5ZIBjQ53lByjJVacOPD76bgda0cFQBRUokGSL7tXktUxQZtFYJJeQmHaw2YXVu0I7Q
1UWgYOepkHdueePipLYv6EZf0LiI5j7Ap6ox8xRkJJf2QJZpPCwUYdxj74KUrDzizLj9PfYM1Yix
sXRYcQd+X3orqEOtB6EfMgNrd/wFWHNAKuJX6NlLRxKgT2FIKevstP+kkUFiQA+3/Ca60mljBeZY
LVy6wIWlXkiqmI1J/TExmFs9hDbmk3oUrxmxYen9I64cr0Gh1jtWMO+xQX2iQglkH5L3baoQHpkY
pl7NkeZHF/o8HcKTcNULrXXTceivbV9N031gzVoi2ZhliX8KMfa58yUOzltE5/agnxZUTo+Mbquk
B6gNmeeWajEvM4ESQceVg6Pihy6YhBNaRCn9Idn7RTAgwAKjCR3NJgaUcwfONGy2dTXNF53y0rVQ
r/eDaiz8VZYVcVfbglYIamZmPfPsFDHvPNliq9DQoOpI7yvqsOInUiPEqVJoCm6IfzLnZyN+L8DG
LlVFD5sdUTB4wYSChXVUsTg+BrN0ibKU0Lec3DYCPrQSN0HQHhbwHG4N1L7uUErPcXTLwyG+dFqD
3mzonVr+gV6UEN+i5aYWUEVA3JpqBdUCxYgYidtSY9DHpynw6Uj4i0hCbeSQaDfdYRunlOQ9AaV+
V/AYl2KpzNxW0EJCDg91IufVp3Q0LjAbj4pgic674sSPaxK9qlaZRc9cKbD+2S54bIet7xfqYCKS
ZObgGQMNy2diQKmTX3cqIvIodGtvZ8KTtSmhEie3Y8ScLb/iuLDVGf4owQQTUFKAKiz+fASeHVm1
O7PeW1coKqpoLjoupJhP1lyjpBaapPoIBFfIsdkjyHTkK1aD1AHt/tFm9nBKQQgkmvh7Ch+sV9Jl
o9FfvbVkaSCC46W82ohon2+GFRbtyl7iaJWSESVAma5CUxgmLVg982N7hhwmuSK0+zoNJ3y/i9m8
ueu9F/wYnJGGrJAR/hCbGawTO4Bvvz3jEh0NUncbFyAxAldqAs8EtWUgbk3//zybrbzpqaC0QSrR
4ZrRZH9sSTShL9F9q/p1TJJBNx8uVGg1sRDywaC/9bwcCMdFVPJf32EDM4iIIsoorFMz6r78xZbx
9whXmBjhstreEYk/mt2XGj0aQpAhDeybBkrC3g2CqB45eB6f7OblPwQOGpX/HrN2I4Bs5GYKxEqk
OVYJkXNntVbTZyjcVRYZIgQ2nAK3MLXHR06Mqg/UlWc6ji9RjKcKBgijKz/nleEm2lp7DnsH1uqH
wq2ElXhhaEA/IKa4LJM8UyvmyOmEe/gk0Wftf0WYVI7jU/QSaawKhlnEhGxUtHSW8s/ViJ92vQHM
3VnJhsYTNt63jzYxjv78UnUAvkCHb6PaNJ4U04a7kkJYfnNsan+s08OCYlT/e720hZTQBcZeO2sc
rIl8eH7o+28Ec2Es32qIK4ucwbySEvhjjGgkJslQYWoHyvaE5QoRzv1r/tolEcdVT3Pw2jfXy5fu
3IREnEaKWxp+50kLgp7yTZQ71R3ToE49MjLtVTDuyHLwh74w7awDwQKuKIrYQFbS97nIBlp4On6W
bpAK0PNzBXJlRMX/hBbCbWvrm3wQ3zVLctTldB1ZsB6+lVXrAHX4e6AxF3QV6cb/6Y9n98sv7Rkt
LYHtDFAgkdub7yzhJoHjuL4MSNm8/WpcLEr/SUHArSR8l0hSd8+I32nRqKUnxf9pCrK7CA6Tx7N8
iA1fSFMtK16RFDeJgZ1apiGp2Bxj0KuqoMqeLfim5E0QakdW/medyRBvVX3KC8qw7mlXHb3rKvvs
NVZO3Jr7E1/tzvTzs6rZ/+WeNMKkyZaXqXWrFUVB/o8l9FfF5Kud+HvwVz50o8WA0UKa9VsDOSSI
oCVR88boJwllcPWKkx5CQSpC4cJxeDyzPBy6F/n+hircUjnpl+ECsfuwWRmNORTA/mzkvM6Qh3LM
cAIKalbYubXwkjEtl/WMS92R8G13mG5lO+/mtO17GJMyGSXTa5L2yeao7EEtski3PvGfovXBXLaP
v0TGqeYTadUUILz8puKDNGnkrVcX4j5zzUSRAxnCSYSoks8t7mAPjMFAa7gA2j30K/wQ5es/7/1E
ClEdJ5XCHC+1UPbkkeqWVpiRXpPpUFvtITt5ppN2+piKyOhRxA3Fv/wOiykhBl9wTnyEpDLfM83M
BHtTnOmicW2NsHzY5FLEoPYo7eX5ABqq+04VixXNNRzTTbvI2hzVeGEk0650VpaECDx3NSJYQrcG
OYqO+gwnsOVm0mThyrEXWAb2b7YLgkfFVC210gchAUtrZcPrWcICyBH2SrI+nltAkAMmC7Ern+Yh
ab0HhEF6xWM7x2B/VXsD0OyFXWzljfVizqZr0RHbL6YwcqlPIGOwMR+flys/fK6JUXPQ/XKqxIVd
8O9xItFt6rMTkp6iunMO3iIXXhDE+O9mwAkdvYRPE8Jn8KQhy3EciCvuDcSIJiA6Xj1R+l+HCC3v
bwrk41B9KELtpaccUKkdvb3KfvtW5FBcCDBwDWOfCU5n/28uu3/xeSvdPh9uilOeYwJIGikWo8/R
JDrvVWj8ctm+KJBa1Z7BF3DVMVYEe5L1CkGQ7t58cUgg2z4s2NCEfeErUwb075IaNDo7xt45ZJrJ
CMEEQwJ5lk84PMEFjKEaXyFFWNXfeCFHjy6sJ8ry2QB/rlBJ/YXRHPhDi6z7olbZ5E99JJSbQn3e
fVvXKhbAIHP/S0et6yG5LzdnjlkB6NrAjV4Q0YqwhY6GnYnuMz87A0K+HVp7DGe3o4bh28sUGPhN
+o3fcaVGfRUkdGjTWalaS3sUZanLZJ8Uf1RaaGT/72ikiRC96SKS+lhiykcbsZTH+XuzRF16nANZ
ah/1zgD1ln5Gq1bCMa6uIGS9bAXfaIvWJg61Dpjnxbs3WTWeaDdl/7wTydOhmabYewaVyZDyAKlW
XM8xJOgposZB8W+zcxLoK4u5te3b2EAevq9aUc03IRzkqSZywA4+SsB+lpjpY4Xc5MoLnMQpkuC+
XtrHaS91D6UnJucHtTVFNnHXYWdGu87vyCwD9Yh7NaQTLbjSdAufeomijJfCdFDlyFC/sr/IyHZX
dGJMzBuAEtCAItAtsxPSmr9QxmNKtxj4aL88wQqPpurQ8uT26UQFQmUt1cKU69EKZ/YgbPqg5z7u
mpZRHWvaTuBL7G1NMew9kWqSWZLijTlhbLcN55KIHe9R7S6IM9KlzxMOQegBwBJzcirifwP2wwK3
RLFHeibHdGY8xXmjRzEonRldFkzEMuvCRrSiWdJLuRzCCsKDydAN6Ku7lc7QzYaMn9yVksRbhyjQ
xtBq6ZcWXlVkG2sEFvMeroU8n8WvukKiNMWXJC7jfit0gGpfeSRHH8m9urUY+Fv/+LWnlwQqQJBV
FPB+TkdC+/MQEYZqs7Eq8Bc2wzfDMrT89qaij4LUDM0PdTt15IYdnCqe4W8Kq01/8G/MIIKgvmZX
hSVJeh7XTeInoa+myWDhWI8DwVoXsGvx8E3i4KogmUDUYb072wXODCo+GewULnB70zgMnBgGXu9J
RpflVoKXnezNp2pq3eaGCh1wi3lOQM+ZgnBz2O+0m+6TD/AVhfLPpIMohbgRy4IFLm8aiTlIpWBM
IrZ8vq+S6OGCA/0USvl5l73JyccQqfFZ6TAb3LyW5iYMxggaRf7yL1IhOHxIjW+yce5qM8YATgtq
UBVmz1zCP9awE6x0SYoeYNg3uE0dsQCw6uRLG87fPgHA+9l0lUBQtAi3koSf1CkDf2CNhMKDeup1
7awonEOwpDt14bSE41aLURStRZKI9B7TugsfMwMGa2vy4mhmQ5dRrJ0Yhn1kfYm5DVC7gnaG3v1m
NxQS24cFASruqFx4FUgPSwREG1JGSCLYY1TKzCeHYOx3I7qiwbn8vxRb5Moije902ky6x7FJ+nJu
aymvAkTFGwdS2T6IBuvrlz0U1qYXVtcTEqDx9r/+hygKPp/l30RTB+RqUmUtU3BD5it0vvF+9v12
yZcH31ihVKyeqI90nLFDa66Q6qBTBPVLEk9CWGlkHeOaboqqV/8fD1aVXi6qf2FvTil/YokOdOk6
gtTcw7vYltRLoA3LWMv0nHoCaT6N/CUrrx3IOKzWgJD7JL7gmJG6upm+uhgaNRhrcFL0HJs5A9tY
dreSMgbO3GPkE450DnJSDDjAfT6bOOLOctmW6S5NvSBjZrCaTMRkLOLAekFnapnsL4z2hnOtWBGq
ishA9KzAp0DAKAkfFS/FRhmOPnkOpWIcN47W5VG/KCoh2CT84XjgqYMmRnonIhXHVGPIeOK8uLd4
7ZgH2YVh8mKm5ef1JRNntzQJkuRKE7VbqfY31X0z0hSZGXxacYnq8ErDMW9/jyuqGTOdfDYqnrfO
Vb7/cQRO4MCaZAg0m+1UTPP8+MJKmKsxRWGAd4nTKUsxHbEdYaVocxqkTKYwWt6A0DarCNIbw9yS
A7FqQohvRY6P/36YhZPXqkvNS5eflFdI0tKT2G22/KWpXBWQ0dKeRcF8yVa9Ls19dvx2rLCcyLgO
WdxGVRmDprMZdVRL2TYbCLvEPaYYDK0rhmNgnF0Jqo981YxFzPJ+MVBqK1d+LzNGTy91pI6yp/9n
Wjk31SoQZC/fpPxDgzmar2Q6mKspnwWNzx0amLe4xNX/MtNVswS72JLoTaRLn6KOKljMkejlvwcV
qObiLKxv8eym9ftiQj6LoO6Tk1nykUfP/omkBJzZoyuBMy7Z9W3HCh8FuDgofGLXAjZes4BMqv+/
7j6Z+2DnaKgS7Us2FXWMp7ClpeNhU8BiriBxcDIlEG/AexPrGH8D3edjpn7k1HvmrQ+WlHvisNYy
NHDUycqQFeIuyLoJcjQLEI7zNUjFrd16LatJIpsguDIysUk4DWS4ts6zi0dpSZZXpEJwrDDATKDe
q6eRhfbWxlxWtpfG7AVF/v77qfcUcVPJ9ARm70ZnARiGWUrz+t/AG9k85ceP73MOqSwqbq8DuLB4
LhvVSDeDT2WSlfcvNE/kIHQlsOKqmt4vVW/X2gXxeurPR0UyMC+N+KyTu7YlAwtEB3xxv9QluLt9
2yCDtQBd7axX4QllhfwFjMVbpskwk+cfIMsibEhW47ErFqDXj7HIeCM/+ElZceFKGYrdUJyxHex1
eg4VV7rBjYiwo9eAQrqLILoIRPr8woe4yZEe7GkO+DctATHKcZKeay2ycqcOnVZGVKtZPqL46PSQ
OIH0zc6O6lx/Reltrxl2upATx/kG9vwoEtLBXJu5eplSPjlGsin1xw0I4vWFkSQr8LAUQXg1DtzY
UjLEfPrvYgH4yJw6fPb0cD8yr3D2dcSJ5JVt4GN3mz8QHY76J8FVQ/sCTRgg1gj/S+NlhwD9HfQa
JSD8KxLtVdvWrhJwJY5ZuwosOsTIN+Y1+U0ndYiwO235hkWJR4ZXBR8lOiqC5oi296bC4Kg+x7la
c16pUlXHtcmCFJssdUpNC5BzUJDuQt9jLOPXr1Mlh3H/iACgWzAz+408i2mU9NevjKaHHRuqwrqk
8MibF3N3WcMaqppnFrcZeCkDRQCAvDqrmc8iPXpKV1IRG8Ir9OkQ/5URlxIdk+wqe7Ey2Gtaj6dP
Z0Td99GYFnSeuD2jrY3knvDmmeRNqWvUh1CCZzWJsAx+EhYq8N9jYtQxMd82YrLFl9m505INNimF
d4bLX00DhnHIzLnBBmHgP6L2CzPW88F4FtjflsoKW9Mv4urAmaxRGVC/kpKfHLiccMwsLSHQvkHJ
H35bLnNKRs3xsK68sxfN+4DDD+4lj1QVrnhDZDMPIZcGElCxF0wIZX6NZizy71sKY8zzm5xRucWP
FoS/0nBBjOeoMRraGNeX1tEP1cPhR8OktfEy1D5rDxH3Y/+bARngqCHi/no3zHyJdGkWfRjxIbWa
5GMYtopPAIjT+EUQ4HKFmpUqvHj7G6NALHM3vmjojlBnQOVbfihFrJphQyMwuHTBVw+f4tFVsOnU
yhsEQHXSiIKN4DoUZrF3RTHVjc5aavPCalyd8PA3cZ8FJZL7c0QHQ8T2daIdqUXbYvqCHgvCoCaA
dm+uA8GY2yJe0et4izbruwfB63r3kVai3dbYAmcWHzzqhrbGKbUcKdnpBC3QHrEHiNdbxLYAF/r4
EIqsTJPNN/DdV1bt2OD23Qh0TGyo3vbdV7Yvs5UEnwx/qbEOQFcycK2IMhBCIjPC3MHdfeVccMRK
rTcFoR/ZhzMnTVLYcC/gafpbrnaESYvhbt83E1NYGVEhZwfvDhxFAJbaxGBw5Z/oiBuGvm4hx5i4
a1ONXFmsS47ihedgukcpzeqB9Cqbd3hrxZkzJIOa51lP5dQjhoyaHwZRa0jMLFc3CKvIdRMO1Vp3
18P2tqz3aymxHwnvUWRkRgVKijURACp6eCNIfdtAenSthEvynsCDKX42UTUfIB2GGl7SaYwUL2dv
00S3qnMaOQncOLMaQ+Z9DVvOP5pabrjblQ3P0QeUU9x0mbOv5BW6QDpBM0uu8DtDQfLL6F/m4mJM
zE1kr7XaklJj2SQ59SaUt4Hu4PsSC7NiB+ANYLnG7M+tvy/0kP/Q0HS/bqW7g/wnm4NMM6CMBaIN
BPWOPd5hfE+53vurf6x8UCgNeLMiQxGlxrZ+yh8V9lFGH0HnId/0h+LR81D5MgH0UOkgrPo3pJIz
iILMrEdEdpkCyCbaTzsS0+d78BHOsLJv/lG/+/qeMx/aPB7wTNcePGGIvbKgeyYp12ikeA65LEp0
pzFG2yNPg2XptcuG3FXGV0jsBBC1SQW7gwsyflZZWV2nQWvyjRSD++5ofBI6aJ4IsBajmm0NhjYw
objtTRGltMoiWiktt9IlPt6ZkAdoOhOs+h2QDZWfDk3BYFpmW55Zf//KHPmxtudrYZgcYt/1Dk6I
Z72ynK7TpLCbK6RdIpNyeVYg23BMzf5Czq6I8O6YLlXq4U46Z6lNEIhqXgELJPBvF8TqjlOF3NAg
KOAnk5kNl43e96u7Cid8qRgF/WFd7xedZkvt2Wi1eT9I7HOxrm5d62fwvWQWBEJEqXmz2iAUFz/D
xWXzTuiMpI1QA0SLFy2ng4lMZBvjuWlmZFFaGkEQApczHwqTEPWhbfoBRwcyk33sFzU+IVRVjP2p
IjKfjFEtWlFhKSSisWAJ8RLdIOzMwXGJx8YpqGNVo/bIadP08JtJIAqRG4a/So6DIz2YUGraDzMf
tLHzfuydttGe35gmTGcWyuvU/JixdHIk5IkYUBHC7OCgWF03SJ5k4O2/ezPZPgXLlj6aiieJArl+
tfXQ794YAqy7W1iFfUuu78RLniyE+UXLovNUol/MmrCeUC6DqTJ7jgWAhsphRlfUIGRhq9l2UlOC
4mm8srghVwuyBjUW+C1etglsfvxe/DEB16LugQaI/6JQpPi3FfsOgfiE7yfRMyXhinRszXCzr71o
iN97oPmXat5rjlTUcDTinkMZaCidCaxpQoKUylJtJhc47cn0dC+XiE1sba3WQq99XD6lnOZ8eFwY
7cwP34nnoI4QFnWUKh0el0QmwEPmrdG1+/whdJpYG+ZoZ1EkQhKZkxVIGEjbypyaCTwj12Q1yXeE
59xYZwm8NlWaqyNopUZmS9zpue4gvoW4EUZaFfiegdAX9K4AAVlnaxyFwyPeDDBPR8PRTOA/Iwse
rxlhXDByv7pZvywHVpIv5YNQiICSpRCfIVA/mKTeTOR0g8ZxWfAv9y1olSL4X6rv30iU0mk5i1My
OHIXxrzgyYe0d90kHuQ+pZLE3u01x6IfrE0Zq9aD0/6CPGrtc7kWZs/PuuFuENHs8pFsc2fJ45nD
V9gXxpptldKM7AfpvGyEL6WGbFcGFThXXDiD6KCUgTyQ+9uKfAxJcw9UhAPbesT/fTlaiiTF0RkN
mxMVbNczthb24FxCMDvfWMcxHopLe1hdAbx5n7EW5tv0rDsoIK3BJhwj1pnyl5H02xTK9Ta0Ljvk
9MjCw9LPFB9hwW9yEx9dgVZNwygaEw5NI0j8inv9HCE866MSz58h8xEJXMOu++8TeRMLj0iDdKSk
Qhvu2eJuJslactjm1Ia4Ncvo8CBvOf8cF3I+g2WivEtp0s+Xj0p6+UKptmgDaJQadIOnaBZ+T5iK
GhuL+WqpUV1j/7RSFQ3ZXVE4jj7np2BC5fKmy/YALy5BeMFMq1S46/6so8nF9Q+rAuBruUb11CQp
3M9KQ2STshajNtIQ5R3AIWTaLc5+s0I1S9qtkT0Z339mUp1DKr7QHD0/eXfZ4pr2J8O9er1/YNK5
hWn8aM9rgdi8/0IS0WztR6v49VGeuIlxZ9VkqtxZgu4z5RKL3D48OeLS11nwdfgA81JkmnUCO4EQ
1vMBEVtw6G1eo1+/sYGzsUWim2bI2TqnIwrAvaq2Fxfike/aWRifRDBEyansjUy2+N8oFHCkqY0w
E9nenlXfLPWZxV4l9nuM/tE+pVX0ZQE8RFRFupSb2JDqtMS6rk7uj5rh7JGdI6DiGE5F1z3bhZn1
jbKGsGK24HOhWKMZ8exFejZZBBS4p67j7yheMgrFxnzUSemriyOyYkNh5MN27I/1mBGLFtuFCWjG
ZN6RnfgFSP6YWfEgmjoMZcqNXH8PSIWoWIGkerttPHWM+cRobvyE5lqIaONiAI7bM7cU4U4Vihe9
Q7IW8JLbNvQixl03OqbVFaYo4R6P29bpZ1lc8kEg1xejdF43bBkQQfyde0jnWeX5yub2m9GbS08x
Z3z5iuM0RbLD3f/HGevtmiI7lazr1kV527Bj1JNsBTf0Fd2mzL77HT0TFVUAWiBSJauxdRPqGHGd
Lj+sZXyQ/nve42n8jY8vCvjK6txWfB7bmYWKMfVkkUmloiuqwBf9XaPucG1Zfry7hUVhqiyoixtd
PY3UYZhqk+pOzAXBYjmtZlLj9auFzAFGLM3+3lux7tAuiGYUmJqjCRgxFNhpyCK3eEmU1+3hFjDN
+3MIuF10gJm0hZ7dqoz5+MJRXjVUWwtOTDtgl2h2rlSQFijkDKlKHiX/T2SelQRZZXiDnydX8JeG
QzivV0fSYagwUW4MQS7yvu5hmHCPRc92G1eSGE9WGc4vT31ocS94astxO2JPR2jkvZSwrVG8sMty
G9NXlnPWaOtl/EcWLTwFe7BvtlvqSWUVy9+ly4PEaMKTXdzVW8STjx3PygWuGgZuZUsbwBYWZCH9
rJeB0Gz1Vh3EXEVmW6wSOoW9DZa7aR9PE61gcqORGwc2t7LaizZV0IhL0Io9USPueB8xJFXQ8b3K
AlTVidrfAIUgJPFXKA8jfkWYBblSj6IYLR+ZSH8snXcFsHd41r+MFyAzrUgENU+arzQgBD7I5lke
lIdVFQPvTzU89s9+V0Qxu+xg02+guPOivola4bdr8KWn06eoimwJ91LsByfI0EZ94zGgFIz830fX
HAR9RbW4BFFixYpug+49p0eEl3FIKGHmuYWcvREUBpAP4KUOAyk0G1vSId+KvU5c/vpTdpjmoU2t
DbU+HZuFHsrj37Qcp6E+v6rzmEBVCk0oraxH9uRo4Z6vKvbH/liFjYbtogmhfpFbPB3BIMztYNXm
QbqKQVeTERjdjHho2h8dYGDUMrpvrnVgS5Iap34uvfZycO8Z7h1f9Dcx71PK5/6lD8naBGF1YvaI
q8+uK9vNPjfPnq2hrJNFPMgOdzFHBAi8PZYBC/yEgPsrtIGOy/YOpvNwGkYh12rTFn1D93psp8LQ
nBCUX/539rP7HKmwYgG8CBl2VS52Z9IctZXPo86uXneYAfleKe4Q4VJ2dwsVLlYZ8xijBQnYtuPs
/8QikwFf8X1wU46U5Xk7ulXbbV5MYAbmD17I7IYjYAuaf0mjwYMf2z4OJRlHRQjdAvzqiCDijAbL
aNjmNdLhq3NuVQyog3nCczWT5Lxqiv2js8jPOEX28GBzN6xX+y6KpiDpqWzcJ9RBQpFmMTjKf6mC
kEinQRAIGmGXx8qbf31CFsJfjevF2QRdxQJFBMMI+JRdfdxaZImIoXxBBSWylH0cxoij0dF2gV9+
Rj40CPxVL6Vt7mpLr5GFZfYY6zavqyZGscL5K1NiurEh6ah9W1qN+lNbzOWHN7aE9oyMO+UtfZpa
ikddI7D4XCRJgVjqszzwt6Z8/4uXAgadhCFB3Qr/5TE1214leitQyphpFUXH3zCZiJoWS8NP/XLG
r/Y/z80Nbx/s/L15QHhZo3rccvK18lbp2h0juZZf21S1LOmizl9GAGubfWfeRneG1GD3ws2jkwKm
nJ6k3qxmy9keZ/pusRNl0GZG+B5zv1wlxU5e6zXfQ0hlH+laeatq+DrUcPXkxDASWummePyoR84e
8QsTOf2qbqw2fagXwHFcL0rodKLPOpQV5MaCFapGtYRP2IxWzL3Vmr1mBpaRD2Esl2BQosafTIaM
7b52cIluJ2QK5KM87jTIWxMGLAPJeSr3Yi7O+rqcK+a8zkUKs41JZXwleTMKaIEiou26U0Z9xzQv
+ECakPN+ijzJg0QeKWQi6g3XtH5nyVqKqw6GYWitS+2RlWshJ+yGaeamZHtjBldDIZ+owJ9vc7bn
47OZkMQ4WH3NcCAW46esw3K8U5m7ObYqIYOSUerhanB7RuRYF1Hc9RSNndfZB/y8iwF6GqFBgNql
tqRiIIf+h3NLj9OQvP/97y3da74mS4BFMGy2TuYvxrTpQuGTgYrdlsFu6Rh04rkW/WAcm0ERBd55
9wifhWWy2V2cIWUMDQ24AvEqfTeLeg0l+6Bj8cheqB+SJ5goVhIq5gEFZycu5NayDR0K+qyquoih
IAYQ06y310kGc6utXNiVCyHS0j97KCNPC/FMFrk3RjRlr5rRGiMTxtzgiFRqkgJavo05kXvkMfUU
7NSrHlwnIsBjYjtVg2WB9iI2+1DDcpY3RTyD1t6OhoIDBYMo4ptZODjHCYO0maiAiLq9zjS8sxNf
4xRvSwlvsbWdMeShRyTjZ1dArylFnUHFOrQwTdcdDRox1dxHMHnDhtOIREIjiBq9+eNSlJ5+KxgF
I+pyxZp49Si6X1/rss87BKhdCjo+17/FWknnCUocIYAOoyzEmCqGE8Hw58mqgZwuaFbQ1ia8civo
z2/XNMI1NSViB4aeiTisYq3ekNuzt2KSHC4E45osIIPPqMITV4wNX52ZT6DnXF1c2i57sgl8HG+Y
0MrIjxY8t1SlWbYK7MHMdGGMI/fws3DH+UvkdEndbfhdcv8rtf1itz4etZ1UxKW5h1PJXXISOnDE
JmKMxBhHocRfAPGf5MhLFxTL4LH7YSrCZyL6tDc1yK4CdPeyOYY9SB5y3GtUg79/hoGFqZju0b1D
McjRVCPxT9S74ktqo7prNTkvaEh1n/hBwXqzfaGpbye/5dRD+dn9osP9J1A8Td3LjcsGxKKdjZeo
Th7bbjZ6d8NssbHmMUftpQFjv645P0uXz0A9bSJrUZHG9qWvk49MEygjghZjl0eI8P3co98U4R1N
cC27NfczOtioF6ixquyjEQ8ssYeHUesIQJIoLB8Jw5Ys+dSjNqiYfvXCXvxz9zliMiL7d4gjwS6I
D5Y2X30cwb6/iaVKnnA120uTtPzEtfqSutNkkaLP4fUAD/WizyBXI/ud8/+Sc1OpBnZpHlOxiDxn
11ZcB4ErzPDYdTIYQpYUmXgc1Zr3DC/rwfk+77E+wjeY5XIKwQNSnvpPXclxFq4akt5w8DziOafP
8RYcF0yjB6MYct4GK9lX3lVpXWXMgVmrIJ16EbrlSk29Xz6V5OahmXQx5Mqi/PBUD4cUf4N/RIIj
hywzdXSrPQskUxsjTHddt5H+n3pOjjpdiO3FPkxwBuZinlIoP9W2A5Pz8wi2Lb1niBdwdcPg8LMN
lIPuA+V9wKz/ztak4KLqEmK3rAVNHW7m5b0cf8F1YTaIXlxGlUsxjluCQ51r3hYhPKN2S6JWn3kt
+xTRI+iEiAq74obopDrU1B6vrSL3KDfACsesjhkd3YplU2ULvrsvyWw/C4kt/d9QtDsQvJCKLmEI
34m0h9WsCJllCiFmmT5YNlo56GQUxVVfDMMzhh5sKOli/uNHqbuqcLXQkdZUVJ6pW4og34YaJ39u
JaS71hUXOBuxMMpL68QExScBiXA+FYWLL6GKi8P9QibevCyrcn+SGBnB5QWtPW6NZUOhKKRRGDoS
NBDIEd8MJ0B48ASEXaE84A8w8xDZuhZuWaxhwE85hNWRt4Sc8a9yI5ZvyeenyRm4EZaavtCWzIq3
7ODul6RkTQ7+LJB+XP7VfRHqGzKQnoR/ULjmUqV/905NnaQaowarTUnOoMP+pjI0PeSWzUPGxdo+
SBwCGDi+jjpqKBQUtzVwc6BYV8mWIv6rXvbCYgz/Wd4UY8dcac0IWursbLwkOs7qHeKBm8tOdxFP
kBaCyr3qCyXgloTANaALa1aQ8QVfulPxtRBk2E9phNFO5nHFORlElNwRVa+DUAOj4pP7M/jomV5x
HNPEJk4ux0kC4gng1VfIJ4eHpljORKyRc7fJPnghDnApHrSbKv6MWjacyl4+G/3nmnykK1z7/B9Y
e+gwMX5f9jvoQC7ltfe1WmMbN8JkweKUlcqXsNnGQAHwRn+MamQclKlTTEyA03/iLu1fZWgxxshF
q8f4HsWFxMP77rsoWp5d8cPQwNJfUCta50Qg+dRKLtsi1ygTTbhOkWuqDbjyV21zFusUfYRUDkGY
Y4hNHPJwgUiQeqZtcRJ6CcydNvJFtaE8bODwbnOuTviUsHBMuM1IwTn2oTDRDKc1opkEHr7h4r/4
PwWpoK/qmvlblnL/1FsnMRjcbH2FEH6U2n3I/5LZx8UdBtL+R/3XuURKtoJc1OWOtQeERwTdBCPB
dTcC4T0dADu4a8sUIJ1THtnYs/np+LQPl307jqzLciqFOBm1MzjdialKiXLUI4ENJPV+qRYt7yoe
Pp4WclAB6f7LKktbljsnEhYdPrklICA/8wpV+9odq+Xza2TxZ4AqrJww9qUq9ags5AJ4WJ2mouc4
iP78zN8XS/E0k23dqqtX6XC9ts2EtczG4/oyf2YIqzVAAJCM1UkNkFHDyCrInKaFqgW0qW30iR9G
XPyIilPsTVVJ2WoHr2sGI7ZhkU61qzwUW68BcCZ8GIWlFSqiousnKnEOIxxHAYwQMQvNvvwRwe7E
5JU+uRUkKaaJ3OPHR0zFOiiZNNeJ7W3aNE/j6mjgbpLiOzsLMuwyHhqxsO13h3UsqXn8W2Xbx0KU
vLMz4HZ04QYAXu77rIJYZVyIqdrDMQL5xDjPGEe1NiQmH8Hq9INhEvGWatNX7nR56LSjN/ZXu8HA
83x7xfr7zh0QNWuJdL+SKMkOsqqaC5RTTJLJ+exDA4Sif/EcC8jjLu8pNL2suWtwzZnVVzxjkqzF
w5iE7XC1W+W6FJ0dAA1+jENch3Zc8/W/EWY12UUw3PdAaxJwAoshXPOdvesO+0fuPAPOQruykrq1
nh6Yn6cdHXrbvCid1hBhSV3j/tippKioj+8G5Bz8SIWfw1nr6n6ybHZRPPvHzrOOAPzzqw5WnJdl
00RepK4xlsbXV2LtXc0mjLwXD9uO3/dkzFmYtXY9f9h0XBdOAc+kD0QNShwrxHolkrjIal/C9etS
SYj5L5rPCXa6/kyYoEbzmGhFNp3kbNlo/AY0XgVbAGplL7WK7vKkwC3cw2tqWOCUdVrOlQArlflW
qavRyB8ge4VW2C/99Dg42RP3g9TXO5xfVPnvQM30+RxKfcgRvsulcT0Sf1LBjJZQSyiraXAW40LJ
DWh/8KdcFpN1ZH/cvpYY/fPjeULdtwnYjxmNySFWRzS+LILAGMuG6t+CFib8wg5wBl+zO/1fVbqy
8QjWJ+DWSKYFHOL2Y0MwIaSE8maDtOFcpLGrkxFV0BfvO4ojmiW9fydV9SeOdfhEzChet9Lm0f63
g7AAG//Io1J6EObcWHxGmH8SpE+uK/LcGH13cpz7RcXe8IOWeUclo69uEMwDATFP02vKe8xVm4LC
XrrZdQ7YyExlIpZ0ATlB0UG07ovMDAwy+dXtB0H4hU/8RqUVeGb/GpMEmTQMCqeEcJFK5w/n9qLQ
UC1ld8bKS9O2vVezFXk5T8u9hhiEVquwyRnAvxZkcPQGp+FnvMVb/PxaGqaVDoSFhohcSzGTKNSQ
+KW1dz8RSb60KjbQMTbXEGulHZsyZcCt4+RH4rYqqHLZDF6v/l6KFO/15tbQElKd97V2+0WHabHp
ZvMz9wRA0I+Mo9krPpCJ+xNOwMdlmztHWaX4ru5reiJizLU4vD8kSJhh1Lo4Y7fD0hndBmVTHiht
Pqqf+pGZnL4twEYro6e+X94hpdqxrXrKbBLyMzbrjvrSwbei25UQtwhPj5OJ8hdLbTegq6ObPTNX
8+o6zQFZaL525yenh++i1/f4lJK2xpVxcHtTcnynv1oWBBmoqiw4Y96zZJlIJ87owwkXbhiKJZ0A
NaL5fsYL92Vi/rKmVU9Xti7xy2FpcKeQAFTMzLzVOSJaFvBtqfAc3lK01jvA/CN7eDMB8Y62qt2G
DJxY8+/094TpXOh6/hcuFmeCH6NcSZnrCCgDCstBMOz+E9fncqKZNvtI2v3MgvzuT76ltMceV0sd
ft64ttb472jl9Qq0Q+hiXWm/rdYh5xASuZZSvFmotPL/O847AOcDHkbqNfN2TQ+Dp/rzKE/8HkdF
gLyRuDRz33nb4Cp91bOeDM8650bqUYZUIKVnZTBzD1HZMig+EnQghvG5qR1iVopMbKQmfkWw/MxA
DVKKPYgbC+0n/B8mn5o2S+MbXXz+Lg9VscCBCKbNgoDVS4PdZj+kkxTHgLOHv8EOO7+Thv0ApxWY
7w2ySQoh5jFKFF+T+TLUdpx29JbsYlna9MBUGhedSHHoY5cebSUvkZVTzXzNNNBkhbz55NzAHF76
hhFxsrq7PNvNUsOQVMXWiUyYMp8Bm5LrJnJ4xtQ6GEqPQLzNCfAzG5criwhbnBGwkmGQPVCEmZc8
G4WULopW+DuMRyF8+xiFtMeTPW7EPhoq7eBnFlycHM3ZwLBiKhQqt4enfd+rSCuGsNRACzRwUxR7
PlIIDbPhDU6B1GyPKy/0Flv3BY9JKrvEMNVzXTQCGUCUHppmNNlAMyfx0yBnlk34hIF46MvBZFtt
Ir4nnUknYIhMS51R0giPuhxmZwH/PtUNpWoW9wbrzZPvbvxKbQtfCaCVXu7aU25KWJEBVUh2p321
c7YyccZf9M0pJWpA/tIPwegYWQOLwNtECX8DzSbowkiqNqrYV8YUd86wKuwtTOT0hgoKIPdKr1Tt
nUB3XdKCSFKuazcP5vZ6w577aGsjybWL43iAHX1tU4BABG/yNs0jNaXz/dCFB9msqg6V367BHJ4r
j4yn/EA5C2SbGwHXYQACWVAs0F8QCZwYiE/dlrB5VHST5DiN/D26PrF89LaHk8nsOhcIAvIuIJ1e
CMeDe8gwXlV3JHDdLfVDaAcMEoVT1WRUO2tX0yiz7psnd4JBnbYZlwbwUoDu5w9M/fhEvf4KecwO
2wI8safjlcA6mEwqIZRi4UhF0uhixaJLkjXJFtMgGhaqsLrPC5jkl2YPZIkY71kOPEJweJc/DpTK
SKFMIj732A3jtpa9efR9UgUztGlE5SfSLO0t2GX4mrvdN432uhqC6mjMuIobXfGbvmV5O0YhzbJg
hMA8pXhjsJpWAkFXOv03X9glV/oUbrNzsmKW3Bq7jkNa4A9/pt1cgdpknqRWjn74VAHAawGuGzdE
romNEZHLFr1SRXGh0UoYdn6wdkdAQyLpPGjDdRS0W7wcfdTFSr1m4EK1UBMv6uEtFmco0glkEcoZ
8vKbki7t3B7/3fJLSoSLll2CF6feKvxNTw5ikF6iGtVygvWIiIJgdUfAPHhQbIH/g6R56bEiLecu
T5yxRyZT77BTcE4keswz3ZvtSI9nuTpWyexdDUsWbQyZIGNetyWCAiwECLI9/BMex4Jr02t0835/
QcSGCJYCsnrOZxgDhtaCrQBDB3a3rTMkzSmdXFLRglwLHmgGw548AfeIxk22NjylwcSjBMgRCEsM
/VZ2D0sc47R3qNX0OnDG/nZtkv0ktMsVPoFjeTtATRTkNul3X7COHiONk1ntOOig5VL2+xcfzDM5
gYKCjH2VwerzQAsJKaOmliCtwogCBtdPEoZ9A+8OWG01l1i+uWJXtl0XBskkxWsyFz0pAREgKq+b
Fy/YlJBs23HVh2Kbg/r/3idcAM94GS8AHNB9Hf6fhAwDiEOaC4s8OG9kmgGYL9/vuPvS1WgTztxt
K3V8KiLzOZykFwvjtIvY5MonNvW2qskh5UD3N5lStJKG273CPTr4i/fvZvlAAdJK+iCErb6pnaBc
qlEZDxGShOfSRAa68pKvEKcTeujdTVQ+mQwiv1/OIPiiGJdYUTwxwL007XtSyKsyw+f4Dww7Wzm9
iJT2hQ6BgBBIhyxMzeQzNWgzVfdhk7fklNxqd+QsC8Ni5hindS/bq5gOY9FG5V8Q7WNhBfgkXDIx
Zgj64GS1GFG5p9zAc1quyelvxTuqMMAnOj30tbI6Gn9tbwGQCFyc3ZCDT+SqIZm3d5qho2So5idk
ZOWcb/ShHIFe+AT+tHBi2M4ZfHP4Z9pHBoiLXZdhht9rXmKA+cOyp/KVSJV4sXe0mCyXv3avGTH7
+A7OLyQsj44j7gsPXEbR3vChlsamewYeFAXv9ckpWUxP9d2nzOK/b5k0IFEyG9qUohLJd3UBNQUa
Nknr2aB3WED5Nmr+1OiI/3Sc+TEqOevjetuO4Cl7J7fzwTY16HYcuU+X5HYxrSnfKuoS80ecWQ/F
S+bj9cUrQIFu6aYvTW76997IePmMAHw+p2YvSkv1ZP0oj3vkV33oCFwewD6Vd4Y7tuoInbA6rLmW
zgeyr8H0w7bLv37apDgxrlpFgb/Swx/Ns4hk1ByP2JJDsxZpC3NRx9RndopTRxbQ3d1enJWFker5
MUDtD/hlszWdm2RfVs7WLkh+1eEhpb71eWHVVYE7JBBsbr7cmQA5n8PLqsP/e55vJoMbTDdpKxTC
iKYt9jLC7vErC58728zY4E5n5MxGrCqRjcSI6eeFW/gZa0RA4stIP3vAfmF6Dz3QZBA7ICNdkBwL
cdh2FTU1zpKQWtfgP+5l3Dl9cxG3efYOFpWmE5kDVAIahgxlN4b+EBR+Bbkm7nOiXa4v0hlSM+uF
a6Nt0T4xGM2WbZvfbKU9xi/BuSK982LuOX/g5U2mOWywEwsVinJauTUE8URz5ZvWjgR0DNT+JuTT
GGac+cpmTPb4ubARmXtmjyy33li8JDaX01IdqPdzcYtzsv3pYdeQcf7r2OZjwpQQxJGvJ0aCqI0j
hokxVoi707ov5k4KBeyu1NflxBzlncsrFLb98pcee7sycdcbO7Ow9nuehoFoKBuE4A0oxq58pDYq
Fx85mttPz8SAB7rCH7/Gg++VxVFzeNlDndfeSePRnNl2fmjwJWFa9nqehiCQYURX6FImKvYfQcRR
18jr9/ifsY0IqpDgwP/umhUzt/E40WPIZR/41t0V73I96RSBI4mVF9aKAva9UFcUMFcEFCLlOpx5
3JD4HZaN8okiZmZPqqksDz+24LeZALeWfeQAi4z/knjbvl+Svb4n4o/9h8wzNis6eqSWGr6XQDVu
bKQ457COlRjAySrR8AtisnoPPtKGr7dfbpNT0Tz28wfsQNc4VuE+MS93STKtnxPSZV1L8OLMrxCI
3Ap/SbLdCZNWFDygJ0eriSJK1gP2BIdmB9mRG+xJEO5bj6nAd9JNpEfaUq+MwKgJggmoAgPqq9OH
myP7s0Wp/kvvXowrXlgJA4zoLWabvyWWKvUuaxVgIt1iOqRO6GjJixD4nXAHb5tdsWsl9++VmDti
A/aKcpR0PWRKkFOzbDpLEx1Mcg9l49ff7S9LvBipOmUwhRESIRS9QPV4+YItAdEgBhjIwg4FafXe
gxustmN9exgIyo19CKZKmuwYNanDBCeD50RuFen52EH1T4xv048V/m4sxStuZKc1NxsFtBGMN7Ln
XWjfowG9ust6IFONik35VlW0op6uxKAbI5hwgayUoxiyn5I6gpZdBtEjG84hetqNVrLhbTkkVb4K
4CcoLvXVKu+OpMLSO9KGzj2V3jq9omK4xfmvyqGEe3XxcdidE9NbhkWarfJJdSoWhJlXHYw3v6Dt
JBpBd399WY0saPjjs4flBf3tGKvQsDEBE7C+OLeu+Prss6411zkbYVC4iRkP0hhLUcdE8lv4NVbZ
KdnflO2pVBqg/malhQvFVWEUA5VPDiLKcVfiHjUxYfpqy0EwjwVJ8IvBCArjbjiQ90hC5Yl89mQi
XWprgLUer7t8kD2v/AHEYMIUhfLzOvVXHxl/DKSMm6BELvJA4yj+bNK4RBoJH/nPy59Yc1fq3IcQ
0Smg5pCv8zDTXJJ+Vn2jMd40c7uFmGoVRjnpgva+3Lxj/3w+C4Z68wx4NKFyTMrpMzsoSdUqsDF/
kcV6PJRDNgEZeG1bkHbGNusvAOIMFmgSR1nHs6slz1/16FXPtgOpq8WYSk63e0E5/+fdsiWlkiFn
2V7Kt2nBWKWvpQRtIZIgK0rLsSbX4YMvZUHcCPTe/v4gP3JcZSRzwWkPzEkWj7mwSrKg3TXhh/JI
xAFS2Dw8687lm4JL0esS1Isg1LAHh5EDmXCQA03TN06061oelFtXYSc95rj+FgeTOAcw+Ss+LtuK
aUKaDdFAMx1FKOJMEP6eYu3g5SpjtF6vNv2RmB2ApOlOJhsovgGisx6Hd9EliFpOygVGRxdfKt71
de+SX9NQxHIfhLi/M5x8Zn5coTtznyjMwJfrhUBRud1NKG7oi2IMNmtin67yj7qpimc/gYtXZ8ya
NLjUGl2ofIfIjrEHNAtDMrpuLCFqDVbPA0uAgxyJ3+aOxJzOw8IaN07Dcre/IVepTE3vMXUajBma
N72j8ecUwKtzQTE9OpqxEHSQ83jL5gBXofa96W7dJSaZfrCTMnEjtUr4z+RqaBE14B6LOJ505X6I
ozrNYXvDexH5QAa5IozuHqFL8NEQUAQvUuyp8+Vwtvo8yZ7Adfc2qbVD0Azz1Fo2xOmaRFTmucdC
WXpWysl20cIe1ZbIBQc/+tNzmmSW/VJjClulYwlGgymFjviwe6rKCK1sqGUsnvEkgo/USFQByVS5
Bdo2pULiwTkzY/bu5JQgcD1+W/NBBqqeGqBCp7lzI8gr1mIwJOqCTG26IIfXl0UhYeEjtTxbnpI+
fbdFa5urBrXSR5epGlRDIb97s65NQO8HsN0Uc/wbwxAMo47cXW+3KfqorKXnbCku3Li2lavN4F6t
VgS1IHbnwl4T/rIACsdZc5pTicJ2Iij5U1j1xKjjdmzGeD0JY4l09i3deO77bjKMPBODgXXf4bU+
70swZAfbdmW63CdCwmfUgV1VRVXdyQMSMj4PlftSrdKsSHVbsWIss9X2iTEBusFuGj4Zgu48RCIg
qhgDyi2UePQ+veoDErnKhJMrmAltqLSZMUaz3r3sbt8a0Bbs5UVJUazNghA1a1r1wMiGeiFFM3+H
8S7oZj03ScyX7P2XfEVL+0F/4ex6xz+ftZpyjC81NH8mj53HozSbBmYBUV3qBy0BxA6CNblPTzux
vJC23KRtUe5sSMq4OyGl72aGz1sk5OqGVw/YsXzLDzeg9WIPfBxxSZbmxJRNHjKH4ntUzcjR9tK/
xr5qbG5egkE7mMhB+v3gUFNeWI5xOYm67YC5ceoXUQz7v/nTgLdIMZonBQLmgDYihSIPlZ9KS/Qw
iW6a6fmQWt0U6AptjnKnIMo0vTIFNO/2cZVGPRGAny6pm6P+7qPNGNTd01e4MFON3WRuUnwDsSRE
SUy+bvQlytakLasyJ1hOESTYzJPikFuo5Vb4ay0Zf47TR5vVxTvfdwVGpD8tp4eA3TMm3YSLoI0W
FghbQTojWq256fPTt7nTnWG/ZAbOYuGMgEsEaYeHJvFce9q6gucLIKiNjree2tVYdHFMWHc6/pOn
JmoPPY5Hd36TCCJkvwR77ILUggucKBNIKaxoAwQaKjh/Rl+pOtoDbvWmqhjSxTKgioF6SLPl2Pks
oherqaWNm5G47z8aaSFmGWQzWRl+wiJAjFgE17KqAtTbIih/7JxtCVRaZNvJXqzWU0jBi8RuGrZt
I0z9qoSg6U9AoDtusq5qxATtdG2IwFYIjIc/0+CPR5sygJpxXKIFlE+1rxulx+wHKQac/rVHl8n/
6c3xhYE7m200AzGyk4cFEljqgAu+3/AknExskKAHi13J/1pb2YbrNRB71UFlHfKBvdJlHPCYFj1W
iDYhB79UoRJL1tvs5eHM5hmN+LCBy75MxiCOYzbrcDGWczkIAiqRQK/SzV/IKIvy32HfOtB38Zxg
GpSqm3eJLnXyCUOzIVvy04Pm45BKH0WQOB6u8wXdPGdQ7zb6LEX/ZJiSSQTudKie3iabQ9ij2qsu
fnBzoML4DIiYJImIRF7qx0lHRnPQCBkcXIw48cZIKXnFabSpFmj9kTKoNuc5OluLU2ZhzfCRCUBg
rD4NXoe+VgQTQEGxWChyc1QdJhz2w/fA4jX0cdGte6sFT8IFMQ02h1GGLfpPShjp/JoJjsG3Ne5w
4gwPIDxRLNv/Zt7k8155pCo7CG98l16WOFITAEcSzRg4QhCFydBgIfbNt7O735020Q4u9vBDju/E
z8w/F8DlcSE/yQVGVeXo37plkvwhkdH0gAau65qcT5B59USzZfyeMv9nHRqfGtmPshylwLYclxzD
h1CeZJ9/KDWBNyn9V4VQ0AB4uVrTU7f7T1YDUVulZVv53+137T35SkEAHnkI8iwBWFQxKOq5Y37s
eVGSuh1KU/q/OdnJzxFg2i+DOvIWK6Hj3ZQz8r5M/AUbSktdbXP9dDXYINwMK7EdxzTll5WXsVIX
TdvwUkurTGMGuVUUovNPvOzLR9e3EFYQqil4U1kv8QsV1Tr6ZhCAL4dLlin/eKUp6rKq6l2K7lsA
+XbM2rri2auIZt7H1UFNSuWigTpuqq0qkx9kmNHN0MIq5DO3bxa0xI4NIYAO5gZ+7imlBogpVGOQ
cL+12IP1Lg+XuDHCGxLGILnzsoHp4Y6UftdZ9YZJVonGpMINZCczF8jigKpT81JXhj2CHI/KEdXj
iBzGscTw9JRYoKF10sSP6oIEA9TF7YOh/q8WfA5qgEX06xL3RTaYjueChDmDx6KdkECbfBO5DzxB
Cyb3Bzjr9bXHsw4yhm5mTUZhkoYBURT/gLpnBYRKiU/If9Ik++XZ4vpmZKI2EW8YMksYP85P3S31
UXiduOCw5+v64t/5hpYRhp8B0s9biwhMZ3Ahq6p85AU2VrPe80bAMVTYLoO+9hOdQgJT5kPBWP6I
6q1lt1m/DNbj4Saf0C7MdIh4mOMunj3/XAVhBzQZZDViNxn3tm59xAukvZ/OU/B4eGkvIfIHFVAe
N8ySoYXwN7ldPG6cb/lWoJ3TEwczm33+aziuNVZgVUvPTg7G0eFJn5i+u9m0mDwpd6fWcefWWd8N
y94sdh4YdyBGjCaKPCMmeHLLCrC8rEoN+Bmc0l6aMvzyLLVjlMCLBQzFM86GCH5omamP0N2C/qcX
uLNwJwPPt8YyQzQ+npELuAjTsvELYwUgnDRVQdkjqIkdar1XO8XNf40YYfcHZJYxahmeGcFEFtIm
LJxAsO7q2XSbayFHaaq8ek+OkW+yVA0GjweH7AiaLn1WEILiHd8QDmtg7woSz4AgL3jFtvv7ReFY
f2Ti5oWEqwCgii0dyexIQtgCzrjSqEj0VvUuF3bu7UT0aj/QNNK/XHzMxCXpyrGan59Ygyo/muLy
LHp8Ogeke/+LRdxR4oqGbtnvg2VCDvvB3ae3lDdokkcC3ci9+ZR9gwLHHz0UeIaJ1YMC7RgE6oeS
i3yHO1COsTDV6OmSfmf1ih+udFDu4eQIU1yUFpDZ3UYGE7OcnFfapvkGEJ92iSwgY/O6enwhmdmy
pNMVEDbsJZNeBehMNCTdd+wa3/6n8H6tJwbe6MTA8lOVcyugyEkjsCStEuKikIK2AYsMy2bVx0jo
yL0JarLbQKwjaX9hzb+7WO26kZ6ZJkkPAhHJQT9+fZecjEW4YAn5S1fDoQ1Ah1Ru3oM6X/IlALlP
yhafDbobYzcreEFrmwvN0NFFODULIqIzZza4tcDSTbtarRDEEz4oVXUJwK/Px3/2H7VjceMp70O1
llrJsS3Ij7dVHc6F+vdMbAqfsN4oLmzJ7Zz8LIPt6bwHoB5z5mIJWRIKI7noxFxDNUvNWXkXjmMJ
E2NsZeqXtJIUi0jytPKQ3cgjxES99nue/dnFFVn0oGejeLzLqxdmnQz0CBwdy6+N/l0lG0xjKGYn
eXF3CsnlMomn8Hf4SbeLvRQ9I+j+lNwsf2Mmgs/iaWPKC8AlsR4icH3LEYZNc/1U9TGG4QjXKpr9
OkokSIv6dDYdmhszjEtTrlz0gMvrIeplYmcWxD6uR5BYbbtXNOdgDGE4vzb/EWDOquKtzhuTpJk9
euPSYG/ys5Sg4PJlOPSm/fZc+qvzQV6BznBpKWuaNH0koAazclSZs9ApoMDKRm0OJj4o6PkG2CWe
Q/amycU98tAovYNk/nj6QJum5DKc4b27aymgZDYT8Ttv1AjFZFGadEGBUFwZp414vkhfwnYEyGKk
Y6gaYPUb7JWhGtI45Xtd2I9F9na4lkdTv7UUTW7rslS/xdB1tueI1qxB9gFlI8Z4fpjB5CZtNXSH
/WZdfkKzuRgf3GwZFedik/KDXLfxhP3PKkTlaSPtGbRdlRVRLoO5paVXq5noYVXSaPwlWM9X/O3I
GqS9neDW9OLwQxjDpfXhFdZ4ruNEYquwV+o/XnRzfKn4i+uwd7/evmmVgUQx79Nbp53odPU6VvqB
B4MIkd0AP9YEo8++chdOdeuQwgtuShyr3GoamBsA+9i3ssmhocNYgV+JKICcSlKEjPlhuxaG/wlA
09jccs8u4dnsFfpXrL1q9Z1MV8TziFw9/cwHn/Y1QD200FfR5Z0PX8imZUdpiUpjJMrzesN9QjYt
N63UBKyAidIeN/eaPS9PV6mnsaHgIj/Xd62ukr4V83Atg1KKWDsAHMKSL9m1fmFWFP84u2IAhG+y
/S7IGBxD3daT8KQqrpZwPC8pBinFn0LVyy6OwuiuddSkOjlYpl2yNiic+V0Lze5iUyB/6xEO9K1f
I18sUsXcMoP/vGe5VHcuhsJxzLnGjcZD1Ztv8GyjR0MgCrFnLK0od6gKGXtVE54VGnT9aJ5tbblD
tYxJ1ALb96oiSlQFJarLu2wvq/n72y5JZHO/wzakoj2fx3RGAbqEphhyrIyTollj+/Rn1oUoT22u
HAuhpy+ZvZ0pf8FCrg0EvoSI9ERru/eVY/8ZlvMek2JX72pAh3ivl/7PWU3a2F4y10QlS9mB//wz
li/ABcRb464rsb/70mJEzkaITeQnyAZGP3O8xSQ4E9UTDQxX6Gd2EI9EeI/HuBstXi4pmMBgcUqu
IRG0nOc5m/zASWSps6mF/u472hupvh1+sx5b1LtcZBWIBd03/ffejoKymVsWhrRRrGSseqKzudl8
8rfKdCC6zkPaaSzEt16yiaO9E8H+qT+YUU1rV1vYwC80MmI2hr9EyIy0wDm0YPt/uIRk8npDndEE
r9SgrmBQotReqym+1sIW42Za+YZaS2yrmilt3W7IjtDZV9CFySOaFYQP5pZ/2AsqluqxS3VX1BoB
y94RLtrGCuZIIIfGxj9JTVS38ihbp44IjYc6vVNB2cdVhKD3obgw3+fKrL3+pvR3FOIuA35CDZbf
b81NQKB8yWlnXCUOH6PJNOvQg6hZltxxM4qbqzuySt9qjP14xVu4ysanp9kWmWOUGqN75Mez+hZd
gBrDuAnDrAy81kU6XX7uZfQLUFCmKYDJ8itueQXqRXKGss76LwqNwD+Ksa01ZLq4v1/ofDwYCfGx
5Lf2dwzb538L9KRxcyhGm+O+dIE0hndQ/lPD+WX8ORIJylZ9gqpgbF5TfWqZkIKQeK1zw+leEXuH
kBXkQdScrmX0qLXRkSvif/ThnDoG3FwKXRcG6ULyvJ8mR7+oM8rqwQNDNkVEFBCogXlODimrMM0L
yqVbz/FXwQGTyZoQCnXWGdHH02WGzlu6280OobB34gms65Y66iEin9D4MnXLPSOy/wLr32X7xlCd
GfxMCecXOQrOXxWOKvFwx4ZQwI30tYvm/jlNp8hsyZtXxkFEOkTY26OzVQMvrOhtyt/sEf7jlsWS
5dsFn5pGYy73eUdaytgSMwHVeW7GaM8vcb5CdoajpsHGJBthykwFMHB09T1YJ+HE3J5OG1r9NbY2
8BQL66dBfMKEM0UJ2bhIFrbhz9uQ3ruPe6GzDkK5m7mYa6JBDvENMzo8qsD1VNyPyZEWDeQOwNEF
bre86tCwQa13rKvRoBjp5pFMRz+Ex+OADLF/qAOHC8YluypFRhBPO5siXn0Jb2htPjXSAju+bi6L
Zx5Lid5Ls69CbYl2OBoFXaSh+bYJ7bYXkB83qPFo9WP/Lgjxbzg7ZpUqEK7AwouskiYbmUJheDNi
3Wn/Ny/ki5QzNIXrJXioR99uNKfV3i6fN1UZ1pk+lTxXDQkZXeFvx4kMun4LuL7Z1j3xeiQGRfYw
uxPKbR8OnAa3ty0143rzDGTPUhws2DArrG4GKSNH0R1X/o1ANJnsgT+2OAnPkN46Fy/MKeub78+i
v1bOhFC9zDe3yCdgXDfX3f5HsAy/YfvNGTMEN4+zSrtyZ8ix0ISFdC9RIMCC3NCiNT8OgmPtvWse
aMI1eWuglba36cDFDWDIbmWSy7yMWum4M4RxN7X6CynR86RjpxEj9RwBg5L80r8h8BUvh5ajuVad
YKeEUMbRqDe0Pniu4b9WY328qDUeVc/ilf2YVhg9zw9ogy6Ux34R5heuUX/j+toqJ3aJwBYsHmnb
WF6W5/zul6pfJf8d8G+QDknqZovEVpfXnbOS+MbWQJaNBviWJc4hx1N3ohlldyizkF/GNYe8U6ij
uLL13ZLfR2R6VcaFeG7PoFZL5y6QeTvW21ineBKD2kK7AGlo53CaFYp4Di3fOochxrjCLg68zTMD
7UCrvkxC8xDOMPqQIzTQAx4+HcaX/szm4nEBSvGVOP0vqQaF4DiNAPx5TP/ZG/v0WLJZaUEZ+1sB
ugEI+5fGmUD1mg931/GQo/p78YdOfTzIAyC4gYmOaviTLxYOV+WXrp4UITpwpTC+De3Ip3cUiE7B
3XymZOauzvHJC2Akrr342jROAC/dFxuL2Y0bLik0p7lSofv3njho9rM/dxumnCpFT6cUWY6o7dcb
7fu2SAA4KdBNhQl1Oel9gXYcaIvpVGvPTGoh/Ux89jm3gK6I4KsRDXGPyVf9y7Xc+gq3gYz3I13B
aIDFbS2ZueJJDlMrEg8tBSEc6M7H0nBE8gjnkJFOBq+U4+CQeGqgI7cdFWcQixTmsevaajcIStKE
h0G9Hf7DVMMMfP1wJa5hRM9X6O/vot79Fwu3kKgacjODUe/YrzdF50GMTcmnsPYYJVxCELnxxhlg
1RjbC/4Wh4M2RnpGAYDIy/bLeva8I/DLiwnEQm/T0y8MiKhlMDgbT/+0aQonX1fwWuCg8Ih6nWZS
4D+P8R+qWWkhrmph3KL2B/c5czYNYsx207CH/uqG+6Wnvx1/3XNa3zZ+xBClekNZzvQARwgFLoBr
2CFM+2VHLR7QSuimvqrHRr4G3cpsC50OK37iRJfwJB1aOLdpQO4zuhXPb6d3k/71ryg4lkhK+nCa
8zUFi32dRGL43OqXA+PJy3NkWPxbLmj30jKeFGe0iJffTCjjZhKopC152D7TvwJ7BpleMi/DxAMy
KLaFhXjpjFQyEuG312DoGaeUUQ03U4LzLR8S4VZAP4VcQcvVMh6tAHmxpmtgkvdaVb1JYsGouYun
oISl0nsI+utwonSJVcgZrljcpg6xjyh359gq8bMiC+zWin22oHoRqPFV29lUoWRkJohWBzzjwFnC
1vuJH7ifEzAEaLCFF6lTWzZy6zpUMS/uxHLK/Zf5ZhXvbGtUh82K20lIuDqZoQnQ9LlkABoW0vpf
5TyBXLSNdONXsfgCPI5d4q9X1NMxE+88/MsSd6FKQMBqa8fbTeuVpYHg1+xG/5pT7yDkUtqPbcPq
J4oiq+qOE93cUa+rOd++zdXXkGws/BhbCLV8HSPRRmcGjGxhbR3cqyCyR0EEkHKZRqGzRPNcqJsm
Tcak50U2COtYsFLaOBkuF1lMs3XMMXzyNfJxw486vQbIAY8KuUzoHLSuYxp5Jvn5DDMpkHAukuQ8
037i4t2UO+QGPhZ9mdLZxmqeCGP1664K4kvk5XqbVWoVq0CbhBZzcKl+PJBASorDtWAxvLU8NNWw
/l1tcUM5G+8AXcO3e6DKlqa7YzRcySB4NsYOof/paJIk2fIgwGVZQcTZQ5DAWMZHxMVIjJmVxShc
Yc/7DX+zhDTOKIgBSsS4k1gWnG/sm80A6goPPW4N+wN/wdgsGs8dzzyyGGYp4pbyuz8qShhlbEQA
pDeNvyCXDlktJFaBRiXWrJrV7mNTcy7eniVrDGJrDpRwwPwsrwYyBMJ6CIIF0dLWqa1oKpQZ8ZCo
AaQNSs+eila5FvI9yL4HxsIBW7WVnXNXT5HUvgiCVprUTB86654hEKFY0/9bnmLF9KNKyek72zLF
p/a4+nXZeqo2NlmxKRfFLV34qNDzrpzRo8fZ9b8e2AbS9CdbYbKPMJCFCXJUZuz4AWReIEgfbXBD
6j22we9k4Bzj6lRsVJwgAVHhfgUrp5Rr0sG0N3mOQYZAiPPXijhC+q3H9fBlEUDyfOHkYJjmmO0D
93C1BMcqackn3HMdSoe49Ev4viJWAQ9HcnFDBUZ6BPMskAqq/wm9/wee2k7v3qo04Scdm1KN3Zwx
qj7r7KHevIX1lkjNwvZbTnkgmXeHIxO/zs8xZC0BCt7yuZ+QAmhB+wBCPf7sTvv/TCXaJ2j94lWC
xxkECKqUlT3w5QoSjNkHNCWllMspwJCxx46KlIAMVRHwfWlbHi3bhSG7tt6akMC/L+oaK8kFgBiy
RHp0oo7tcdf1jtTuxL7pjzS1Tw1uOVT1KgT5f7wvM4TgUG/NQU1E9RzaSQF4+e0Imd2cloyiHraF
EMM0SkcBL8MX/N04kKuRgaqwBMMyXuAgMgIBwChbhuZmBLrGPySB8Q/+Xh6seLqBdOiW/jHpYC8a
uLT2Gx/hMuf5GGW6tIMPsJxFWOGN3SHgNYUpyBEtp3stqSjecFp166+TZ0ASDgAQIeeyc8U88nkF
NhhzOA9G9WHCIHAuqZCAdm1YnQ2SknRMFt76ryk2PSj+Y/rj8UxhnL6Tp6p0Q+89yJOE/BrRY3Zo
DmOdWR69WEQCpFn5VT/hKTMYN7cB7m5kxIu7TA5FPwVZizfqsnaUWubtizd3PKoNnw7i1iX58RPQ
aUHMDRX9VhtdvP5GNJjybWdEjf5HSPjnF6pm9a0dfC5jpEU2oYZNgJw5HQceZuaxVGXTQkK/ZepP
1/++NOLjaipJTKGgTZn+nlrcroSX6/rFa/upsLjd8xbBdTVaSaS4oKYglcdIjFYUZnMaN1ulHwkl
d2N44e884u8sSixLtibrV8JAg9pGIek/xOe8wAyyLb2tMeielbLwXWiHy18z7AjMMqyg6LstS4y4
kjJao0ikcoVHV8oAp1OM2TIyNmvi1ZKxqH6AcxEzp+KCzoeScQckm7cUSgSEP7SAEApZnIGGmhHh
u3691UNeLQoAD0krz4KREb51lTiqsDbUx8Ery/9GA/PJ7d75I0q3b//DoJcQ+iBesnv7FJkRJRoY
gWay/vrSnXR6hMAqJ72ro9bpJtOVKkmbF5FEErszSqd+m3dekowjgctbkQotIgYVG8vRYMA4ohwo
RWD3XFThGBkWQbSztumvnU2K3L0JQApI6LBn+RKVyHICyqSEWQmFlHCvP+jXxqGKAmU4Ys7dSqRQ
Ru0ekPluJUgt0W8cRQJbyhx0LH3Jqi7gpRLE8RQbzHkyk32mVlTHh+TbjpJFRwiWx2+h5WMdhRIo
r95J16o8cZBvX9761AqDKwWL+pjv5567R4chnHmuOXCgPvE97mU/WsgMaMcBSHmvU4vRH7ZqBVyx
BKvz3HgOCxVUnFa+YCiKl3TXYW1ICIQMMatkGR7e27lcjvZ6F+fJ+gxdnIQQdrypxSfZ4HKHfCBb
xyaisbo/cx2vM37I0I2Opl0S9GAR1lEm+kU+p+RRrQ87BHieI8Nq/uWzVHloSnL2zRNNeEsHUkBX
gEy+dmIKsFtKKTG36k2WwuzO/4haA9ZsvN719M1iAjSiBZDvK2r3dmESBZ4y/vfOxVdl538Fkhra
+5CADpTcPcQZ6jRnkWO62oucx0VTyu01PNdUIkVMMBLH2Fm1pdVs4TnVARCgoLO3KiJs2VDppxp9
m/AHMsM2E9Bo27a+bBnvS8jqYT0jvF3SLNf6qSoSZN4+fwi9nVssUblq0wH2wf/z/ovKRqYhPW1e
SiGdO1WVW6+rszPfZe9lmBNF8L0DKBzxMaw/j92Md3DBvn7/W3Dz1jY3DphmAIsWeNO05194f4oe
vU8GPVMRJO+9s8DEAmSRQev8Bf7ewkvB6R0wtdjtipJcqzy3l5jSokr9Ng6LjjTsplV9miloxPOj
qjPTtakVd4TpkvCUEfXRhEPcaoPspXyGOupW52jtbutvNCsglnu6twtmCZcy+VDwsWHPXJ69ciVi
GqSqU+/qgpYMA0Opf5gGp6BfwSBve72gJFckwE8Dw6nxLL1/GGr8dvPHwVbudNsp/Kjo7AM+AevY
u+i+apDpxS3Rg+02YpOecKNAKmFS3p5pJ1paLTTCyQ20FcDaDU1dCM/+9n5lZFwtIWrYBiU+VhXi
0fRdImOnU7Ap8Fvt2Q2NiiwnHmi5ViknfPVjXh2u5DPu0FL8uHxxB5tjq3wnFYQ64xS+qIlM/nQq
HySI7mwRjxPsgm1DNZ+CTDx8vAkjcg3Vx3vGOCbGz+2ad3IHdBYjEBP1imPpRqVXU5VJ7dDKGIan
hW+T0gTNd5IrAkffLbGccBKbKdNDeQEN5VHa6WOBGdJW1dGZLO2qfHUFB3jkOD5urgHgCU5LImpS
zgfkR1p2Gs0cyFXu2okqtDd4yY/Ts7mUsMZ5IKA/PFNKaKFZk6H/BJp1XZbi7Mdv4hC7bvD31pHN
wMrFD+R2KVLMeJOp0RKeKYdn1bWuqAchRaHWnTzei6R2K4lOi1iPEzhOS97v+DJKBU4XClTRY+rv
sDlLZQuHKl05su/Jp+wppsqjkCto92SuVDp5axlrLgNw7nRM0k9MTgMfb4UTMZpkJ5sephzKFpIW
mtwf3av8BkGDmKHcqotLBJe8wofMQVN9sbjJp8MofCBAu6bJ4EG3Zp3fwWVmPCtX0LCvweuT6+pU
IZnG/6FUZZN7dKPc/FgQjy7z3sdk9SWkcBdkSDPxjzuJigdNd5ojR1nXUouTdGi4i6IMXXE+FQ/a
ZM3m1NsQez6/65Ynd2Lu/QMi89DQYw/Zk3OzslskG4ZWG9z8xUvX2CPX6TRYrISEjyqkKgxUR8jd
tCZAGb335H/hS5ks4aFPtLBshGnRPiPczT6fWMc0hGnfdXnWIjljyM8Zu4GkEdy92il2hhV7CPna
/tfGefci7D5X/IyHCvcILeX1Pa1yAuZHi4cxAACxm7WHS4rNuwRQhwfhY7lNKnO8gFOnDJmzzAfu
Bui1u1F1qEEiWXQLPOjwGsUP5Dx8DyAivksYYVBSCNfiBSmk5gq+riFtR5KHU/idCfARmWFsVPg8
i9zKqtlpFwVU6HxQmr6Bv3SfhTqovlZWl3K7AiKg2MTMml4HHWHYPUTFotI0GWQ2wgmKxf1vyJfZ
Z5L4yTeC1WRmrwKpL6+bVLokQzNbhbtlEaDh1UMibcv/dQTBqPBwbjiI0RPWcFUsdlRtw6ggUv+u
HU0DrZ+/5bL6nMptUSWBsE8X/Y5fINvacfmvL6nxB2wG3M7rVgtlhgQUl/Uo8tEPMyimIXrFtYDy
sU1UbXijZSGvZR/d4V/QsL5j5Nk7AB4wm/qjaQlhYJJAkPkEnm4/hLiHGkWnEiU3SiR9Ci+x68uF
A7Y9exjgqOfm5rAyPmr0/r0CRio6y2n0GOLr+CuO/6A0CzJzu0/iQvTOh7Nn6WZ8egxkFp5pmRgx
xzC/giGv1PBQ4fzpgvJ6JGZmq/ik5YjzyOGQDwEwJpF8BLcBoZE2acN5/Z7z2mWeqWBaNVbGB4Zj
7AtAKp4SNFOBhIvY02bpATcMkG+qHewUOZ2B9AX46qlsDNU4EoffVBTjfzmTaIu3IWSWWbejx0qx
Lka0HnFk9Z+8Yal+S5ogrBlI5vq1EhGDDEkJKbDr/JMqIZVn3AUiTyfwa6uV9VYHn7Ai9AcaLalA
4i562Up/3KvjRIIDVbCM8H3w2SnT2o3GmkbBXmSuOnl3cThUUnHNJTZL6LgVvLu3jJqM1kBu+M0l
L/JXd7zJz9KGELstv3/pvw2l9YJkJ/kPjUK3ZqjY73jidGHPsgr61KZ8VU7rSzIj1iv6OQfisnIO
CpPN3mymtSq3jZUaiRFulpTaIkv1Ormsahg9A5qjmo4UaYztdATk6VHbyjzX9xen5YEthcW3U3zO
7jx6ErZWN+sALn5dIXkUhGfOx1nwkt/rwM1C7DTN2cWMbyOmim5Ahc2P7WSpNjB6tBf5gxDlPDpc
AblovDohX14uRtaIGRmoa0+mO5dgHOGiqYa2SF1akmKFUmejF1Jlljsbl3Zezdxr89tSRu1/VYzx
086O5Va+MqJCAV7fOWcMDgX0Tjrdhs5v4ErfFyX5rGnp//B24PbCKyNuIxreC8JksNVMOSiRQf+m
39J3tJVjO0ltect4Sd6V1wW3ya5eXrPIORPNvxQF1i9XlZGHLiPLAbVC/ZvOlKoD8Q1QUkPb0iyk
26c9o5bgz6XAIFQZtrl9KvE+bXGIbKmKCrOylHpB5K6U7WS49cAZK5CIGsEre4TAGe8Mhq4O7J5o
qHjMiIT4Zzxqdb2GcoukftOEbmdwR59ks+WYp5Pp3iXSDup2TDuwGP3fIG0yjyvifREkn0VYl2cM
B5Yw8BkLKAWdmsbpLENuiVEQmlDSPl4jEk6r8D+d72Sle+MtEMgJVxeF5NETw9p9jYrgLUhB5Y4L
MC3yf/i3QhJgs68ztSU5RFwnIcuwAErTq0m4sJf/grFEM+LakEJ/D0U78a8a+3PEW1z0rEcH5YCH
HmEPWu6hLQG7VvFRPsBRthJVPIx0DJwGyKndiSF+XmkQxxytG/d51wxkWYYWwptr7LTPkQGpTkOa
XW7gmgO3NU0V+xYOZSIeByPFtWFOZ9LBS93fZ9PRJIm8/PkDyBqpBaQsV1yiIbLD/Csv3XGwcTRP
FnOJmQity7G5MJSAWccSjGsOjv0D2qPWdqfxEaHbUJ1gOEhtSd/Nk/VUQL2o4s51ZEHvXBjanseR
11wQR0YSBcp4CzYheernX5fg1Nl9YgzkpZUtN2SxQaMN2+LJOgAqHekGLSnLZFADRNvfY05exVfL
5ubxqQWAUwfJh5oLdmsj7Od7lFuVU+QN4h87DvbVGEUCH0rHP/6uO/Stxx87556xV7ec2IhXEMfc
P+fCkSXzmP1WatbZAEOFNinbSy/ub/tx8tZv4dQW6zuVF5lc7QPi9NqmJ41K+nT6rjaHIzQWgOSF
vAR6gRNBkvvy25IYVw9LUA6dhFNIk7JWk5xRsrZj30hxlMvdh2RjiesqtExgW3h0imz5K2HUN+HN
xNjuYG34KH/8EuFdnOtfq1tzoDLBsvzw2/Uj79DwwZqztDq3UrNIO0k+MGf3lwkv3HTJ6Oq/0j0k
o/pqoGcMlgOydwzCsHfa8Nx9VDjGgH9qCZKp5iWE8rWQLBC52xXw9dr0rqDzuPpush3L4RQNH05L
hgiTKQaPt0sB6+HkvupoYdUymBLaz3tgjPIxw2v1xiPk1sNvxC4qSfkdDUHs+cwwZViSK1k6Tj0g
fYQZUQ7Bm/a1/Dnxkw5raAt1DZb6XEH68AneFTRGHz/ulGLJ5VPtOcuRp6Er7dT6tG5DnWYzp+Oi
0hDMeRQm6YIFv/D5cBc3Gs8s7NU4Q6O2DkyDUSuLY962qtOYzg1fwQQSizHZUGlosxVU4DDB8q4l
hR9/Glko+WVbAUtWfUG4FaAwYaV8iaSyMhe6VeXQk3SVAHiOdoB/+FuZC4p0e7sD0HFau6wKheyi
qaxylBJu/ZXHa6Y2Q3UncSYOpqKIDSVOW7i3WFUYMOK4gnq3s5+K7kUUV8unf1CnlYRm6oCdRLTZ
/xiFMuKPECyozpFYix8M5SIqJ7zVhT0SI0XDTTIrwLb3KYHhG0/rNqKlWuDMFkE+X6IiZsCEPe87
hyPyTYjqkJvDXBh8QUCGWGroh4mHjoNOFV+VhQHD6W46eI6apdbyY66BecbZQbCLUU4akmhkkNXD
KXNfx05UzHMZupF+xVlJJD1Ojcf4yYWewMW5VgzmRTR19KOQbetgh1FNklCfzJeyIBD+P4hdyaOo
1xF2GbTP1AfWKjRSWoD+ky14/dt6jXZqcN+juVPgcdSmvX+dLnNqvyYWEDcuFpPCdU+i27CPXZQ/
bRmeokwb4d6chZFMb0VydhKaYcK0eEutFhoGQfEMjUnl3CMtanC3h05R9nGRDAcopKg6vsw6DMB5
GX098/u9DI2ip4uRqcQiESGglm3XaxlC12GwcdU/+4XF6HiyLpMqmA5Mf509ytRktdzxHv8EekrO
Bm0DmQ36xaARP+hslil9/7/r7R1ceHQn+TNyVOcEf9tlN+jY5CuUTlc+Ovec9e7X3NOjAZmBek4j
vbdi3mfaBxir0cEClTIyUnjrk5I6U6wEoJr/PIIIIPKDY2OSy0Mw5zCpyc7m7TXeo9BKuXBQ/Jfo
yE3uAv4y7R+QP421UqLemb59oFgVVSamCGqGu4U3MQvBwDcwjNkYb73QlBu5aD8ut1IjUv549kaR
zlsNiSnuSDV9BvljyxzV013Vb1LulSpxJjG3YiV7zHuPQZigu41RyaAQL9QhrCUnN6FbQELOMJtk
yM61SLGZNLBHU6h5/KvLYlCY1NSuX/DHggy004906squkG6pcBAuRqzUTzMJciEs8uqL4rJw3FhG
MXx4rRmKQrs8YkeY8fNMEfoj4lhC1l2fYhm69iR9BxMueqcoFXJ2v7OL0cz1p874bi46qtTQgf9v
WMBeFJLYLgn3HPv1zcFG3DIvou+vonGn1cbQQkyHQQ+FlLuGoork7a3nIFo5XHLnQE5o/sekqZ2W
a5RL7bHshehNJhFFfGMsPGmGXOvoaoD/1XW5JHjoRU1Ts/EcnDT91DpIazcwsjzdfJ1hBURpQEx/
di4/IRJjs49xka2n0iJ6oftcIcdTOzNmnbqSuxr904AKnJ5wLQrqch0BUeq+MvoPemJ3Io5/BMCn
OC2CUIVcCj0JJ524x+1OcCdCJ5EImjNOJkdulw1lQEpj8YbpL5FfMjiLNrye/rflGAp2Ecs9WHBB
pJ199rT2UGSz/yPY/YwLyiph39rcPtRt3xWeLS+pYTG/Klho1vUxd63ngxtva3JSM+D70A1f4BkC
X4xGsrZDE9VV0cmARtqWk4n1ODnq6fvF9EjEl8zRzLAiv65D3RErgtIfYYFa+hrX2iwYHjHNOKkX
yn65xad47jaKzYYtzFp7MO/HthW+3GJGG/8/eWQ33l00L0DrcNSJguGMeLopBbYh0xnZxNqkhweD
Kh38SDpgxAEfOZsN1IOdUDZxHi7fB+vDRdztMqqedc1LbtJMSR5DLZ+93goHzWtHiz1j0D8ptWRN
np57xhBn5KjVe/Ex0Fa4tVHNwUinr74lLbMYj0aPVM5BhqAJO93TDWq1WQVf5PVIhLq6Jqn8KU1Q
xdODbaKjHcVEfDvtQgRbwKnLS/dQ1bh17ESdZQ4AHRkJTnWsjYxjWXybNM+/54jjvMW1ygSScovk
yZjf7cXdNUTz5ctJ9zGd4Bon1yzooAxiCtaNYsrn4Tcdfm9hmGDN1PJ3llnvqjkDrnAhjWrMEGEy
SVLOgjBVS6qONe6nxzJADaFYQDFoqa6k9PooYf3TybY95fESfwS9m5LrjSr/N1TfbIkS6/6OW5zn
L0tCdyC0JoK+GlioPVu8eWi3wZb56cVJhT1LN12Szv3YRSOy8tEz9ZRYIxtqvqE40keVosWcoOJ5
YFcZP3jEq4XWDgEA0csgvnlexPyzj9ilUKlK3uVOqxQrfthT3FKephq9MpJSSz/QewAK1JksBDKy
HKJ2PXnZ5VmhNFs4Bn253H0Luq4b0wSsWDqG2bUGYIE8qyvD8qk6E3qCFTxmQqSR/2fIaGkRrS+s
RByR1+3dw2wkUwIm5ktuWCOC8AtCeNuIDJTMqPOealiQMwEg3LlZe93E1Ku2BGpyIWmAut/3fn8a
qWfuEiOfkzJtbhZghDzjEa9PY8KhUtBzW777EpbrNEsCVLNP0lDLzJUDYdinuUdzwDsKIIuvX/YO
59eIM3XDI1gVWvEOm1S1WkT2B00N66cTSAmkR0lmYefFfxeV+AjOgRft8p6V2qQa3PwrA35v/oUe
fBfMyJmxq3G75QDNe9YqJtfzn1MExIUspfikRZKHLdxyt86TYTX3o1Q9I8mw8en6b3OR0B3JcA1C
6UyaEfPZaIIwGtWT+zoKGZzXersLJdbmyGLAko+sDqk8qPsZg+D3lTT//iFZijtsnQFVJu0n7zDS
+afDZMULQmVqvTX0lr/QkeRTMAa7O0lTQuf7ymkrLGAbFNFMmhhU4CWGlcfzZ+gmcZHkPLrkuXzn
o7ZPZdcQvCjc6pVXcI1dhZ+ktD7empLhY86LkyqawVkDpHqLX+nXb9KRDjxVbPGLsmdTPUlFonac
WS0ojRN/5SMjcg5hPXskVTeiN0hVvyALUwalcAaegt/Y3m2I8hN+e7vTnF9L6khypR5sVPOn2s9B
sCYxkLunm0tfb+rXckPg4eBRiLN0uLogI9Rw0+GHWAFxoYFQDwzv1GBBDXQPj51/dtBvGlqp+DJm
wTm55TB/vZDKrQSFS5qhrdGPAgGI9CPyyMrJYvdOYAcomAtD9W8HHhtysQMEgto+kPVbbAe3TK9D
1JOrpmVWLPwlsQDIqGTJq6hWvb6JGiuFJ139LKpAgS8cEynzIRG4OfuIjfw0QJGXzpOkGfyUT2dx
VzLY7HHclSrs28oLHaAL9APHQ3+FQ4gp+Cgd5s1ntP8X8q8EM0bl57hnaGFhKpiympL1SrnJbk6E
OtD594hRSSHlOZk2Xs1AU9BOemecxgzMj5hAPcK2gzdJsPE+e6oTeSl6rZ4BLjcqDArYdhtVoLZs
WtTam4SqG6nhxxkNEQpPUk2VxB/IwGFQEgC3mx0PzODA0ywAcdixU/Z+MOmGVaAfKbWE46p/2jfo
1/c43HnpHAZ0/Th9pcAzxC0I0Xgzyx0XBRNOglMSCkY4vv8F/Cvqn9oO8VJsfn23ZJs5NI7T0GEO
LJjdLol+TBqlVd0cD9yNbojIXtXdSU3RifYBb9/ociLG8FCdMo3UpaqBtqOvfvZySoVKFe/kNzBv
VgXojL8zlp+DrWaSOKoaA5OjoWbG49QhoLczuROeWlSVrUDZhJSMAzYhSXjLY3ONKI2nYSyc8S2W
4YE/E8fLlNeZC5hv3On/+3TPq5q9LU5zvu1j0ar/Gee3Q0j4GaBZ/N5eE9lHV0WFUEX8cKck8Erh
oUL9WDSCdIKbZ03knyaw4SZ5gRZ3pEmGvFsFpT9jc4KgtHeK5SadoL952W0rpI7GwmaIIQGxyczK
uGpI6XQryt66+FZKPeXABK3tw6GmU0RMTUA/wdMOXqJVNAURWlIzIToNEQ06oM8oh8EfzDiPUYNb
Mxzkrlz+Lnc+XA6Yr/xUZ19qH4Bs0+1N0yRdEeAsrIl31cuUbsJf14skLAFzJn60Qu5LrjyTAQ/N
tb601EtUcVBWnDhZgHGObD/RogjFelTYtyBFEST9DWhRYppchuIB13lgz05wrbfhLDGz3FYqCI/B
8kyloYMOB47GznvrK7gTHftS1VGl8m5r4jdolI5YCfCefe/VPn9/FXTKQWBhoNcjLnFhASJ4QPNJ
JDib03nyo2FQKs/u4frWNX9kd9c+lM9B4WofK4EzugVv5aexlcRKGuTMNVzJqcvWM1yfxueESXtV
ipqTjfdXeOvT3TVuoCRROxlBof0lhADQ043JpIxxSincdm6PwNY0bcIf+hP5irl2+7rxXw1Pojun
t1Y4x2ytQp6zgoEA3QdCoh9bdB4kr3IE9Fb+v2fXpALG+PzlbNjw/mzOnhvdesAITczNSf3lKP8J
ptSiYXn3aZjoPhraQoshBHaPiELH97ThnmnXD2TS2mQWJGj+F+DYztQbh7pJ5gQkOWK4VEs8+Mw9
KGYKH8YxOou2APUvuiXEf5XyeTpUUz1CH1+U4R6h4YhrjgrLvC3TA85mX10ySoWevIulgaCsI0Aq
B27qDIiBcDdcj6Y2AGYhTYtx6xzlQVsGebHGculK0w/LFjqIP+a0gJUNdLIYR2ZJnPnp/QR3heGd
sMjnvXQIfdDJcwS4NkgZieuNMFixdQbd0uNCWf0DfmCRWVpr2xySM2kUOqHt/q8hq7UBioMPoA4/
ZQyvF7t/mZhglt8CwEkpRjIV6VjBDcLIWBLF1uvCHGn3oSRV7iVbbRMRbD5OiqKo3s4CuRUadwpO
MjZ9IabCwHMyfwsoab+ipRIsV4GGkIl82sF0sPFIJN3Uvcek1wgPnI0xcy3zjbAEPDrZi0he0fbk
KXwlekw5p8ErH40iGfAmt4wtzWg96/OPdjgBrHod5yE584+tbVwhM1SlvIoQClg5AUwvncilLGNv
pjH/fB6IvcMaEYeMHU4npbHutO6+mG0CkWbANpMscXZu48nT1T8kfUQNYx4yio0s9rUlCxY5XOZC
yyUXUKYcdRBiU8mQlN/p2Z6N5OnPIw4wwxYx0IQnwdPa2cJI/GoXgricDF8zZwn6yRmkGcRes28n
U/cgnDvr4gT9UBmYgQo58w4AHWiplOTZGoMcu+BbR1tZ7Y9+AV6Cy+N7P5RCxzG2XnGJb+z+WAgh
NXFhY7br3o3Hjk53jARlLEGnWMp1c9e6IJJav0ly+usdsKUgI5SFwRUqdDkDBDLbcmfyBgkfS5Gc
3F8LsrQy6fzSk9lJVYFnwzv7DXzPd+6zC4mKPJQlh/4KeR5yzfGXo1zmmWgG0mPsXXtRnhxWCPk3
uG/5twOsffC6cvmNlrTIab4UHjpDE3/4ulCxSO/eox1GAYJ7mieu+tu1RqRIbdm3jcV8G+lshXP7
V70aEFQAWK08SwMSQ4S5UHJHxJRdGfiDMOUjnH/uMIvMRvm0XZaoHlVyMrsJRFQ0+3ocJYCPxMOS
bLSQF/k05tHzgV5zHLfzJagQ4/k/yPMPJEwvMbk1MLr6rViAYLsX3V6OcuyenrWxIH2cwnHHUfke
z9IDBUyqpt4rHUJvu48pgUnb0cw9Z/4iV4J/JHmEC45l7j+ZKKc/aO3lnlzhys90VR5JUE2gWciw
VzbWDcifNRx5pezAfLmsgQaHyFS0VkBLNlD4h84FmV2sWZqB5BoOSrskVLhj1c9ZnA1ERuJHVv8d
HDkeVML6EGNE+GISoY/ClMBeaK2/u4oTYZAP7PJccUPgJU+3I4dRdTFjlwUBA51ybJkqwT2JgTYx
LYGo9zFTumpy91aEwCCaWIGwbubAkP0YprmK+iGGb6Cn4JRcwqBlutILpOQ58Whbh985UbX1H0Qd
uK/Mz0gG68eWJIpsVE5vb/5y/7PcLCLnIF6jn+D4Pq50TZIIYRX6k3YUIxWQ6V7avhEhpQoZB6kF
1XcF9Lx0oH7zUCrw9RDKZJlbuL8dGPPfddN0sqytywgzS3kyeczGc8kXqlAgUC2qTm4KexqX1oo+
l6iqk+BBHxvTaG6W2N3W+UK1d1A+3KhtPYxviN43xJOBQ0oMVHClXGuB0SYaZSnNFPiawZLpx16U
m1jQ7BeHvZLlXafCHM3vFiEkv5v7TQ0wpYCKYJ04HUPPZwi2agBYrfnHnz1tYMvaiUJmJGsqt5lP
dM7F7kdlT7YrwpV7L+ZBwfVhY+VTiuNztJmvWFcJH4m2n40qYaoA/8KuUhH4Xow1CrgYudqdDR3e
WW9oeRl37DqVohksMWj41nsNzu5izmscQq34lx6LAaOit6+og5nEbz2sBGoA4hA85aniCBcbpenO
2YzJ30VUFhOKwZgmnwzdN7bFEJAB+2/kLIagv53StzqhYRuE1MAjpN+mDTKLB7uDxkVZ7RZUBECy
1ktNJyT0vDF3Py3uhYkarNkjXkphUZsf2Giy7YyH/DugcxGrfaysuT16rblQZyJ0HBvBjaPDC1aD
iE97I8omg2pLzAmjtgUH/7MvFWciU+bEkL9abV1tTt+ng1Aq6EF7vts5JxbpRJG/J4JsjSu4TVhZ
L6wI8AFW+BwDISNIlWj08EFXeWoit1GajKCiLDGtcLdOLl/RlSh7Im5hdxIieheg0y6aiAgstd27
BmZ0gYW19E/1YiQjfyDjqtnBOThll/PzPOYFIMEB1LpzaOgaTebVGIM1H8RFocJXAvPrkeJ/+SJZ
G15WKfM9bSGXCXdgMMvWTmzi8cRUxWltdB3RjO+hFsI4Xqtb0qbqh3ktaaeDWI1ksWDk4ilJ3zDm
ekji5O3BGi5JRcizDJaxy7296szJ8XPZccElveOSgvm/bH1kd+v5GIsGayxLZ4hrv4ILbuBCVVxF
VVOm4HDrrCky7NBcW6mE9xqkxK/OfcsgM9Sb6mwCfZhpS903DrVUnF2O6ez35jwvQiUKYUhbs6za
AGaHqCJoCkX7BqkoOGmPxlSQJwKdusq7ArEjS03pyICUuUeTGcOF7FydHspVR5AlnjCkJMSQgBO7
PifWONPzmPmHw1H0jkNqhexnhqHUhexbziA1gBIxFiMpqJkobVsnH5W19JHqoclGpcH1BsbULqhD
dlgUFlTnAuP9Ng1z8WFku0bHn5Gg9USRy7gwniI28IqXtXNEUMzrzKL0c12vVP4PmUttpxZlQ6gr
HsyrdblDFgLNlspxA+KBrxJ/bvWz0Uh96/HN7Wrgxe97aWU6woSCkLFfU+J+NnpGJUdxtlUxen0d
TjdgGxeDkRg4KHOPQ0GX1N2Zj/hbX2PED4eJNh2RnkRHR6VLyUjqjsCdv8ozMkMmo9b3W81HR9CE
3VhsqgtlXPP4vh2yLXxhHusaBlPvfpu/EhUXatOqn18ci1EJh+SgHzaU0YrsR6uiXaZCtBLpPiKk
PRlpaTFs+/vpVtv1Yf+TXLY6YmhiWy0jAMy2l2dlCdthdAwB43a4fp/GydhBq0wKjD6auVcefiPd
1y04gLlxLYOYVuYHGR9V2nSQYbbk9X87XIrKY7EmvLqrCIhjQWzvxIAowPH+SYAtUjJhcmOHLNtv
pp1LNMdZ4pwKiB59NOytfD5w7Ixj2HlQK4D3yaUPiKFeLW39Mn/2O8kRkQJQEo2/zIVIUTJKfQDs
MZACWlpZDaXpz/POLZHIH2KkH8Wnur+nwJc1XcZ/xPsABTGaFi13bnoMa+38sdL+FwCMkFHGuKp1
ZpkcOkt45Td7UzbrSx3UmsJLx+ZrKzKBb00vTlnK+OEIXEAdLpq4KEn+tudRo75q6NG91pPqDgCI
pIUFA5uKOmeLY+L5ZSKoIiNKr6UdeOVzzx+J6c8/5BK4OjEI9iQM06Uz1gtdVU9QF5tGADuYD7si
GxGQtXVtDG2tlXBjQBSNsCnsmaaCFVhIS3xjxyoc1H9ft2+qxo+UfUL9bMwA7CWsvmdRqcAqeoKe
5bHhUyAfGeqOID+mns9PWvAiIXqAb9tLEc6Vsle6pbTp38Gseq26f5l8zVQu6em2KUpgyy5355uh
005F6EXwlgrZZYL6ZUFax/21sN+gYOR/OiSFSV3GoMZlZfJchoYg/CL56K0pve1w4RmdUaBX5kp4
CNFbf9YFCaXmzf0Z8AWp3Y0tymjrHkHu0gDP1dFnhZjXFOUvtHZ+NyhWikZCUNXWytx6mt28mJUf
9tKbUGyEdixtwM2CsJMl0kgblzI0gAtwC8FbZj/QPO9tQFfJHUP2ArrjbHM35N3i4qriv0jDzjf3
hIIRnUCAUXD3ezyvP97vLznWwygyxWnwMtiJpUW33/zVSa/ABSHsKWKSf8dwAegg6FOvJhGMy+sv
l5h9u/HEwsrkTJ5hnHtpXr5TnYcH0AcK5Am93xNKt/637MooYsNwtCGSBogpJ9FyFmtKHr/trrKI
+1wzmklKecPyrKsZw1+JT61xbfGnV3TVnZDV2BrysF3wPqrt4DUekULjma4n8Jrzu5FowyEcdnP/
ZZNDwPHOeU3sTueAlaYHxEJ/LwGf8bKa8jYPBYr5vFAEyDslgTi0Lsr/+OxmULF0euIUaS4zhgks
abtpd+7n7Qq8gINpx4cGk2I7QRBFRfVwLENqKJHPmKXg+rNVW258bXzVanvTdFPJrkJnkwTZ/usH
88nCdccDZJzb8TxiczvvgYLwyOH4EnnS3yZ5USqSKT/f7YvJ/UiGg6TVWRWStql7DCHaI7aE75Cl
aS3/WitI52X0dXJg38G3os/h8J1yVCeIx4+uz2MakZR18e54+tdmPRMWGKyc7xfDGMQHgmUcPCHj
BzYtCgT6SMiD7QZ4mJ0LpEzZoF+Cx6g+Wdube/w/icWNQNU6QWQv+u81kaizJkZ0wwAHFWhEplSk
n2GHNTEq62l1yICJ1ed32iEnI4k5CCbwbr+FLRh9cxo5GnRVar66mbfaXd79uFYIqMeBIqz7yOt9
8IAwpxLgUpmGBtjFLMUOOnDIg6VWBXhQBcgtxXsC5/GkoSEG25ud09emLRWXTeIm3oOaEJfjWuS3
WAe+SbXSaXuGJCNWSmvWqv47f06q2vRRMWToWPaoy9woOCHXkgrsAAvzFdTR3VAUOq11Hu5sK1ob
VspF5vehEplA7tzYxIcgsknLf/SBUKs70cdC527aZ7uLgkxsPh3ZJmKZV07jSSnPrx9Bkr0KSaSI
kSLRtv93OEKLK+LkkFbB4JTbo24UtEXQaK3IuTCaukDq+7hI7+lauh5/aq0oKwCevlYEchgbhexc
bGXRz18R9ZxQiXVaPRXrhqB0Z/Gtbhc2h/gPOfzaq0wN9tqy0tpLENzLIZW02UDvVIkebsEmTPnk
3Cy9H0vUY/VXZEutIfECsFahLQrS5DvWld+rnjSDolzfasYCQZg0+O6wGNUpzIfQNYBMkMLuni7a
WAXT3GKh4/2ioUGkjZleJgM57loyjfV9nXsH4eSHFHiqQbkSYx3uUtmGp5u0HAmQ5Lfjp1ycS9xQ
eQO7EMB+nLPSoWek7crW3sJrtY3x0hCJNQzvM2iZJ5uKQBq2r22wkJqowjIOJbVgFA5ipoeLBa/Z
gxftXIUQx7Hfb2Lvv9HMMnk4FrKOp9ab6ewOTigecZDkmgXGrReX7lCGCjkqOJh4xxoXbbpS/H1C
uUOAlzVGA2N+VbqTJXFjTkgej7omTkw5Xn8zUnAyBl/WqXs+gE7z7V/nD2f+n+UFC5Ad3DUbYoj3
E/9TXbtjOPk8pc36qUqfqfgMiiNbmh2sLnqaBJrFTloG52Nd7fNl7FjqJK3IyYpX4fFY0DgKJk7b
4ZprcvQl2fMGnnNIvLOWSUUVdRk7fj343YzUvmVdrTaa6wrfXcvQW1w6oRm7y2WO3+smnMKigEXR
Gd0I/3HIQ2Zsi0seoxlNiLbzB97MLnCOFLeb2Etcd5XGjL2/wqPi7++NV3hLkGJpx3EYrbqWrWOq
W1V/8MeeaxmE/+i2k8aNUip24viNrtFmEGSF39T9+HvqeGxNPMLUU8/mC9TE+tM+N54ir9W25+bu
dY/hA8Ombg47JxOpRuxNqT1qOvGkm/xmBLXQFDI3IB64AA5cT2Nuu4swutIbRXJ7ky8Uy65P3XgE
9PslCI/iayyhPZmca1TFAIVQfh+p1P0eenKFK+XWb00ykgIhUG31g8oQTabingyFwA7lOo5VuzuE
ZIDthTStKKnfwJnzvL686K5f5lv5gp/RYMdsOKrH8k5G6qOjYigJ25l7NHasCyZkt9PyQ9mWBLqA
glrT44Pvs9GaCwH2ak2ot6GQk++33QV2MI6DwRfpwos1ko4Twqi0gIw6VFFQwmngtuCAXqT+33Gj
AZSMZlIS4/zUj9IJHPJ/oieEcun2CRajrp2oQa6yTiyMf+jnqwii2QOJzZciFJU01Ztf9QrT9938
GlvXbSu5wJeZCdFcm5xzaoFoAGniPI/qkwxTxUk4uBjDtPh3gEWPHGlpK3nh1kjYId3x6l2KTel6
aN2u1Q2ab28CZ3i4kNz9kVzSM6FztI2eSNzPFIWuMb8yTvTy+CdCzVHmDPOkTNNUnMYv/Jf1phc/
muyh/xDZ+LoxL4i3Rpxq4EMfcZnDkL4G6IrwJe5rlsBf1bzCInkY8p56R1BvA0lShXhWvm2iPRrI
Gv/eWgtyDvq/NY2wpunpYol7cNt20hc0B3ZSGMNn04cjYU8/HWwsdB7GwZSLdthVIBIBZQOohAOH
w1Zk8fDM89lq0Ctdkzw1pfFMmcrekKqYvMCfGLO7JwFZl4B2E8WoHqPFeSVLX4J7+FCfemBU2Id8
rIsZOncmUtWVjha/+pZnZ1vsxe+FT+UpbHqgBKeLLi5ajU7MdL0X8IhoJKwocaP9H/rYXTpCwZST
HTn4Y7TC47uZBVVzKHyCY4EoUbRqCkAS3bV0tYjwE/6jMetM1sfMlgFIBGKzasstCp5KgG0RiQkD
JT9/ihMZKVgn9VzFhzuQEc4PWI0Jk53WOK4jdpUaojaSPcCwQixj6VxCijpuiXOaxFzDaetV4nF2
maGbAOV7DnD+G0YVgPzbnaM2+EONgdENCq6DJsc/5tsC9dq9p2Jil7YQaVtHXaBQ4oxznGSNTLgr
vrJ81zMjcY0W/nFUxQ2GoTdTmyUmUOWjduwyfbXuqAdrOOUsUDpdrkHx6o5R+jtuShEt4TmKonK+
JViFI73KrHA0vVLMlsHoxSedBS5Uv3utRgsfGc7sCqQ8AgnT7XEbGlPXx9FURKzWBN6fM1CvJU1z
+vRiryG9wLJKnv3UL1s1TW5bIbb/hqHeMVxm+aqQcA2pZUzR44OH2zyl3w5WRMhj23YoD2d22tCQ
rzXCZ0Q2pIBIZw2B53GN7fOg0oqzAtx7snlmvO33RwK1isGIbQGX7Jd46gzN1wjMzEElB32rYxTy
42xiETg4MyZNtM7M6aAe/P5Qcwd9b93RiVNbGhXEss48eL2YRif/lXnsieXsy0ern98sZoMv71vg
bXDQ58bCtkqe+wba49+vPTB8cRF5pSGfzIwfFSfcGlOPez2Z7iPNHOotqhc740Jb4ZdoBLkjmGBZ
Z9rahQOq2zv2XcGCCSMUtVpVm6LK6rgYEgV8LuvWoyhuwY0AlVWZpLyufvFAda9/HGk/NoxfVNae
qPt7AfZkjQiBQrZpr+6A6pVpWvuYP0ZpsJ+BaP2qEQPr6GVkXGzQzBxj/Ln4yD3uwgGsvz7uRDxL
LDEr8rIJfSy5amHO77diXwRgVtwS/FNSFkSmSjIh2Ze9pyL9InkV7/UMgFZqNI7RM0aZHQ5cc39t
RQ1MYDwVP51Lx8TmkcB8n0BmAGiLJuYKrS6rgPxwr4yf1wOfQOQ+MWauy1rHEMdCgVih7mNFD70/
Mo+KKrjIRj9cKqSH+T9yfYg7isC3JkNLXajsf708xohEK8ushSyNfqpSGfPwpmm39ghNhq63dZmD
ltDY1xuL6cYsyMBJRqDRips+isEuzi7zPICsNHBnE3ffR24GKn+ye8jJnwmVDAWSdM7LskGyBKoT
rnCHXLKJVFfDAtYZJuFiRsP9FSwEN383cEZdBCyuscjXrvWW0bvyEoCRrw4iyAiepGFyGlCFvvQQ
5z0JCh3f+AsOaMYxiqhqJrRf9A2zHkt6hby9v+zRftDn2VcTKLnIkYL+cVru028N3Bz76cWRCj17
4+3X4KPZ6KwYtyXtpJ4kpoShEjUKKtfKF7GzlIqbSRWEdEgKh+CojMhw7MyXA1zIt+4C3fd/e6rv
EmeUYs41gRLC13duMZZV7OKVmTwVRRJ2s2EEXk5+XRehUWDMzEBHmbAhISUAQg/zMNZtzR3tR1Dq
ZDdOHcI202Plo+pU/S690jD82FZDXCS0EMzzc1xmcsQp/F6iIhSPhZBJd9dzaAH8glK+lP/qMoOv
6Bx9bM0nT4lZXaYY99jX+Mwfz9suOpV4BMmU+UQ85LTiA8zKOymfWMWplDm6aJFkNymE6NFA4ZCh
Shih7GyNt2MvwU5SB8HSnjE6Ek/3v3I3xkS9Mx53Kl9sj+1vD8Wnihi6ErAsecUle0Dii5OLpqmF
gGw7afXiWJsdGuakiwGi8jP8BDMPXJ+vYv77WlzUasKVPIVsMIVEjmGAtUIXRBRDn+p9Cxbe/cfg
CZgZW4ouMHnn6Ko9ZHP9QEm1lzg4Hoc1R7sV7bGc3t1v6kUxriREIokepjo87K2znmYIjcFJrwcc
6jHV+D1NmjakDmIlWvjWlTrksLCAEPpjtPSeTS6DPY8BvTsNv9k8A5dz5282GNryFd4pDZDZkPTJ
OhCytatGfEJ0H/Mj9l1HdL/jLohMkJmhJLuDfgyhhoId/6AmdWQ7yFjk1P3f6OidJcyfK3vLPwlE
gkFOQ/iQ1GKzsxSDHq6TI5mXEr1AlJWPzS4gnMSD86uz5lfetvPJugXKwjq9+ZhPnhpqy5d/i4nL
7bfvUPwMGNLBxijjH22tlcT9NhVoRsGaepXShFLmSelfBNauz3UemrMTmw33+W6S0Kr7jNXmP78M
vW8gnGEmFYwhAiV7gVE8jzxFpXbe5UpMKJfjBnJjHhzIynJphGj5xojmI55bJoubrcASboaqjUPz
E2cYjs1f90IaAh46T2LT/7eVAZOuF4ctWUGXhpjoj+hI+rrB+ffWye9CSz308kSA3H7qUA6Q7mlx
Inc8CSVF533GtdHrEMngkEipk4+R0MeN011hwYE+oLokNTNdv+Kx0SXSix/YhpiGesso7bMxba5i
X26RLWHQuG2V9Jn4ndFaqbr2wQLI9T4vlfs8zykTXt9Y4ikgc/kI1+HNJbd8thhTjPW3GMsKBH2P
6eTzPnASL4ni3PFsCMnMCN5veezpY63jsp/WKRyPG5UPlCpHgomn8902LkEDcz6Tp25+2lzlF8kV
kzy9DYWGqFXx47RjcCreOpnNc0Hd8pNDHwKldCTUzhlknXiZQG96EXZZSpj4pbvfWdavHuhY4ZGS
eW1MwGe7ZMyIvHZebMUNVpnfzzRZjo1cQzEER4NFqHBOJRioPTUJ12wQXNepVhmVi2XRgPwZO9Wh
pqmEi3+bY2cE6s/T7gKPqjipCJsAXfCjkofO9Oap4M+iSDbt6pSD1Ee7MBsFy1xI3jo2uwtO8gSw
aVm+yYJyHW0m7xjNrqvi4PSuCyv+qPF0xaQ9Vr2BipLhxFWHbXMpyXNQLXf6iCjBHlNZD0d4dfQ8
x8/Ce6uo9p0pYMJf/hOcSW8LU6norINuVCvJz9ysz6ss32HRWTlMDtUp2qHKR+t9kWKT0ZgfW8eq
a/9BmLWMGr2fOHBJE0PgNgZHPPwaKlVEziW3bwDfQkkwBsJ+X+MR0oOtZTeVZOsOqqyBsLFM67NV
1ZRMyRB49ytuGC33GoXjLWX/qtgZ9CguJ6cqbkPi7zoKX8Tcsbo5E/dXUecKODORsRMMihuHjNco
Z1u4MuE7uY+/VCj1c5tW1WVhIrTt7o3BJy9YkPxlMbiz2KCObLhpx9kK+6mH+l++c+YQkpgvC+fG
GvtYiLWrLBlGyD6BPRAvVfJ1ZxKfe0WVTs0l0iWgl6J/7b7eww9bG87/SS2fjNdJ09gr5qjAjwRg
B7cQcdL83ssiDORsPDlJ2UGqfXVM5wVUWiUPPfcCkior0Fz5CR1+Uu4H/2QQR4c8Jf5kXpb1SVIx
DGGyB8W2m9mTdEjHiDSCaZJIUFEg7lwrg1KUFqttwvyfJ1wnxhVJZ8lYrHLWMPCNdFZqPGyMZWlR
0EudrMcrMZIBH4hh/D3LZ1ZL0DSz/QYNey7pthV9DytEw/YM98kZFUkT6qI+KyGapxkSuR/ReHVG
aBjU/nmMQxI5/jIaMdFj/1pPIgADIDv0LHbSDV8lJhErvsvOzOCp+ja9P1APa8ToRmx+bZbGgz+O
ztku7CV8or6qsobE9R0jN1iVFPxXtDtIJgFp+Rqy3pFOcwzl+1IbdXTTOu44vW7FBoBPwQgr4SYN
K9r1hxiMDGmY42NYv65RVA/J9LulfTvKlMJIkvVBvBiQgBah8VjR3htYOtiDqUfmPctN92wSbo6y
LDLfiOmYS/7C78xD/FEX+kInMRA+1VWYHDxekMvItasSeCLhuUJx5yCBY7CGctremCqxJkuXsFl9
1Xfjq6GJdLzjzLouHaMVuPhUW8dDwWXMM34hnEnlUebq+wJgUhy2hW/yeObqRzWOy+8PWpMA09RA
tPfjpxjy0ZU82ECe5GculbC5BtLA5K7OfcerTDNB3fyIps/43puklt2j1cXv1gqu3jM9pi91awOz
7jvFkGGsTgppfMyX+eEagVbEuboZ6PQ/an91sEoaPJrByQBMidHm+6gzGVDNUygKD1d/7xTnd+aB
emjY3dy9AzroBW05oE1oXo9QC61nTprIFevABKuUno/RngLX4+4mWlUsiEicniRGSByOgtEWNNPT
CpzGiWMBeNgNrSY3X/H2n/9TH1sfDSTCzx70SgSxXXyVodldjW9bDyM8q4jZH+DdSZf+AYM+Bfhj
Cl+UmTrzjmxB6mG7AU0RXUDw/VZFzyR5gVJ5xGeM+MNETM45EvtMz/pdBnVN5tMV8XbxWLqWOBtJ
6kKP74vr7gwOVRHOuyVMe+bdlb3HkuFr0OjmB/v0fiVPEOL3dTKYNhslKtQro9WQlM0w2x75WcZe
wQC6hYXQinoyJXE0q442wYImxROG537xRCfFG+AZIgZVHNxRGeaez74BrXxU+R+SZ+pg0Jv7xtQp
FvPJ0rjWv8JW5m0kUy9nskwpr3U3epy14qzdekr1hGaq4ZNCNqXcyd8YXwzIimAIyKABVMzPfhnn
sdUSx/tKa17TEx7O9keLL8x9Iq1X2Z5GONAP6eoAqQqiP0Jb/nUDQZ1R7Kgq5e9ZJYJ/9MAFr7Zi
WYPBankQ5o97gUSK/ZW9HkGlHnfqNCUe60ENk52Nar+70l4KFQ8oDoMIxnnZR/Ep3FgL/Cte6AnN
ccn8+l0DxyVijvqn3OAfdgKCcmCzox10zKVE+TbPrcl9KmzCy98zKEQvRXcqtiP2S0Mdudy+EOiQ
xe0oHRzVqc13YTHeVZNNBdtoiX7Q4uTTbqdBsInrWAU1cgWxpkagJSlTQCNyyZsiEcywT758CjHS
nlpPj2Sd35Py3B+Efutb4WNbJZCehz96OjrwdzLPbZ9RKqm1H9jiCgR7SRTquCDmA5ZZ1XL+XPOW
pd3Z9xiRmzIwu2eRDF78TwQL5n77ubjiYd8MTPi3RMxHUCif+JKk3ZsTwvdHvTFl9HgAhKDLHuDa
gwlkjnGpGVnPffQyZ4CXLqJYZg6SyqAgJTaOP1vjOGbnmIPTMse7XcjXKetNBISCdBln5iP44JyO
sO9+XQiHuIjnLT66KHdC1SaG2rPPP/HkJkX4LhVgHEXDMMmaQiMO2BI9TZYoAqhFiMvPLuAXIfZD
pSzHyVAXwsz0cw2YmK+m4p6y8+v2NlHpQMtL9ZDkkLdyWcAQWmyEUZODc8kC2b21EnqAa5uATMD4
iduPUGqn0vMViOQgWnGJ9hswnyjULe3DG1CKRAj1cLFHzAWtYEM4hkjjf9SE5HWMvwrco18NVrUk
/ZCVHLDa7wvqEjm0TchxxSHgE4aoVDS4XUdG8xfv4rpd3rUPdYMdlZIo5JQ/8ZH8t8B/nsb1llaM
ltxHF0eqKHSU2ygW7VI6Y0Ty4/xig0rQsOGu5oxVHElVggtt85tNTB3yh9tOjkQHOVrNMqcJ5WGv
JsVeL40ZD3wKx1o5euKj0vjl+FEm6gzfIkGg0czpKhCkwlH/NxcKHqC5wK8ezhYGvvHkBVwGlnPP
x7li/d3y3MMK9PQcNtS0YtOzsoO/cX8SNhHoV46AtRKHJzXsTX0ima9tSr2YT5VD3FOWQ8Y6VuiV
0SvziMnPTGEvkUqHhlfIud2lvkiwORnbh0PPJZpLh/Br96M+2z38515H5OKLeBVcNphUmrn7cHP0
XL3Z/ZRABJQJnHzhF9iQwtMBH0IXeA3dYC2xI25mhwM5hyctzVxi5qcJt4MnBpQPZR61KaoCw9wQ
v7rAHXgDoY/geKyw0HSc8m/KIz5x9y+kMu3aBqQ6fhRm0k7b3V+IM/ReZo/NKs01H8STj3LbO5T0
+Sysc9KJN9KU97jbiOtHl2DD8zm1F1NieYKWjJuXavwQE/jdA7GDceJtWJaxg3tLD1Tjxv1Mp/kn
yO+M2xLxmUmGFblIRif679hlCu6+bx4Xvhy53R07mnWvetl4hEBAmiHmgd4qauT7BLx8j5kT6az8
b14odxFicEOnniJZGu7ePf3z3Bvovvm3TV/cPixbbqoHvhLUjzwqWoj+tng+mHqgQdJL8Qa0SPTO
csksPTWCbaC+zNcfHsdN1y00GilYyDiQh9uFyTXlcrIwbptI1C0hYcXs6pRtc832XM7qHGJPAfHt
hPtDJevFWdbxGCQIhKWtqZ620kE2BXn5WVa0pMYLxEsZaUqylS+GBCa9MixB1ZnfCeDG7QmZkwjk
vGuevzLa02C+0Z8NXCbyyOp2s7jsiO/8gvMEpPuN1/+tXs1KK+T2P2/ZbDFIhk6DBYnI5jsqpgid
DIe1kqgwebrcqxp/iZi0hTJhPndLbe+nWSyhliPgX74GiQQ3kuNOC36oKbiwnWMFNeKEvtvfKHLh
UnriVPQkk4cjJlzkX/kVsMucxnghjnFXRWP8IRHQOtaO0Sj69JrAUn4Sire66nZ7P5vWyJfAsOZ8
T8tuetakPs/g6sFR3kCv280+DrIZ0sf1xxbRuC+K73HMNut+9d/TDXEj/YiYrbOPmelCT9X6e2kq
yXO5VgDck/eaEeeKCWcHTnA8HuP7nl1v6O7zIWA/FAkKu1pcrAYiFNYK+0BY4/AZFNi7djAxw95/
nj4LIry84C5Kn9s+oRLh7y5C80lS9l314/Ja3Hxt+ShOTS/oeZjWlyQviJWhj3RvkdE1px7nqXwA
Qp16qCjN4ZT87r526cvY03ymE+c3SvOUmGizB8Bc/aaWQ0XE/+k5WFam91lt76nz7w/T92fIvOjk
0E7B5Yjjufd9HbsmsORJSwjTcOPykPrjKuz4n3OESjnt/nhf1NdYjcFXGdIKemiYMkP0IU0bWMCg
qS755I3DZLU49cULirrSY2KDgYqN0fbZom9u67g4PuT0XKCnjD4G4WC/XAVb2ApADodg0+zoGgvy
zs0cB/X8mUnNKC5KSvblDg8Eo8/ndIzLrdLVzho6YZOJQDwtvcWipMUzbwwLEfc8WQ/AQCdocnXQ
JuBCm/EurMwc7oQKkeJq6LCytpg+UcD2qZH3aNutBaAKUjmjKBs6nUewAZoXINgSMyzUS2UgM2h6
cpcWUawE16lDlc9P36gVHs3ZgCi7D7MMqr2Nq0xemd1jlMEoRs1kTkYhsMXzFGqTMVQBNo+2fi3H
FZbxU2GMjuGsORDYYPHdNurux6Q+g86Q5d+3PDlD2on5WxXqegULxeozANP++nwVqonxlDP/HYjC
XcANNeW6BeE3T1UUO710gI1FOfv36xkU88e3IWMK1zDmI6tOJoXQFLzXzvWwrJm6M60xV/f9kuH7
Z0GGqU6b21QZJoeR9dABg09yL4AhenyeUSkPXJqcOKiWI+x/HcukUuaffz1ZHa5NAmY/t7KKY459
dFSWY2gWg6jrid8O+XnQDZKdgaBmq9Bh+Q5JzorWqW9tspllQ2NrYMIctgYiUcWxIsL0fzCYAjIF
P64irJYnwLfNAdmOfuO362d4Zm9CgnMSSxeHadYQTvSfKl0eGCVXTWVN6sBmqbkM1MMiIBH4fIjm
NemzhD+rKLI4OVfxrjNpEyBoHT+AyQpUS+WZHt7yuqstp4MrTKVKNt+R0kLm90NNbziTSdRaEhz3
MJqEHhokO1+tC9eVqbd4+1BAiW2X8Nmxil4ap8FeQzvRx8PPTGVCLXkeQTH2a1zUIfezya+tgV+1
B/AroU49+WWUQDBaH3CqGiz63CfymPm8idgUHox8GppyJl5oni29aXOEXn7ceEoeg8rh+alSlmXI
j/XNrdG3zoDip/HFqodSZlEFH85s4WLJ2i5ph3QeQdFgcKioTccQLypmER5UUVk7nYoIR2Nh5Pd+
TGdJaa4Kop5EZJp79HDo+QczxI2i+qvrv6KLQYRnb1GLiwMI4+X3PTCUdDAic7YJrwdW7NC6Cu49
g27ehC0wJt9KoMicrbvtIVBrt1lys0qHhEzmuNceMJ8r0ZJIcOQBpW7tIrUTHY5rmdUcxB+uy2B+
tj+2CSa/7ooBe+4ERt2ONBYghbzJn/gjxU7DoBDJxweeAT6mj30PwqA1G0SVajVtE9nyVV1mDd+u
ed2EuPU5/5QjDzFGrzzYcg1mDi2oaYRUxoCZeqQl6GoFTcn3gwfuPqjmsx2HKWPfo+9q2yIyAUm/
4UV886FxZj+5TarQOJbl47MSRV78O4PEX6mFkfi9hBj05MI/l8bbXBZk+siAXrZCcN7YE13Wj5Al
w/cmlUz0xPia7oOJkue66NJ7NqFPgc8bJM5+eaHhYlvzWQ7u7k7XMlr0UI52Kx+sWtuUsDL/ooz5
RV7qnuHgkjD99rg95AR0GoHl15Q6VOOjEtja9Pk22mZEoVe8HdhVdHCHbn3X4Ko4ARFYvoVeDvfh
b1hc/2vAr7cRHYVKP0lYDmNUFUa+P7aN2lokzVdJrSZAgiJpzbRxl5Ro+l8zIJLM4EYI0mbuPHoF
k+Xoi5fatvk8izncKRfFKAv3Uull4uGNpFx1Ge9GQ09XWsnrgRSN7YpdDY56IfnNvvS+pjEpL1Uj
CI4VYi+YW2HijKn0cQjSWXfH2etsXLLBndvN92c5JKIYJvkYDs+v266CqMmnzCFPEon3kgo7G/tz
txkcSFhEjnk38me5bmEP1/0cZ1vZrQarHYPif5L9z2VMz5GsnnvWXxqPnBvFupx0hMzF5vm9N074
lbojECF4IqTSgtBjqIKwNfScZxd5LmydWMEvdKsu8MezGD9CQhcpbL/aQqNmt4fDl0CQzr+rfpT0
GX2gmiUS56l03/4Cg0fefNtu8tB/0PAmb4iE5H0T130m2fcgxTh29lwckcYQpjOA74yWJJhSakw3
KcUrQJ/b21ze1a6lQ9HyK1UP2PHi6gM7tH+cVvFIkJQz1QrN6GezPZqy7t3KM/HVTnDcorAzdJN2
nv7xXIMpjEq4djQ+xpQxg6lzyUPiaBRmpQwOYZiiQgSpO6zqCO55C+ii2xkrgbpb40PgcHL1sfaD
0vaDTSoQiOCtkIFi1yFgkITzqy7DQARcfejTgRocJHvEjcZ2vbjTtBb3mkpq6j/3Sp//EVRBLkhq
+0IC2ROq9MZVZe0HUQwOBUSBUGElFCTa4p14zg9hIljmNUX1jjKqAC1O5SAvdHQEt+NvfhBqaS9O
9R6aWsQg2mg0aR1N9are9O1Z4kF40s+xEaTrUYCRKZHAqW3YlXFbVeveya8uIh/5AwdEo1z9K1aB
H2jaO6aXr5W/R1rkchZZt4zFJUMG/qgWsMMDa9ve72qnDHIpB5ZYx7RdneG5fP9kAJIQREXOAbS9
c902gao27/NSjXGh/mXeIV6Zl+/wRO3RXJSu4zd9Ss/+zJLnmYQ4xY+tgPyRaK+VFaT8lx10Oidw
BmJZY3Duy9aoCcicyi+4V7WPNCeArumZ/OPg24vVg67ba03b4qVaRoMltONVzMMM//JInic9UbXG
0i0H0V+c30Hfgx5Q9vkCuBYykXSS2w2qpsRvFX9xzMsJWlUaAINSuqdx5FWZsrF0q3ZTELEhJctC
PnKwn1GnIu4TG8/Cgw0a2EcF3bdLW/pTjnwimdqNfFu7ORmo1LTty0SVHRsCKlHu/5gpvYPAJnq4
e6PmymZr+32NY9qxuYMe4+6Z4uZTfE1qkh8e65MJgmRCKl31QRij42n02V1w4kpln3rx7Dp4r0Xm
1PNsUqqcrLFWDat+PLrJp411CDyHWNSHPw0Ogofc5wdX1Nu3WNlwSbL6fNnI7y1LTYH75cqJK5wY
Etky4H66hO4Vn9RC92VRj7C1YxiE7p4Fcy4Fu1XU2k0Z7QRLNKb3dCw0RG/4mn7z9rDdGBHY+tkP
lpYPjq3l4XCEMh6CSF1/KpaVU6w78pcwsbjNpcRdMGrcTjl1zOCcbc6Kp5Cw3qQ+Fs+I/nIWHyIV
WFiY/eV0gLEgDM+ZYWgtx2B9ERgx3g/Y6emTNuym81RwqBwN0YBGHbxp9T1OD+t8OUudYe/676pg
ez+BPXY6xBEfXkuYXHd0mBdhqaG0K8UiP2P+fd/PqdVRI0tJwuDwBP1RgqcFAj3SeRkWWSPiYKLG
8bCSz0/uLMl3/PIoTLB2O5Pp/HskJgT7BlZKxQPTec0oxcVT3inEiqOSMQRjGoG2rPkaWXQ8X3x5
XmCo2IY+Qle0A0PUimrKvME18TB2bXz62VGazt3JFznuGIt7aUKLOekWins3fIXTMRAMqLCGeY42
B32xdAoVZGb79G11P570yqKJvneDSUg7rekKDdFkqn0/aHs+Pyr9OFSfipRSY2PI/sjnCGLRo2bR
kRLZ6RcSpsoXkEEgYO7ch34eT977E5sVY7iAoN+AXFuu56wGp1H1Htnx6KZI2NGZIlbv1ZTCHCvz
o/SXRyYNZr9nDk2ATYdwA+krOKaAT4Jm51tHYb6AmkRbzJ+7fQjK+78rzKT291jNzvfnVDj/rLQ4
UnQ1iQ49KVCQtbwP1G8cJ9kt/SGps0CRC918qEq5cNLjKLd3EP4ZPbZTeYBn1TzejrxGya9FQp5b
Q+fSAuZCgsthu+3BLiQWwpKNsReajQ0wXvx+4bJBoasw/LABdPtbS+RS2ppg/vJH6A0chrGGhRQ9
MQ0dn+DEl7Gtabhngx0ZFmrDDvcsFOEO99mm9YOxq86fas6i11WQ/kRDv4y+f6Pl1hvHvwUObL1m
s8JvG812zm0gnwOPeShzdbkptE8+rCWHGyu+TNx/jwR1klDJOUTmy2KjyYbc/BK0geaVo41e86h+
kiLgP1bf9zIM3CpD/OCaCBhTum7FeptRp3WzOc7AmkQEaKpGWmVeSbee7VYi9ltclA1BYwWWk4g7
OZd4uZ+WdMC+zl1CiWlmouSSjfbPT3PRkVdxq9VYoBMTE/qPjDRW5KRMwNrTP7kGVH5/zqY7ztEQ
0c/kYHXjJp5QUghncb1y212YNs8geGgaYu2NjuFwGgiOS5iqrQofHH9O+y7nUOBvj1ZiA6IGvoTI
WSS0hPMPX6vryOI3eTr54fZH6oJ+6c97EskDQdugSQp1RXDhLVu+idfI27hYr9I1SMzNuqwr6eVy
Nv1pktfRNNS1ji+uBIkjxGT++lV2snlzbSA7DwJRtUahpt0/ya0V07EaNK1Tyvc+mxPddLUvxCpD
YTbcnP8IcT2Us5BLIS71qo2Ukvd6it2ryPRl+ddGyhO4l/Ka3L9PY1ML2upcqopTOI0Bqi6Mlm8t
uIrmxOxF5f99uggFs1eK63XtvvH5bvv9OGJbhLrpVgQrMjMTxi5zTS1rCj76USnsBXp5xDmUkqJ+
Rf4sREVOAFTmt1LtHVhhUXCcdKEEMyCF+fX+SGG92wBX1kP8iJ/ZA8suz/bzycTiNSSm3DGluS/f
5LBgr1zT3GEfdfKrghRSWNz3FeqpnMbzWMVIaO5I6AIEgxypcY/aEw/VAOJIW1Mhh5K4wIlk9ijz
avaUL93Pe7IdfAykNq6LD1gttz6tTPA9drqo11dVD+bqDeg8TRJviIKEXkRSPEQpDnB51LxBVcCl
hWYmQsFbHL37ukOjbvHpecrymCxaqox5a66GLf8CaA2Mvpq7fiiZRZf+Mlx4o5hHMawsW00NABPo
rGFrBgcspShjQxpGGOyBZGgJttNtenC6y3n4pIAd4o7XY/B2rrkQCgFue4LuETCAfW5g8znO0kv0
UljRD5uwComnO4Md+c11JZIjMAk1x66pyFgqdclkLgdlWM4aQlFhb3dI1+cTNk3RiGMvkoTTs7tW
X6Q931EfoDtX0t+Yzskxl7/BobzURKYMBBSh/QYZJOI9bV8jLm+yaGNiVYXB98NtExWvD5S2quTo
xWtHDRZn1/WsNkOVOGAUmB+MexbIE0JuQDTUqNE2b7YyndUGfgNhrBp3aOwgNWCw8jth+fsDC0QV
XuDe6N7ViPqZvPupj7+iWEiMaaoIGOuYa7S2vUvg1yYSypMCHwYdwBhb3ZFDhndFqQzb6OSf07Qm
6fHBkqNwkalK1kifsd07E12XgPClPEqHA7dcKnM9FgshTvXORYbf7X2ivaz0KbvosH2+5u6Qx2H5
oCUBYazcqPVsfdhLUIYpE953D2N5KAC4wl2r88wqk41HNk6yLzwuX9isy9ZXgjdDyr6c7/JjiRWJ
KMd8+oTtq6vzfJgCu+rcUO43nXY01x6sPk21qryBrF4as1Kr1/KSxkmpEuwV2qV/RsgLZgY34fUM
kCkoz2SJ9CMOl8pKxDYeTt1dEm58yD+rVKEN+uZmKBk8SKJhNVaARtnZFVKLL2bGKv2WQT043F54
0oT4yyzv9gyWZWqssfg/RIlmblVlGBh8IuQoaFtpXHryL9mWZ8YyxDGr0uF15CCwtmfp0Uiq/9Cf
5dSIpT3VzFxGMnK9koBJy/UKYuZv2BTg9ch3Bjy4Gy692neyG2ZKSTYq8B5niwG8J/FE4jTohrhB
ASnPqf+y8cNT/+GfxBAms68GxsjFD6Pgo/uM5LkqDzlIrOw3UwhU6au8WpvB6TIzGRiBLk344Gsl
xfIug0US4vO3lU8RstYNNzSqaqvRJSpXLpE9/gXmod3n1UQ15/1Keuv1W3fHUNHgUQ/vFLEC7cp2
1CbwM7+wWHEefHlJqQo8fZsSRQ/Y6NnHaeIA4KA/lUsjngltgQKAOMOy8Ip4OzlN2e37q8u4aknZ
umMG32Knso1vzBeK+8C73rLnBGDns2sZzBrcOwRlDE5MbXmqn53oFQim3AJOb95LzJw9ahrotTxx
YYTrxrYxYv8KYTSLuy5hv9n0CY9YZ4Iw7ZC7pz/WhfEt6Q6rej/LK7Q3SzfyVZkvDR4rD0OGALtE
ZpNgsuazjNIGGS4zYS5IgpfKr5ydcRHdotfGtKCaA4qY3ceGYhmW4CdpA291qpdcQtO3USvabF8D
42CFc3MX6Ab3xmFKs5zhNrUcnPbhteACnWShGQLf88oAQ5vP+4TH2V/DrBidCW5f8n07FycEYcr5
U4AORn7rghEbpI+6x7QUZ9OrP1qtKzEaiYsI6mVis8ri2guWGVaBVJ7cCciWXQOvdd7UVOel1Nxn
x6NMLJA4O0PTOTfddWqTg6UciuPiVMiLF4WaCaI+oSHq01TIimKmvsL/2CcgV/5YD0xxToPspSxx
WRUGmVnRVrPK2sT9RiGZzZvAM/Jb6/WRAfxfc12lXJLTPbHjBvNe5rV4l2bcLoTub0e1fyM2MkK/
J1eOxqK9yjYMC9XtBE9O/M7fCwolVfTjzl3X6KWIIZFFLfI5BHYqnbWxxLWiQC91nk37FzrVuPh1
uFRTcHAp27dZFpsmr7B++0B8b1ARHHGvFJ2OdBKRe/6ZGA/83JwEFYvW6nMr9qFIQdC7o7QqxMCB
EY8BMTm2jxLHaEl2duUyrel5LAJndpCTOtvO7UrUgMwr5iUy68qAXeFPh9xksT7kQSG7/o7nV6pF
hM6VeZBgiPPmSn0GQgfGELuXJWEtO2b1m4d4Lf+1slJdd4Sz7Vjpg8LTNhuHJ+Yh/gngY4+uRhlY
Sm+2TKOnebMEgoHxlSar+6RicaeGQdB8TG2UQYkut6W1FHPX5upMWdUrkCYsbU2/VjAeqmxev6rB
2UfKe+gACv2QIuO8ZRLctm27oOvz5axvQV5LT4hRb0cHDInU+A6qIHvC91c3F1cp28MjunW/jiIq
j6GMxeeOQgFhAAwKC1jy8ndZ0Udch1TmWfcIzzTvomDUk3Dy0CINk2GngTy+aZBEQFFp3TUMryo/
Z1hyN2ikj/behOuSdJL124CBhsEIB7B9dBne1IMD05Ox8Np/sMhL03I2dHCE3mQVm6LMyQ4U4/WX
1D2dtctMISxs817ePGJZ/Dy/O6iR0Gln1rr3Uh642iWyWoYYErzxtzgqDQBHwjJ4N8acNgZiQgSp
IUyv+//1gKsPBR4336GpLeZcK9WEHv/N7ZVHUEHfTnLbwE5dGaa7D+mSiCK/IB1l1lxeXSewD3p0
DBl7saYjVSeZrIb4ze4NJ3JAkyfP7RYdcHtF1x0/lsxdZJSH1x4E64YgSPmmvkEUVIcRNctpv6fO
9NO3uZcUj9feUB4FuP1mkLfXbvVWEtq36M7N4QzMYhj756NXrg6vMs6fFNhyo+q/Pq91Rs6ateZi
YKRQjTnnFp5CKlJk9kOeCOaaIJ/Q8SRpzJRECNNzRrq9A310bxydP5Zbo8FivSlvbKwfaf7YEYcH
tRydqLpMxrbOmOBs9N1TLYhkvcEibhQ56J8jELUeFtn+15q+LghM+5F2v07UtX/w6C+vT2nlYcWt
ejVebYW6O7cgOQNZfbeV3xYn6BCReFr5fSYvhwDVba7v1lF8hpqoJCDEE+3GPK3nLBmE74m1IfEv
XWxxdDlah1MdJWGzLuKtfe94U5gg0ehoIyeJQPKkAoauH7rPFgKLHl/Rdk56iGvwyTHjHUpyNv4U
hAkwSypuwrel8zk4CY2gStVXwsBlO/TnVwdGJzzvCUSGcp4UMjuvs61hgaQvIVfLKx1zzCc4Wcp6
tES/MR9LISngKTDQLF2E8T2oUsYvREzwF7vxWlxZ+xeD9enJbtY5abzaltb3fxPAguxJUff9fcBX
7H0fgC0HxNwOwT9vVbezn+R2GLLB5LV3np+3WJ9rLZQandKXMfvPJNXo2vXz7fG+/LC1CaQhx0zj
2dNQTNBevSxmIOP2xIIAt3i29V7mhwftDRRbRjTgCeu70DDQqFZv+dW42Z5SZRs1qYbFiwVSBWoc
KXip7Kui+F7zyKizDWEmzg+euxnOPzKKcVFJ5HZ46er3B0zzL+KZGnl5erYNtBb1htQT01bHMJSb
MtwRSJsXTFhfnqUHU3Uc+r3uPD3oZyt4JuY9oemXQ/IIVXJzcuMsx3sCIT35nA+2pN/QpYIABi/Q
WfslzAYhyaPHxDI7JGcreJLa9kEWPNImzwJV5U6QZkDG0nyzGeZ65rJqdMY31ExmGKaxFKZh5DnY
czVinFlqNfLpWp455PSXYGqQ8khRVOj1NbrBjnJxLw1oUGSUguosABeH/WrxdBtiarPz15YHvcFd
nEmP73ZYXxetXzhU5jPXn4l5OUhYpEFXUE8CHjHcUROSpet+bfRUxeJH0r1ZfBOY2DNGei26Ns4q
EV95SpQ4dHTNlgzgLxyNFOPZ0nazBZYRvEi8T1S+QrOI/2ubgbHX2E2C2bNaCvzQ6TvzUVlW2Fri
vcoJfKJJTWZkfewz5wUKTLwv7zlMEqD5QR2CGTgOgwhGd3ANJ4g//aqqQbkeE6UvNkeIdytU4/Ww
bKbLOpoLbozNRFMYwHeP4oW/n1XriU1JcPuSvixxMq6XYeA50qs7BKELfvLwhJpiIl7wgr+ktZlf
Ej4F8hhaUM7r7FM8ugxwrWmOOs8qGd7dJkoMPpn4dtIwTgMP7lVn/yWPkh5rwX/CzG0GnUpT94VY
zPvUHepGHbTiovJ75XkClbhnD6tNSpbUloTsVMdovY0V9OPGz+R5dPgrQCoDto3z/snWJZEP0WvL
bqNsgyMumRgyWsNDSaWz/XyJeZorZxBC+2eL0JtSaZoJCQccFJEm8tk2ADuGG5iB6NcPKI5/UHH6
PrTugTYRkJ3fNCU6BgVGFYGEllglpsUzhdylnoF/P7U6glG6lsBryUmTIstjsnvS5qvjIkH+vIpn
5Timhvojywo8ngq3gqLrP5AVnr0Y5jU6Q+DBUfdq5Ga8ahLKeTwCIvtNW/HYXG92MTl2jFFkOoya
cP2w1/vdBuphQaE/xcyNsM6WH4Cf+YPY/7/pnr5WoIXHG9DtxIXmZfXucKgkQcIrWJfvUyMJ+xN3
Konxujt1zgzLPcwpzn+WaK81wCuxdtyJoinOHIXxXo7jIdcAe2Y9pX8UlX6YFxOduuyjVREjA8o7
WLtfTi25wQWdSepuHusII61zFGAF8fmixRYvUpOPMw5MYrV5nKzbNA/VqFpfurCOuB4UzlHyZbMU
OTdcIs5Alt/0/AL80BecpvAukf4eUBEqMk5KIw2MBdpeaqTitz/PQZEsjUBxkyNBeg92ySxXPBgD
v6gSpxHLN/dYcxjDC8MzQUxLA+Mz9Ot6WNn/kZvyTPyxxSiVzd60/a9UBzI7+HG0QLIusKmgzwq2
q5bZ3pPTFo+FK9hE+fN1fTXB1Nnke+Rq/jHBbsXdjIrv5/dCMToHj6+kP5zk4DkY2M19IpOU7RHV
AatESE2NPwG6LRnhN1D6DGItx29NIEef5XcfHoM9tTr50fp9I7YWAHhMhRVzF3jXoOA2FSxQfkaV
rjGNj2FiKOvGip0vJ8EQrKt6OAByaNqFHirv5xM0AK0qzWD+DZx+qaB17jVYM0R7dJhO98bcpZRd
z5pk/C00WvLJ/qWMzMDqdmRHqGzfA95JI5YhgiliQCdtt2nvED4szz9Ktfwx88YT/fqd/LH5FiFF
OsIu+X41CK7PMijVlCzTmPitPAXR8apuhHu3UTazV5p2rQp15HJerOAz+BG5TDQyAERSDHqs7YJq
OZpcmvmQV0FUpsCOluDKouP68vW3mq2YXP9iV/onRek8SiaSO8zQEbQiUWrDWEyxLtbUwtWyvZ8T
hGo+1Xznw45HdKb9JxotRzaUPeQMozQwzdlGVVZ/3aXccQOrAhRFMIza9TqjUKA2TYiUgGWOK6XO
KO2mj3XNj6eWj0z+QYqcrzRi6UcOkg1Yx712+89KdWvQJaXxhIau3Mb2nsln4btRTd+71kiiFuCI
Ls6TDRwCRnraxjwTArVccTDeKrm7fx2FHLLZxW6D89z0aeU9FAqu4F43af/xFFaLJQSryHeB6+wZ
Gos9XpxIdB7+ovibEZwiLIxmwqAw1C+rEgKYFxwfDBY1ckrJg0k7IGUmMyf+UH4DxnwXDEcLlVp+
UGrLGpC5mA26BuGc0E42n3UyToxwIT8hTjowy/V83KfjCpLUtLZ+aX2L1QYq8Rqs8GhpUQ8VC9en
KPJV4lRKkSAEjrWzspGEde6FLWGiLr1G69fJLA7np8E1+T4rkhrkKqGIxXPBZTPpI2Ep64S00TBf
554gJAMTzgzcbJhzx9HLYxcFgF9cggnerHB5qQZ8VeOrMneRZqgJATBBNnUFlHO7JxyuUJcOFwID
9OHEEhd5vahk5wHUv9aipRQ51R9VSqVHpX1DoHX6fu0R4R5rNXYHrOmbhyhtr2l/AzDDBpwadvDN
zXdodF/RWUA0jp3eAcnVeAA4TLBZULbsmHaEmEDGTIaKfVWW/CLVIVxO96g3IAJqKb9YNwLt7CTW
QmOcyA2P1sQlcx0NkqW2L2nYh2zmjqAEnDICyFyz/b2qosGBqNuBol8vKARFF9iWHIC+NTdWF8Z1
p6cgpgSo1pA7+TKdbbctXRg+vY3WZzaZcKm3eSqOPvTItvJL2OuSKBKz5fwxakJQ4ovb8+8NXZuE
PC1Mw50y32jPSVB9d83pDo6+69NLiC5vDHu0hXbNEt5knLErjyJ0LuMHSL79wSaABnO+jhLOgcTz
LnqaqW3kozQ8MkOpN8Zi1/AapGXZkwejrQYyIR3MqsOzAhyEUMyN2bVwmPGSfQfAJPdcByGpxN51
ctRiKy14wf9YjLYETzu7tP+cifB1pGm+7tMKz82gb0xStXaZtKm1BcThWCG0edUj/pfS103bGzVu
kbggFZRZe7u2QY8ZXf9SWpfNJhazrHKwFEQXfRD9zSaMAXpRbj5J8PYZFNoMW7xrfMwwzEBSnsbU
YIpjRhYI7T2Zwo4GvDrQyYR/HS42sGVmNrlR3IKQMLRX/W6Z634c1Djk4gA2S+k6OYmy7BZHYTjv
VrGUAPPEdJAWFAmGLtRhHRr9osCGK8qQId8wRKQrv1c3L1ADY+c2YmyWvXjpH3c8VtaaUuaMB9Fk
ZiW7z3WSr7wOwuyA6r1klTikN4vZXxBgRKia5otptDXLRatX8m1BiEF2kEhPNpMb811nBQFh1ler
00r8PFdlNkuwIp/R0rfK87HlSB6XNhO3htLwTD/tRjirk3DRo8U6+Vg3CnzAfQbIlar8+wX1b0Nl
R5YtpMB7jpzj2eaXSK+hvElpONbJjSSE2hqt/xhGDYeAxJaRokG/vG+Wb/tucDB3bo58EIz7HS+O
/TUdxhgbFrsAgMaRePL67Z6DnjF6dreJ+ydFYUasnVFKCqu/EQbcoVjS5196oW+07GURM0qIAk0D
8CtndFqRCworEqJIdoHC45HjAG9L565uE+3KZNzHh0iiYdD9ATeUeQ3f1010H8/xNcvrP6A1gPBM
WzjkZQAJq5h7Pa5T4KugDoF4neeSGuHovy7FzqJJrDkAgqeiN8eq3FJNvGhL1btKMwO8xlTiA9PR
vWg8EoK0ut3EDMHjPLZzp0fJh1lBhJpMCRfn/XL220eGhTYV4komQG9Bv76X+mfYwnT6I0ZjThFU
a0CMNqEjgf9zQ8Ep0gVJQSImgoQh5PukQHjD5KZXYIydA60gkghDTWCajtyh9QLTuqmavu5Jilf3
5RxYepGdq5E6wZW0r52dQTzNO5x/SjIrPx+Pee+fpuJlU3xus764uwaRNGJpzSFS2qCNbrTqnc1o
8Ri/ipApntnWrr01L6IKIxooNfz8WlzJbnTEe0eU2q9ASiq4BEeSYKELc/4GYv/8yV3atisOKNuC
ARN7/WvvnDTuF+wNue9Wk9uH6ZMzDokMkBzQfxVsXRrMLAAjf2C2w9Ls5VufZWq6128sBm21cvL+
PW5P2TneKsIRj3JRVaBuSjfPrpmy4fZG+H4jxYh8dWfCb5L22X0tWwId4SGN/W49Fv9OHhdF7oj5
3Ssh1j/Fh022/sT0ZNgriKzzg58vHQacDHuTRk/bz6yzI6r4T5efj97fODYeB21jFIIgELj/UUU7
jaZOZPTc79PMj4pUHoc3XrInPjNqusFjrzsDUapHy61qNGPlv5XdZAmpiVSpAyMHQLX/m5mTStVM
hk4I8o6AH1Dd3crIht1aMFmogk1uJMWDjhMXiQRHLG1UMkGWz1CXogh9RWxd9UX7k9Y1IrnRmVKL
F9QiX393LMjrX9JnOuPooDe/9Qc+AIabiVjcWsyBeChqRUw+DJ6ozi6SXpJ9QgTC5WMLih0z/DPO
lWmwHEGviVKVWYql8nIVIHQud00l7EIS7j2DPItM92ywriXZNXKMXJSdUZTXvo2kJUa6ort4qbvO
/wfkjq+nHiDKnUBI2k6NZ1nBQDaYsa3oj+ylqtvtaza76wrRUfhhqDgm1EOPQ7DkHj6Vy1QSZUUh
RcMi5B8bhHee+o2fi64mx9r1rYGS/wBJoo3D/gG1qJIF6MGgkBLjz2R2ziR9/wwIuewIKEHrgvpL
Jmpt6/VzvFZRbyspj+0gx5gsZNqj8W6ksqWF8kOZElGLJELEEY1Yn/G5usmynarhe6HMmzdrHuyJ
GbroyKzHM6WKxvrsvQUFgw7vBTbrHK58ZeXg27OqV9NBmbwsI6fAOr06xP4nObnurb6K0nq6unGn
L7Qvg+1npzqUkg2TL90CVdipAl3nqX+weyZpIju0I6Lv7MqPskO7DFWsvYScJcb622tGfhRXqnBq
+k2ErqlQI8TF73eh9wfeIrNuvOyPEp67T35kAitBbulq3LeUR/6VUepQi03IhlB3Q7X0A2zmn6hB
j5wXMMkisN0o+UBe5YLlQn8F0XxCGcQhqSJnHsnPSNUWKPYi3bCijxbW3GoA7avgcxZonIaZoS/l
7kGE1NmF6Gtfh30LibaPrmXRowGHFGJ8ejCD1uNqdlt1JIr+J/YDK+kfpJSyL1F1Gjgur8T6EQ00
9ZoLBgq4j3nRZx9HuJbDiCYIdZxPNze6BGh2oFBVQrkPO6PGfI008CUMFLoKL4tuDERkIgTzONPX
7fcxRcHhPCiPHMN88CoPiruoxcz4ltrVearvH0hAHWrurU9+T7ul8j7QzJ8V4Z9bcLS68z0maNuA
/AeyzgQnJalQEnebtQBczCPZoVNOH281Es8zp/K+f6WbRISFh0uA4fA/VpKqdxumffLKNk9JVhT5
Jf9JvDBs6+DX7pNu+W4F0ZX0UvvY7k2ZmCq7LqbsLAKzpbrOxH/KZ5bn8D75Rg63QJZyg7ZcWGvx
hIdeDlxIqIspc521T+PsADk+P8xDVvk8zfHeAzkxdQuwDiskgp+MQNdIhK/M/cXGzLOy1YInVHY4
MtngRGeUKU06Mzp3BrKEezX501mycQ0maggmjcCf8MFXuB5dUHSV3b0ei+FldurJkuFEzyul4yhT
LDtlsgKDl/T0EZjcP66HOxfee+kaTmF7FJjDj91Jl8Ei59QHDEiYGh3h8BwEJI936oQSLnOQuaN1
c5E6Sbkv9OIyBC1fcbwTjPP7n7wyfEOFuAw7Qfs2R2vBLNnoNa4xV3QYGZycNoLbwyiORY6H7+6k
jqtma5f/JCq46oah989VWjJ4y0kpbYB6Uwg2sMusWTHmdEgchYL5mWSDXl8MLQrt6LKvKDP4uOY/
4DmRBH0o4TmZ2b7GafCtFrFJI6sbzdGpamWqDj9YWUaRzuVvQYGMEDlQ+2TzGKg+9SiiSbYxWH20
3jyvwngRm1eqNFNPJp5uKFewbXwqU5ngYAdQ09NVgzZjsLWdBu6BV6feIu/nYGG8xftAD3JnbZJG
3pl8stCpl0nGPBvrUbBqLJQpyvNU45Q6HPdHksuVVsMTucy7uMLxBzhRgUyUAnHkB6HMYH+E6OP8
QlLTXL+khi1iMi7H3pFDUNtjEnjzIN0M7TexDUe1Kl4Nl3eDaY7fJBx1hwZM8ic08SSn+H69RC2/
hTl7ElrztRwAdqUiYsc65aGyaUIft132u+Tdu9ugh3KX0OKn1eOf8abvm2K1uFQuqX7XnEfwGq4w
yWPg5DgyqxgXj+uyaUbReJtCrRI51vp4c10mZuFSidHLgSZGIAtgQGTn/YErePGsRO+RrDo4Nycq
ziwwXnG/Z9BjClbvo23fq9K01l1ypXfExLZhlA4QcXUs6iYWt0xkdbr/Bo4Xh+aHAMGKwlT1Y9cb
gxcpnVLDn5RSFgQNw6nmrq5QHBW0HGtl4JDOwtSo121o5IUyv7YKO7loLS+uVE6LD9domIK3Sm8w
DAtDIMrx3betxnWQXPIFirZzEPzZPFEfMuVgqI8z6cAYlX3eThBfifZvWzdHlJEPt3Vkz2fTuAzb
+GgMZQsE1wb2hye8zG65CWdUg1a2tpvjZkmdozGyI7B5Bs1UpOxjy2BJzelamh2FHARqgkCaoI1a
Z49L8+o4WtrHYvwE6xMhzmNM40C6jePlDYg9x0aSkzDCpFW4JtGa8CakpcYvUp9kl5HSO/mMX/mW
L91Ui8D5/40E9hS3ZeN80KSixD8L1tMqF+RZ4TG4g69rKL0H4W8LVCEmLGnmgKLJPG+t58PnEmsR
KSeXapK6jUd5R7otms2tNXsmIDEtMCEIPq79bRDUJTQTUMS21ztp0FNC6wWtZs31OXVtjZRnBDYT
JueDYfsMLf2H6y1lcY2j4cE4NGAcs6hIcfvQeHUfM6s2vi23U8Q+pVBqP3z+4DodamlsNsrIxR/W
d3Epp9Qbcm7njyQlL0KJcnC+53wfvV1NNHykpmuLOuYSmbXCMAAEVEW/j5wYroUQLDowPzLLerjN
bIv5cIEANqpc3CUmFOuCbjF5zS+6YzTyrw1BN6TX3qHp+obYMVm5mVapndoLNeKqEQ6GqnU/rm2K
qtrwi1m+9avMNkQNnNRrwLK3iP0U17dWuf+wVz/g6WXdSP2c7hswRwsSObFLJSt+gAY7WV6yw00N
VWJnLWNQ2uIQZXX20XmiH5mxFvDEnpn6/HWKMrkGWd3AgyBjUz4KYsuehE4+lot7P11lRm/22pd8
ZKMPqT/d7kLb709HTmJIKUVOHBqQnVEnKBEdVQD+NC/GxHqveNFagVVqNFv9uoRlWoRoNzI5rLCT
woB/OYNYpdIFWsQ1eNk+4FB1qYeOIMiUgZb4KGP52Bme/Ts0H1CQvTbjlF+kWii5luLiIkuJsnh2
8JxZNtdn3yCXWx2+0fjDAtRklVXKACZ40/57VEDapIUdVOSrEViy6PQWL8mPfMciBtTftWh5KXRV
u0jNe0H1dpXb7mj5OBBIKAPKn4cQZkTzBs5HbfOjSxMMqENljQ+fgLZs7r1EOKQb7PzwznQpERZf
qlSTjDcpKhmtISgf7tsLhEq1DWv9/Fkd1ahcEhPc0YRQxf5TJP7anlhRGoOkamog2pt+UETM0j6/
h9EZGxs89Dlzc3ee+29/2h1NaS93UkEJQFYrKqM9mAxS1ujt1C/YK9kItJ5OXsoJdWJFygISFklk
8BVpIsAkGx2StRYRUo+eN6Xv2UrM/5Ja5dmvZxy6qORH3Be3+AmcITYYuGMUlilzFBq+zloDuheT
4iZWSy/2UojS3/mQFpBmSRBsYQ1xz5ILaQ9Xbm7DpLNFpa9SqceW/vMdOLsLdcQMLkHcXzUHjd6z
XS4IMwM8s6ULWrNTGEhZKPWn8Pb0SaQem8ULpMTQ/EXHr56lQfYiUIl8PuWRebxM3G72NFvIDXJV
eLt+nz+UJrPNlsGBIRwzZ3PqLaZP2WJqoUL2UvGscNmSdlpG6nZmvQftiH4O2XN2vHG/xZeYM7jU
7RP6KGQ7jWiXEZxKFaJtjo8hGUvk9m/+PUSodKC/jUrvjxxkD1GXn6YBH6L6OxuwIB1hi/nlz9B5
YdfumRs1YRh40RQR8WysN1EpiT5hgddunb0uupQbGUWvmxRm4611bcEiTp4NGpj5uPx8RChdXov4
IxNV5AT55Z23eJIvJk5M7/7RvIAbOp4JtVcPBlXlGFXe2G5C43y9j1TYxhMjSiIFFq72gWoJo4Ua
gVzZqlDejGAmX5A2WJpWN+9+r9sPSuZ35U44lmA9Xcl9bk+Pe+kmKTBIFcYHNyocId5xngFByM2p
kTdRKVyMPtRMvNPehHfdaiHHHZ0EiGytnyc+XUQhAvN4jmptdELnGswbYqGZYBXApr13UMdmxvbq
jVeH1PndAI36ENaXn0cnbE4ntziP+mxDBK1MS0roFzTIFRjT3YrX/ifzsyRAhugNvRqGBNnLsNJS
FKJlhNfXwjvY8pV+Rqq8GAK/Xm0oZzk61p0v/QOGxRahqhsM2/XuLWNBDOvv1vNRu3yObb+JKBt0
4wM7/fK+mL3aOc9haUr3fTa8PLLsL5iZxehs43YXp7oI9OQG1nhCgC4h2kCjJRZgwJCyb6Kf5KJo
YoqCLNYZvBzurdivfdNMt9L+zFoiSz0+qly+QRzs8l95WB/6h2TH+OdUhGt5kpJbASIs9+yqeY8q
xbFnToPU4GtuF3GllTqpwUCXny1cB3yd7qga36osqFzB0GvTtyMS2ZbYlFJ2mBZKrvNSNhmo6Pl0
AM78uwoB03hp88A00C/3IXpm6nfhpcQz+gv/laPKAhDoW99ecBgZT4CFbd/JoDNDqDzBGUmBRWdI
4ERKubTA2JYp5NLxOa0sM73BPN6kgKEIGnNjM0Dzm+2aH/PL0tcknUiPAigVK+RqeIa7ahmTpnqD
yIPOoP6rjzvmHr1XD35WxlTZmPDHRuWACfdyPQ+ZaBBvKzGZczZxvuMWuJ2CveNWs99svGBe3t7X
WBwl+nh1Oq5cUvL2qeW5i0XNWz3kKVGPnQZ+11egdLljr7PgsHQGTMFx0WqiI/nLcJZwWWToFY6+
lH25QO5I5S5dHGDleLwYJ7RPLeZgb1a/BYDnezIoYCV40IGx/4iYsrcE0NnONjxQNy3JFL/fXdcs
lXXI4ltKmx6zIHuuDWlUa7avDE+tdELIOIjqnRpHiM8iEQSdkUp1JcR9B6QvocK4skK/ppsCkVlN
Sq7C60vpVnG9wlsSEZFdnBsZBpQIsiZvWup2RNyzc9r9ewk4v3luou/fQZV2zKhlMi8uBunJzqYS
cx71PWB35oUI9AyEgKDJsxJIElegfREGf0uHOvxW07opCAwKXsSbe6dJngnrr+EsciNf9HxP8+dv
Z5T4qPOOfrzqV4GlmB/FcGoeXK5SZVH3AfYdRELcyTj30BrG8asprSHNNshbM+cXU7BIWoCHZtCs
MNSJ13xKrytc8GSLhXEq1f2t6WInfkEVbdkyOfuy9EsIBeXRWSOQNHAaI9so/RwoR2xDAwhJ340F
j4HoJYHOkJo6MNz6lIyDz4W+86NPPRJJX3PaP/pR0oBlU122L7GZqPFR8epwrbAdM5ozsgMiDUgu
cl8lbImEsjptRi+nKn+EI0fGnWaGqwLS9v4bd+3SZm0/35Ij4LrHIMplHKca8NfeKo3LLr9pH68U
W3wU94DU/8f3lFFZsGkPsVyOUx2bZbIKWQbNhfM9p88DKZc8aLz/2cD5VS6ozHK5GTWk8cicQTiz
WFPpp49Q9+djloj4emld1HlZqkPrIUXw8uDzsWmDw9kYgJTmMTfML3iz4B4bB6pMvX6hPPPjhK87
OS75LUo44qO8EeNXXJWF/62pXUDdqLS8/a/ahOWEzkQ5ZFyjevTcIeRlnYvPBSaZr2dKOiSw72Hc
bbuBNEvwWweMZZvOV6M2EK4bQozK/vlbGdt3B13aBaifa4Lo1NjkCKEfataaPe/RtbvPipf101ZJ
6gGTlIeneFHIQ+fphyZPrSenpEXoA4/x0EDolbXgI3Fvagme0uzxpyT/4k1aE2V8PxNv3onmMXvk
/boRsKuJxp0rRd6GQ/7v6fA3KShgA/dkdBJY6uhCcrY1NS8auG+gvfVdYrbirZOqKl6ZwSjnYo9O
1g8Qbfhmfj0HxChPmVrPcdyS6zVvHtyCPjVoH+QCoLCK6MddhD7zzLWmUG0YpWYkPLGtn9N4w/BR
niYJ6/73giDue+O8VoJZ6UsZjk3S/h5BhdwhjTz28kVUHEZ3fRe6BS4VN1pmwpXPrd4/MiFjh3Hh
Bdvptobf5zJ4bVRwyRUXo2PaRGHmZy9M6JMy6BQCjpd+JAh/qvLTn7HIcW3DP0cERmteEpj2foqm
ZAhlIVfJ9EzcixJ/8i8S7Fo0/zZZH4BlNB+z46plxh5BSFXCyj4csguDG9p2KPkOSHMmgSwrDRpj
E8mzGnle6v5Fxu7fN8tnJElUAw9LYq84ara6kvSZL6xMfHwralBEyC9HJlaGBJ24I/H1U57zVRvz
Y/lHj19mZyXwHb0NOHfVl9sjIawqW5uhkYuDrnneIvI4Z7V5Bm5WV72XxUnAKUsnBnMyxlVUu1Nk
yH2P6M0VH16mliLUHD9dBYwo2trISOiEhc4vK8xpA5nlhQ54bxflLsY6U3cGcYQFbcZxm/sKaMwe
pz3gX1G8LtBoGoAI5/9+wkHRCaszcMJmeGfNfjO5Rh37YDaSUahTw8HyFuTKJyiXgCDIaD+Svlme
Kqi+TvOwWwFImTL4nkY07dE4Oj1lKEJOWpSKsujjLZVVhSL9p1vp3O0urbsngxbBA5rDe3eK7vOD
S1hlRlXj2u+6cvAJTNakQGbq1Oi4ZM4n3rci2MfhYLRwPqWjac97FcYS2vnspcZreSUlhgAANfe2
jNzl9nuExq2ANkO9d0YHZtpVgsmnboNoAmOAGycgLYQnhfEWayZ++TpYH+di0CIr4tp1AAUIVcQ3
xjRLM2/TKN0zgBdigIPTNrDxgr+SThokO12ZZVlXWnWwAO53inoUd3U7cDrD2U02BSaVoyJsX4Py
F78EDury2ZmdRmhBebwWZmd3AbG0Apr4P1aeYrNqelaYDPhLV7WnBR193M/rAbJ9u/AVz27Bqe5/
NoXNVNSyJFeXX2mby4KZTDvnGFyd8fkC/CGwu7H6h1+E3Za6wAK7pbe+qzZgxOL79V3fZudrzgpH
/9KxKYftw0iJdAdz66KfkJaEB0SbVHbsJ59OdVX8ju021aVkuwi1dXJVror0EV5UDY0rAyfVQ1vk
FGZhCvZBDjxO/72wK3fpqftHM7/8idnwrc0aVOYZmQUgugt7zX0zN6P26PlAzxoOFceWbhwqfZPW
e9ge2U+NbwB9nZKCAc0w4Mh+YpTfpjH2JMlDCCVT2gt7VpEMUs0CCBSRvB32WuFO21+KHCSMxY3+
wy/hU23EKSUdlk+9/laSHwkg1Fs27cU+Zk6479W7ax7X8uPDTUEzyTDT02469bOxCyL5CH/ca6JP
D+/jH/IzxBVtomNbATEEpO9O1g3k4euSnhz8Bb6G4LC+pQ+WRF1XpAPVfjla1jvMdKqZnSNuXNem
YOOhgWomv1plnX13DunnB6uNObsC6xudc+6kBK3ZPjp9mDEm5yLXXl3Fqp7zMgQYq6SnVvi7DwD/
pjUNW6LhIvT44e5zTxeoY84zzGy7CxHOmWgO3bABkyf9R9+G87ZnvByBiMS6TaYW56bKiv9Juz08
HwcUZcwO8mqLqiSacF7V94iEFxIGV6NNZVNSdM+mcfrzDZ2dl2M2VYBcQGhMf0abu59mUlWBIHGY
lvTT4Hazk6FrD51BFRD/WcbzQ56ZpPqriifACkkH42UpuIJzs/0yHNg3HcGZAJmDQIq+cMbXcWna
g/xLn6VAErygTgOePxDXR9KVe/5/+4cmzfeBRoKR6rhQgtDln7J6utdlj7UmeNmvLCFB0NLdYpdd
DTIiguDfMtVJC/yo1qg+agfUvLIvCm81hipzPaxb0GsrxRFMCR4L/tAnJ5ZvZqduUpjISEEMqASd
SG6ymisAvXDVAGehKrvcwBsn6NCD9nrKZVyM7YtM9Gn9MvblVtckE1AUb1i5L+aKIuOK1lCSR6V/
FjPWOKRRiZxiK8RAqAHg1cGSKDH3Pgv3/OwKGgAVbf1xo0jifmzuW8uq3kQfQAyZ/4knycU1wbrG
TF3pLp6nIdIj3iMFlPv5Da/VIgB5t6beXOstTsVgBtEWaXMN4w1xpnHV89Bvl7QQgGm489gsxwZV
JlIZZP1cWtWM7tti+mTsgcq/qACTk50FnFbQnqGE5Bia8/GHPX9kKV/tjDQKDLkG70UWE7qFJWAb
cKl910BkxDLN/oMTksanXAvcQRGlVT34QdNnIm+rb3juezyNKq3XJyxZdOjtGF+2Wfr4LrK3u3us
fGt9xCdVYXqLstC2I/aeiNsscih0LNzt6mdCl+j7DMppEIb81zQEZ+7yRChLFKqHFh36798IdsLf
49KRDgTTqKXxoJtXolpxkC9hNbPLy7uGAV9vLn1P/9+PY4iTcKef6m09T+GYLXukWFps+602W8Iu
4Z4hJcSv/uttAuS5K6jv17kEfs11xT6Tk20Oa44hPKBs0d0GsTl6iokUSJwdFXwMuUroMNrgCiwp
VYz2lu6bFmZboWLDKSeb3P5gGUOJCuwFeZIu/+Luip8/2Po7ip2LhQ0fw5+xILSAIHL5eDn3gN5n
y0I4vcykAd+oYvJ2tXfLBLW9Yr1QTmc8caC8XNm2MMixz6wRgolNjK1IJ+SJRDz4zpvt78xUB0wI
lboZqXizaOQI3mvqSS4tjmoFb9vHOq1Bt2LYNi9jPGJpP4FeIDqi6DDisvqAw+HfEH7qSbvGjKEa
DoLKNKBZBcMOSVCJDJ5VpMKs0y4hWIgD9boYOcvTtA40KcEdZuavljVyNg46VkWCaGVbh1zUWo1z
dx3Y5mVpLlth+s3J+p3wkbgBDfjymBB8X4YOB7BEXUczGAc9HeaDxN8zsb5hihZhiUi8zEhP58LP
7GVlKKxuPFqq/HNq4xdbAg/WkJ+3jxsZalLizFQ5JIg9Fj4S/BYmGUx/5SnQLKptjOcrAhZxWlwp
i6VP8hYWFURze90aslsQAk507OqQpUkISTQkk6B09sEJY9lVePTcy/v1navhXwLCvPzDQDXBaOom
jeuSDoI5+CwtvBNFtyPBeSylzYcFPr0aUivsa2PSLsXAKMdvBJhHNKjgA0HMtibSB8EL3/8CYfZt
pT202lv/4gmWQiq/y1OUuUhQPG3k5PQaP0AQtBSmGkaXpiWH5uIafvwrcCbB2SJm0lD1TxzFcs6s
2t/nKuzhF1RuT9lKS1VVVcBeX+N+JtxP01wk6VTt3duzWcoDszhnBk8s0AWSpNLS0j/FTfr7dJkc
GUiT6QgSvOJVyQLiEqVrCwzDKuZAAKrHLpjMMDdEN47snawl/UFDeIimH8mIh47Cpp7bOsYKuScE
YNuZYkGS5dCJYFPjGr3E+yi05YhCvsmjGBFqjuwhIH4BA/wVUiS0Yy8Sj8HJvdzZHJy9jUci99Vv
8y95JUDECNs5bageL3Y/mM5W9/UQ2iCilGLcPQ2idxaAZuBr0qCy5WofR/ipR/Qym9ep5lND9zRu
fiR2q5iylVK8NpSsrcCJDGuV3lWwE44yTiCWVSwRuB3MSC3/SwDeveZyZBaqaiDt/vmtPlb0ZbAM
itxp4MMj1hKAa0eF08tPULlgj8Y4llWOkFrM9/QUq8/EU/yEqQFDpsdBrIqkzBTNJF0vahnCkdDV
QeCsIEGzgSXipxZ8mEngb6epd/FueZxeAtLtJjgC+3muOwYL1OBjri0XAUpeeRef6s7h6Z2aVLNc
2oqVYUub/ZmVd9XliB9qByaZIpkUKzUsEVnYS1vBMn2lwpcOD1F7ptUEbG9QpApe861CpFQijCbL
8w3BiK5uLGUrTs8+UXQFZcM3QeQSaaOfA+o/oxs9cWe38g8Bf49QbepV5D0VuF/Yprv6MhnFE01/
5cbjWO4GaDPzDGqz0pAkrEjgs9WVOGUh2G8J8kDHlurStZmR2qp26jD0BOl+ZoJRZWD/nvC/HJhB
KHx7Rli6OZe2RsKQAzUoYO1gtFrr5XOJyCaXgoBvyhJBD4tFzX1HzjH7eTGb+FlNzgqXKORdVP6l
FvQerUA3+52VD1YvqUZS3j0tchn05x80ceVwGSZOow1yps1f+SvAvwdEYpoa+vLcDc4S082tbkHd
WGdHg0myFuIoZIW7R+L6qfYHVP65ncLXRwfaDNwiLbPFA0c+oZHFMuML5n6QPr2a5x9iv/dILhOw
etcSidjtIOIvBE9D8gQISHBven54+h8DBKTqWsrAu9/bobyiGfL1cejuArLrEyTRsjOCRlEzflvz
kWsHlC5o0jbeSY69iKdYlz8In2+4RbE1/ZL/pNgfAodpqOfCsu4CQcGksoGE/NwyqMJ5eeJZH4+w
GjvJdS8lO7b9uCN8rFvSGX/9BvmbcFtvPu7Mp4ti1+fERCezGEHtk+kCSCEY7k0rP+AMao60sBws
FHsh3JwhwhQ+3pT7uBXMpKo1vsnt1Hvp3zZP8HKl9mAKxh/+Oit9b8xzT104I+DfGjaiKSQhMvYM
WeVtZgjq8EU4ofTdVKGLNljBMfJEhkhBK+O790RTDHSgWn2Z9bC+jJAgnw/pz4ZIl+dr1sn/BXkT
xutmcBtkCEbp8FhWhGA/AgUFxWW5V1Q2nDJFwUxRKQo/FGj3j9mBr/kteNGbmjQhDXFgv9Pfo3aX
pZXNc0LJvabEmsQYrSLCWEx+qFOin8Y3dbqeBCpu81lP8XlDZ6NFrDjumn5Pv54UPdq1JOlekUwr
Z6r+RXIvzYCF/KPl3dhmItpGCcwSYz2FW6T3eX35XXfGhqdhkFvlIn87TuwwWVng2cU/2u9ajnPo
2atw5YrK+dMWod11GyPJNpZwUqTAm1Cqg3o8xgXJXR3aCC62PkjdQ9MhI4cdH2KLiZlG+LUsQckl
UGQL+WEqzxYWC+tMHCJjZ20kmozuW4OOz9v9u7CB09sDjVKTbbQ2TdzQOkH29GSntBpwo7SAHjYY
6CejqcRJOEDhH1CAieqp0/nHZ4iOkv1dF7K0874ROBeLCuy7VF5Ys+elZEx9tjh9nDF2y556mhvM
P1KIZ5sf5kfXh3qzUdO9Iu2ijNmCvjmargtvrOst3o1hR/XY/8zSGAF8mdlDxyMSR/+Klr16MeHh
A0RkDAVGOE2f9vYRaXXRSvv9Yt68f4wAm2bcGNd2FE5LNYw0ExUWPa01V63rjNJDKXFVpJjkcxod
nV7wk8x/JtbDbLrduCUEd6zPVBm0DUq58qGv8tFm+Mdqn+b98OuctbeJWT0+MeX6MmnPsMM1UqP6
haRRZLZAbD60u1ZJUw/15bnuwA8xFRPhd0lyf57vRc8+MkNwQGXIYDnvkzSls+KIKTC+VxaTN2xc
2I/RsNfXXmUQqGLEdgyyjUCCigE3DA+A7WH6Lx7SmDKQbMO03IP4gk3LGtG6WLGwlifPw0W1Uzgq
qtX6wXyzPpDqengoehydZQ30ssrLXPLoELRacAKMP1Pnh2tWxW9l7Mvt1s6XBa8+2ASBgWpdUGgD
sxqxrAWf1mZh00T1jNMz3dKGiXITKn9frb7Zh0MoMAeCyjVDF80N1GvobQ2OJjklKEmZ7YA8hrlW
YUTVXVMLFTVILfCXrdL1xGyeFnhuqKHGt7x3gLsuW853vkV7evbwWZir9DmgZkdSKHABCu/6R7Cf
u3BSXmAz3c9tHlhHdSNmA2GrSnbX7m+hZBRoQjegE0RXagq24GETrxZj0kqOnCfohWYPHyPhRs5z
pDZ8aZ1KZbToF+5fFTSu6+fT9CgLxD8fJVK5YpWjq+d47XnyjuTfMSQVSyGKTMdbWGoGWB9E7TRa
DdeD15eG9woatNRK/5i+CIhWVSzPctfscYzABo1oXrNdtSd23JEJ1ImYSuWpVWRNMTiRy7y/qYQK
F6AoNu4VmRCzrWrB8xZzZE0ISa34kSNquKTTiOzFPBdpvP2m3GNL4KqKSrxXKxNGBFFVubkLq3YN
CPwBfX3TwdLOwhXhzwE+xJZDrkl8o8L+pTQ6icHLxvQU0b6hmXAkbkKwDP/D0sxefoPeVs9XsQ4Y
Om0YDdussoQRprpvjjtDwiTSeb2CVoLJLiGJ9yOeDaR8wYp5QPw2tfwPG9CmicsRJhT3F8XxVlQM
JHvBvdOw8FBDeFujJaUkuznOv3xj7bKEG4yrzzt9ooT4cmVtFw2WsR5eeIOpQs4WCKMtIFdLrXV3
wQ+9dwuZXJpmkUzUdRkXWu+7MM9+r/xBoNm1UuqPJe7dXuNtSiDUBV+9N1BDPaS3L2UlevMHxxyC
tWAKTgcUnca5hlt9Gn/wG7lBbSeVtk8fyWRyfWzy1g9axji2EmCxKyZTROe1XBZRpnA5OVILFMhX
+/R9gARgQfIuGom9oahLTA/rK4dmw7GEKFpGG3s1evBD4o6OIRfYohU1HdEJJcevP113Hr+FX5It
Ck3qrmgXjbPiKm350iKLJyIEt3XnmbqIKQKf6uiUZSZw9sWx3F+G93pNvB92kRIrhkwD7bc+C1Wv
wqV8NN/jCAv8C4ZZztypVHqP//eU06TJ+8Bqtp8J4OGoXoqLfhN4o0foLIA8QZHK8G6olzbNfb+Q
1AwVZAWdFpwVKk9ZF9AQm42UtRfTjc3Gd7cwZnJmt1NcLzgi92sNU7gcuDrUNmADtwOgN1suF6D/
yG+KmdeO1voqQszXsVhVBE6QtSBmX8pTiAOzk9rMpwOIFf7WusF1EOVTlOTBm64QkJ64/IUArok5
fl2mhok0vgrMPtThBrU4zD/nwEt0NL9lrJ6wwBds30G41HpxHsvMe4qkIXtO9BhpoNRW88qyD8XP
d7YRoH+riNs+3+ciYPf2+xnbyHc1H7Ufj+yf80WtPbOJsqHAAua2YnFHyZzJak6UWJMgi4nGohna
rVKUj8uLCH07lLwc0YYpPUstpeVWe1gaRexCyzZBPJXhVHdSFhWvDsjZQss/rJnRUTg6a3P4pn9i
mSZUYC0/9e5lFJ5gI4TgSyYrn5Rsu52J+1SH3EtfyfqYogZqFXy/Nv83FFZHf3ImwGJgrmrNzl3U
EgcKVhYrrgu8hZYORNree+LKLiWcJ3ojBFXuAdz37BBd6CnS5lik/8uRINO7EZmym1zg+Kq3e74U
JWhkbfs32O2GefHaUTOAnOD6OWIwxlhNv/qNKaUPSfVOEyQDzXH8CoB/df4fBiEPiSJ/Q5fKfkL0
J/aQogj44UzOpX1VoeyIyk7qMbmtBBk1htnMDNb+Rod4Wmql+7gXV/KsEY3N0TaYj+TT1tW/VUhh
36MKQU5NqTJG7FjJmhdAsgXblvrKkHVm/EB/lRnKrfCC5hcXNAT06KgPG6yHjtau0O+2H6mLWdDZ
ZDgaPpbaoXvsOCtjSOdL/juOr4ztM2a9XNQrOYo/4owMYzl9IJOlpYF4RmFIuFb9awJ4lxgcj4fB
Q+k2PesuQneSekoP9e0plCvibAPyOVQHTUhzeN7DJMTSTl+gdbTQRA0GK+YC7X3YddaQ5Oaqh5Fa
SReVUe6fz5TlH6xr4ry2YQmi+Hf/HqMc0PMvso1rDH76rUHVtNEIOgRZGRlbj4GwOGlmJJcvPc+X
Z3JeG9sF5jcO0OCcKs9sii8uAobR4TwKUsxegdz33FjX3RFTF6qWmbmwLzHXEUhJmQa8B2S8h8Wn
4TG7zbs3KPb81rn48OonYcdDEbx1uBqQxRjHFbqXm2syZtiqaSh9QrgOipOU1h4uDdiFhps21uWE
braKjK9ZhXJN59H7Fegqd6EASJZ52sm+IJTafCrIxr0SDMMVi/XoPK4XNNf6BhssaQoJ9k5H6zjn
B6CgiYaE5wTkk50j++2P6NXXNCTy3Ndc43vizGQNJP8vM43NYn860Y2GCDo1I5c6k+5zcrr5nZUg
e5s7Hmt8N2JVdyfpyzqUjnIvHCpnwTZ1Dn6ZKLVf+16Pu4YjLMVaOaY9t9B2YD9zRCwkpbTvGPK0
2srhdiG7TvOuf4FYAjXKI1tXuCWeoHklNDEL7IxHT3K0J7UzfT7m1vezZD2o4lEWp1qFAFq5oBQN
KM2qWmgtC8RhhrFJXwBnmYDayMSERY46vwrYD4ANdfIyQq2inEx/enHPXGiReyF5EAbpASfN4j9l
zcMpDVF+l++v3USYRN9va8vKzNBqPRlBso9N5h9c1bixVpgD8nKYbdVQYurb/ii5cI2XyM0jbZ7+
dPkST5rJlZaKahMsmuXtfN2nj3oCFU2Ye4Z0+VpXfeZSa7nyXAEkGhJwrthYrNYAfCABEVWErmoq
7EHcOqdZTKM1hRymk9q7W0jlsTj3xa3qxEfRvui4Htq0Kfkn80i+wmI9717pxEZyfCTaQR8hsblP
6TWENHDq5CzKHzxkNgbp5h9bhRr6UtguHo4yfdsQbnircS1I4XjEg7B0Et24FKDs/lGpLVgJWyFH
vzgMyIUglrUDpbQ9ETDbhyFlMJvQdYrUL/oKZhaO4wCgjwxSMAfshW9EhNJ47aUMKarCVRwtx6aX
fI8s/yLe6CMgVXVeizxIOaqfvgPO8QR6bhyZiE7O7xf9fHyUmrxCFVtbMyIJ/93pxd1W1XElvn0u
BzjqfNZfxx1dkTNUebuXctw722d688orhlannVEJhb91gbMF5wFbfLsRHjj7Y0Se5sLwCCnXonQk
RkSsPQXcZVCr98D9XB+NGFpGDQNT23gDxtcmBHGJSP36afL4P1Z9hFYZw7iRF1KJrzXP5NQHJOoS
HtkULrDL/fvCHFi6NgwELnwWPuUxbdZjmuFtvf7YuXlrDdFogpQPvGLnILk0PQdZYWUEGwcOhRcq
tj7d0dvUUNGrhjP+xdF0Dext4HWO17O2hnycdP4q/l7EiLxu2liNSzAIkS/eV/meZPzJEFm+4rBX
7CyD6QAMsFfIbPo2YxvaQQnReIKbiTNRZfyXLtZFpeXogsJVMiJ5JpQo9bHqCbrOP0P7jLKPLeDo
n3ZknJsdnGrrOzumlH3LAq3ysE8ZLlI4hNxomLWaJwE5mXNwqacaLZGNKDw4mxZakMRCUg/Vzdmf
x02pJcfTv0jVB92u1nKnifC8KEpBlP5BEbVySDJBO0Dnj/KKovdjw3ddGCOcIvRjR7j88JeEG9Ve
L3D8V1WWHSDptkcD5iVpKLYNTgC3DSBG2ENlaKJnwRYHE751HZnirUixuJSf5DHLHL6pEw8mM+c2
G6vl0fXN24n5xVSymSMIlhBKd07ry4XiQ+3Ocl84TzbIzgb1YnlrYx4PVnQB3gO2euN176/0Noaa
0wB98lPQWkXJmd8HMV96rImOM8F8WT/zzm32fReBoo0A5KUJT/sHqJv2UU+6AVXXu06m1C7r674q
v0H5exVAfc7WpRzsY7URoyRAYUSY6N3nHSg+6D1cKj0e/zjgIzpJfM+/GutxcsCq+boIaM3Mm2Ar
a+mdDYeP7U4LK+GOqNaUkz/E+QLBnALBct2BoK1Cw57E/QKaUQgWUt5GCsFv/bDhtnRv5/uOYgbf
OCOGRb5SBloAGRGlvFY+B/J33nQCP55ABPjni3p9D1vLWTQH9oNvFk7m6KsjYkxaCF3fhoQCkxDF
h2VmdJbwXvSyr7/7lZKP5nNx0tY6XS87bHxxGSZUD6R0BJ4GBsgO2ExdflGjfJD1YanXw6jvprJq
fSf8TzGYUglkjhPZiWlxLPHAzw4a8uTxflq93AZa80MxcXzv4kRVH8OQbmNU5md0szJlGZnPtkv4
O0ZhcHDRT4Vi/lJCHOp7FOpSh28T8YnntnhGOjgVYNfxlcRPIpoAIlIkv10/VubNXOjGc9GCsrVb
cgZAnUB2AcX2phylMRlmIbTCFcm33ObFSxyY3QDB76tyEw5sKbmiXvPti1UuomDLkJafsHRqqytd
sADrO3Kd/y6Oii3bZHgZFZHNXmsVzTZA85//GaPJM/8RYvxaCO4KEjHHZEeDSPWctpHmAvNtNgWc
fyBYLhQdgnQqWnfuG0tcIBmCn9E5Zj+U3W+Xq/wDNkNwP3MhVjMbgHY0R1/epWDiiWM2ml+xRvSo
zBC0OcW6Bw4Y9ecXr/p5mk/hfrthFz/koOCcC2upIN1vJCGsEVVKWqHj76dZzbud+bH1NDpktvrI
HvD0VGOn6kgP3RzXdlXbRLOSOTFb/fBmUwyfaqjCXp0TxnJXd2m7OzSUqHJmgW4wVdULWYOkZ+MR
kiS+SWKY+aPo5WM4RizOYi9EArZ3mBvp9iXPCQYBZ6Y28T6X6ynlkjaQ/0l1bUP0UO9WUc7O4v/E
gpKFInCcOQJudrbkbsnSqdn5BIb7iKwUjAKyF6zQEZIxdgGhs+CMh4zRN3GU3HRSivckB5NOjRp7
WeOofRDMNKJhSZtGVEZXjWH+Acyf8206gArnJWm4DwzmEzNeXHJUgx9u6I8mz/wXk51snXOukgfr
O9SG2jPBBXCEl3lamngi122ScSTcv0z976NGfHsWnP3CZFTtPXLvdFyBcrNjuDJo7+9MkNDKKq3Z
LGAsWKonv1EG/FWSoChWgjgZbyM+x22b2tUInEJbvDRG8r+x9kmrNfm437krWme0aeKKimfGu0Po
C7mS+yxq5uGxMbolX8AOH50/Xu44+dvxl4I52Sj9EQ0rsE2R/ni2pbii8YF+7cuyxAuYSKjVdlrd
27JmvRgwuPPKttIC8V0hfy8EnfNKhVDMCpQWMFcjaY4pU30fMYT/xUYVg6xngGwgRbTKLiGyXZwF
aVeAvJIJGbQCkbT0WM9E4BHsbGNK6nGsKza09ansSwdPh89tH2RJF+nQdfJlzdtCQUCHu2InW49O
QldHpvIhYIlNcu1GZ6HgLtfadC2xsBroan5rJ7bUPslzD7a+FssmtGQhYcW8HVcdwjHuwuXNIdn1
B02v7B6PqvUNT5Y/k+TpTTcBYK7w8Y5/gfQizJTG6/4EWPQZql2F9ZtnZlD7yU/GLHLT95tqvET/
naGOSX4hs6TMWKknJvqplqj5N1aH5km1ULVXoNVA6h1RiMpEItQau1SuKEVEDgm8e5lvIKaFVqi9
S+l/02W4M4701FZhx2InNkeX4Kjvn4tuLXI57vBdWQ5tOMPadbikjmHS3PFS2g5s0EJz1N+aBWQo
CdXb1K8QSd36npuPg0ks5g19D5b5KqHTEHRGDDklT4hfyzJ8m32SptvVD796kIxrXXvl8KN9m3l1
MQKzKX95Nt7WPwbMZw2h1OFhe+nJKDqNB+9ESmhq6fjx7HiylP8Xyh8lv2LcRqxC8cZoN1UvquRt
9Xb1MqjDUkwiI4JXIgt9RAYvqHREUceI1yutHoUP6ANwWstpawrc72CbuJ7cupIkslDgZ/3S3ayg
FcmYtBfmKGH82p69+pLpmiAkAkVOPa0/PTi/a17B/EVZkJN87UCbSoX7wsnY0vS/mXc9iDaJbsR2
7XizW+52XYaQG2/rOKgItAH4yeljv55juf9QnMXdK2Egh9cg8fwO8p3l9Lad+dBQAYxrnxwJYJGV
HULEXifrxkbEl1PFWfeNmV2OHZ2g/8TmLvZ6cr4MhnQKk9XYFAbhL07mXvnrgiZKUONUGuucb5xd
/paPxvbUXxNs+MGsFNswZwhhwYgXETRute733/11Px93Lktj6UuZXw24dys8xwYdBYUjomQCBS+/
rA1V0WgVvaC1NhCYQyksAflFv11tHb/F4Hm5KOyMn49bU0sDXCVIghlkmBD1UZuZ6WibYOwc5eIl
o4xZqURegAsds1g0ml7TEreoa7+oebdqoyL5CdgysAzW2lK7NK5yoBG0Jnq5osf1KOGzC8NQpra8
Dsh/rzN04U2kt6ms8QIh4c80wnWYDyKKK+VThS+VvEph3Mhv91+fn2gla+nicWy44VImEu12PYRw
35Ss42HUIElN6nkYV4y7PsCWy8L+bVjhdgEjA3emHVBFQKKQli/l6F1d4L9R5WBUkPfu/P/Ep1Hc
lj7yZShIlZ8GXSNZEw7RqN34KZ+2tlQ+8zMd4A9142Z9h/5186ip2PES+EqJ/GGv+EPS2BOcchfY
g2V82yjLLKLSl0LAhvPlYn/wlHHG+/mlMc0V6gL+3P6FnRO6MSyPI2LipQeUSXwjrvbkWqIyXITR
DWlE0G5GbB4X0pTgvwfujvLWhajONG6V+sA3lIzQrl/v+1dnweKCSHAexKi7RefGOly30twVTl2+
lHe8LfW5IaUK+PTHtdbPf0Rv0qSbpSFgX+QOLpTQfNxthBArxTNRE0lNcUpe+HK5Zbql8lGi2/3e
TM6bwrOwDLvDRFVvEf0T7b7t7RFaClPvk07Js0KqeayCNUtAryGYhBqy1ZUS4tog9KcBC/scqHJF
Lc38+BNyaq7CbCigYbPPb4gt10TTn6GI0YO59JWD2hnyraz6Vvdh5oady69aAMLxG2DV8UfiBaVx
0DxIIr+NHXyS+uzrjFTUPfNGkIF/y1M9av3X4Q/pd27+plDOq5IQmYx35WIrq6NxSQY2axZW6xFn
Buzi/1urTTbw0lZKxQfnQ8w/GLK3Pe5LszmY6eaPmvtRinml0iKbue/0/qfMcy4odODmujl1NX6w
yB1/yh0nmAsJ4KRd7YoQrAyP7qpO+KYBxj27kYA8H0XDmksgI97QTF5VQB0gsCYjYiuDNOz7NvpI
PNkN4YGPKJ2lmArlA/MWuGr8TXvuq5cgH5Jepvm1yZr9ofiCt4UFRswiLBT3FgT1NNAHzxGt8CyS
uWOxYQP6Of2PmvYmpP5JkKGSbiplXCxc2KBlfRqgVr+nXVvncHqXpcSePbn76arwrmwKFjWD3hvG
9l245ic3dGkm40tJKux5mD9Sjmd+P2XNsOFHcpRc6meRBxoccxZNmLYGOsOz+fhz8qb2trmUmq0P
l0+w8eC6lioyxUrBjOdGQJZWqn+VccyxsDU0y2HTbeXJcdGcWSYlfwabGlGzhFYckkmRS7FhCIJm
heJicyqgsCCSiCQZE/x4n4+v/pPxhplL+eqWmoc65GUvD3G46FLLl3jeclp8Wq89Km2DVHNUanoX
phk6tNytibEwNy/+wcWzPkqpJjyY44cc/GRRzXriMU4Xqd7G3Y918xFvnxOSoB9nqYrYAnKmvmij
6SClsYnjAIitzJn2TFBVza6/gb8g+33TXZSuQ6Hf6wkbepgeXcLaDTWoC3fv2WwgakSABAAzHQ9W
S4R9XyJJONVncnlYwXjalPYXATsa/sH5pZRhc8eMOjnvH9jOiM2cD0jMfuKZoXC9RC+wMTefUfm4
prRITwf04WwIwYuIzuoZV4XoNWwSh5Nyzw3AYFXkLpWrrgiUrKzVa1Y4ZfO7J/qzM8Q42+VSJboE
lLq77jB31sK3V08HgxZbwf7b+hAUr5D/4DTb0ec+tlzo5Dm7kgqouV7NoOZQwrYgLX37D1lLkfYs
ifFeVmfLj5vdazGlYaJRQB5xb4Luv7ZdOU0V4JpP3fhHOwABKXgiqlm+A5TLAsOb+FSZFHgaIg8B
Sv0eNDJxmP7eywWZexKUUb2NQF/DFJnuhZRlP8equ5aVh94G1LxucbOykIdQu8Xk4micHXlb4R/a
oMMzt+QuZETZTeGfVHKMfGUnUVhIG8Cu69lZygcz9CN70C57AgmwgcsFO/1uRxJNrGST+rZBjmkf
pXsWb7pfzBqi1M0ie9+cHpqcOqUu2ZA/bvwyvV2mokL69bpbuh70WvOsFoGLsdfhPpz1aY1SNJDL
NaIB5rE7wVr3UYoxrxoMnXaXz4g4rY15162Rur+bQFzoYBPi18tY99kyUH5oz85rgexbMGSjDH9e
rO8j6WJimiA+wW6MGvxuHCATgt3dIt4ywZ0MbWb7pUgtPF618pQm3w+rcdqFBo6Nega2IItBN2+/
KR42FVogbhxJJnY/SESETECUWZRqvMbO5Rok2M4Q0Ig1XtvydY5Oa0PsISRi3TOAnrhK4AJXYCED
0IgMYcxWvQ7rdzNu+1xwVM0H1ZvtnNJkTiykj9y9AlEokKVuWGowutWIUBKMttlN+TiDI7x366zv
EJXz1tl/kmoTpgG+xHlSUp0X4rbH3TpIatJpLbkxJ0GaJVYvf8K/2ybVYeJdjb4biAJTMD0mwwty
u1mReib/bFk8ktXZ/6kghL2f9GFzK3acdu+RSwPcGyMQFCtPFjEU+DEhvmAYtqsSSthbz5c3OdFm
A4SL0MBqqh/nuM2TwzzH3+6SLSEQ6zvaIUBdSlnMm+0CLeOdAoH1crUB5+GtXaJEKMrOXo96UkMb
VnuQbcbV5nkxGhwy2VE/eJOct3OB+poCH2HUDikWCGG697xn8W4EKKPRtZ1w7rNuJXdXt3gGC7Jz
fSkno7+UiJfnrjcnvX73KaiRut9A/8joYCsgyXqhT7aqNVbCu0oGhc4sjAjlDASUVnDPTOfXCP2l
PNBFKtv2MC4AfiYlz/iZOwwlhApg8TWa0WOQepW1jCqXG3c0O7kTJiLoipqycByWRqqSxsFlqCcD
8O8H9iO6kFWQOloWB5cPoegFPNxk5AXOp2qXwK7JN7d+mVFRMXFQcxK1QUaRd9ancO/ALwmqO+Pi
Vyis/3Qx2T97FnRa8hOzG7hymbB7cVK29Q/95jCw8JcJO3NWMN4m2qhAQayY04xodu4T4Yq30XGg
fxk+izCVwL0lW43INf1b0yM7PgAneJW3mblNch23UBVz1Mtvl0spx0RBuYk1cK3n2OsTaQE6Y5BT
Bo42/PVQv5A7Lah7cH9afd/VBocWtADImpYh4mHyIwN+kQw3W/BOEgNgw/ziTCu88qoQ8tSMk3mX
8mz3GRi3ME8va6lUvfox73WWjQ2KX1Ls6qqFGT3pd/aWnCyD/f0jXy9Cc1FxuuPzHZ/yPoM2YGr2
PkBNB7q4Xo+A0E5OFhZpScv3zCvAsGNGtl5gSpHb2MHeM3MgiuXzPtNIKVQvYDjsnrXugwbH5Dk5
nPJig8AR3Py/JFbPzMz8qtpfhsi1MMUCThyxZUB3VMTMFVQksfBl/gdYPuxtOdEU9WlFvmzbUtc0
jpc9T24Q7DsQDLX0vZy/MzElpNTeidEOkxZJ0qzjRaYYPXjR7Z+yAGZuI8mBwZiMep1rA0gCKCoo
XXaay9h2VT4ldyOjS+p18MUZtEtsQQhZNBaBQgxQLpkTjMUMYqEXq++wuZWHGtxNBNIHxvf8pKrg
CMAvxFSgdzt/rPJRK74TEUbLlv1/TCvsTGuwn6B0dBZO+NnBlCE7l0RepCRetxGv8VrVQuxfmfkG
0+vT4TH4DexEARVOluVVadN2aAE8rBjrue6iDO7ZgFCpkAOuUrT+KQIa4LTsU5kJ990i0SSzKB+y
HgGU0vozoTsiBkX8BmUsZtqpJMLPjuA3+m6cfLsGa9KhEKKjiN+EzcQI16e9XXTZcV89S092fO3V
HcjRTzzNdATzanuAaZUdPlPRVKYWKenX2oQVNde2YuQ60oxQtdRYS7/3DF+ExQ/FisbpX7B/s0Qi
lG7+sL/MmCzAVeLMn+/YcuxNAetbrdqYAUKQ4LSVL9BiyLe1pQ8nv4H/3XGjpkFT3OS+kuCdQ+1a
eqhp9NTzRuzsgI1bkgMbqxsRfr1uFTsZfmajNI0xQpT6YI/XUSf5iuyRu5msFIFZtSSHypb/+R+b
58wLWqohfrFwwTlupFNAS5n8rkyt6dIqCrgC+3oJPiLlHokp90PQTMPEPE7cuzmBROVnnGTOXB62
y+TRjKTCqHapsc0hqX8MwdGcXtJuPSxY7xHofzX7E+ifWCyNFQddno80ofuB4/ur98Gn/wVbTuvk
zyl36l1N06auA9FahYf5vFI8kEdA8/yvENCO9/itHq6hp+e0Idacm3odgrlesVrYsQGi9hORv+Bx
C8ti2FsBcrDKX03hFEJb3cHe3O82ZOCIakHxj5MgXfAwonke9j3UNoivkvCUsfGl2oneYVnK2TWA
/qInNYNHkJKaLUsIGHztkp2Jj2Shc4IgvYFqabcaBxekceTUMFfoLZwXaOrH8AzOmcGwHq4jd5P4
bl1Y7/BCi/EbvjAoN6r+YOydeEFzL44ZozZPgZbMNxNmAMRGJH9S3xjaa26WzfpbvWfnRb8BugiS
sUAVgE8s71VlbLBxennJgZ7gFPiqTlJqgj9o8VcoAaUTFcUmuAHrwxER7lDcy8/NLSL7N/cIEsCS
IO82Xk5ok92Tzw543kL17+uOb5aQEDxse+cP+u+vAn1Y60xWcmwGS6JqmaEXa/OKHSEw5ZPjuo9h
o/hYzJxvNgzWGIWaOMUd4va8T9/DDnQAuKS+c90MCWi3w5fhpj7AV1vJhkZuwbLZiZnaULR2F19X
50vnIkYfK44KIu4xnOJWUvPxmF9LIuhFoVKpdzhtIw2Ure5N0uoMAomeJqZfA4lsGtK8+TfUs8mj
eHFl5s5qkQM5V3nbpmPKkXjkwrOAurJ4MvDCwot2ElFaph1hocLZFymodGDDgiSsjYJlBXU+zJNV
bqkUYZJKI2KTOXxC9gWCwvg7707SN4+cgzSpyJXUNdAcz9DsHe8XVBbi/k0sKtUh3gcxqYAXHYbN
d1jZV3/KkR5NL6T1ecS0jD0NVRNbDWug0mVW9c+Fvx6IMg1yD/7U3Q3sYzSgVE2n9xe4P3gCV3Na
XBoZxGuaTFLMiU7yAyf9X3blgbotfrr2PtD3iEsGKY3BhagAU/ueMlCN20R0A4HTOmx+aZz0MC59
sh0zY6PiZO/uEb55mczANXG0fbN5msF90L8qvfFTvw9+Jgdr0QF3yRo2Rm2d5DzVTgg6WSMeCiyx
70glql01nQbHWCkvHBjsO32/LmfVYIgocGY+G/wIGT0zEEKBWEesdA2YiJx8+j9hIo+MlD3rJK+U
QXXd94sSlD+uy7NU1oi8K8+x8Ypi8Ou3nuDwKZVIyODHoV9PpjPLI2ZBnS6xXx2ZJvP0SGQk/rr0
p637YzbxU/JbgJkNKtlCyed3KVtNRuuk9BWX8sRrKFDsu01RoTBwnDHAwtqURWQy5uExZmqsrOGV
X9yae88j6Pgr84qjmTS9Y1p94joLBe5f5DyL+G4IYkdNHe+vZp9SdhPRKtt3Qq8YkcD9iB7tWEY6
h1jrDsv/pj5ycuHOwbfVK8daJK8dBtBXYMfpuM8Z35R4mBCodQyrp+4I/bv5QDw8LK+13CaPfRw1
PND4SzvXl0bcof78m580Rbh2aXY+J7vvmMfnxh3rvIes6PR24U4uMJtq+lDyd1bHXzAvjSDvFI3Y
1gJPh8MtcMtmD8qWYT4KQz+Kk05H4Vp078HOSSrpT7dbGitLG8P/BdqD714Bqc/Qmcru6gDHo1di
c5TEG3XFZ4QigRWZFG3IZK6/5/+rAxTd8Q2hvFMCyiOfVg9GRV3PwzAVqqYiQ3GSUh8LcHPqYKb3
4WdhTACG28noU6XrSu3UTouMahxoyMfgbPfDNrlVTxP5CLtc6VOFzX23CpjmSULXOfasrIJErGGb
8/gXuISAjyVWOZobofMGhRjlRLjHnFWyMiHX7MMxviq4PqNFC6HspZc8aY4Oe//i/WWjNuFp31DD
Lywbgjbd4T504C2WOnRp6gHWA6/bsQ6WsUNE4nwXL2EeSfl+A0nXpaw1wWK9szg+ykp11gZirEIK
7OOXkwCgKDTDnF+aixJEhEMGGp1mFfkKLWkMBXb+zeXomkQFGXerZO1t9zsd83M1AjgMO6VkJMhh
d1QLKt38OUXIfsdeyWTNo1EAgyElsoyFNay+fPBJKQp69eCTx9QFMspacHweAEYPvJU5AlVqphqS
bPfmkvmp7zAozP0sOm7Q6QYD34LnVKX+dPHQIhI6m0LhNAiXFM+plCQJEZP0R6QBL7hkWo/7NCXN
pUT8VINq6Gi7f9vPNUE0o5TOSdQleCOJGMgv3Nxe4bzeYnMRO7TuSOrl4OphiFYwLRWzgkG6yLn3
bFiW77c9UlOWkcAlzLqh7hH30fCrxrZSQsB+cyctIXBRZlh4OkuX/Cpigu0l/hzq7WxamkCkT8+4
G+IrWia2yFdSFoOLg9vWUxF472G/sMajm79LJXe80y53q8xOReQust3BIpn1vlfdiOYPubNNs0aq
2RUfXc9BphpxVBsUerWr8QBmOnFVy/dJSTTyktJZoHxHR9wQcb8N1XEi3BqL3hkz4EjPQLTLt7ME
6dxhOv48UE/jGinrmWB2x49ATeS0+0oyEEF4OW7HuYNRu8MX3qYeElaXU+98UoZqrbUikMr9RfxG
OZdXhvFGeGHzdQvba51LYuO4DlD+kCOB6bUmwg/uJLYZn+nLNznNNiRjEzqu6kU06TIlxvcp5+qq
/g7LQZeRCkdItw8noc4uUPtc8eeAYy7P32f/pGakMa9/qgpM3Z+rKiT2aHLwxaOqBy0dtrCcsjZT
0q8vNX/Nzr//mL8KfiJ7aPjLBiKnpVDgQNI4kEkMnpU9tnkT8JJKDvShHPXhpYJ2r5PBmOu9CI37
Tt9TN1YhbvZlKCflXsUBvE1lc++6nsFEBlyLFmhJy/WrH7tWh0w9kq7OksjkzyQv8wxx2nR3CFk6
rGRTNU/yNStk7yo/mp55Zvo8ppmgbZwRIA1WqL9E3da83oS9mfhUkdbRxB85tvR3Trr1EZlntYf9
aZcHbHqvnTj2v/UO1jxjUR5TUbfm14kZ2QL6ZEl3gB0IoMJUYshpwr00MQjOmMM9vN9mdENr+uFt
RqT+ilbLsdSt52fv/fMT/g3m+hVLLHqBbTnh+ovHDpX7r1ykjR9pbIEEiMjIIGyP7d+ugBY1diNH
G8TZdvos+j8OpA6RZuUKiK9FOGDt5NtdZUKXfHl9HWR6nI95CQXVItOHJ66b31io42ugij/btXYa
GTEuOnxhIqNaokA0hdDGNtrb/yc37J7V19X3a2CeroGungFL8z4HVPoTzomqyHWiw4HuO06GBVeX
pFB5juIYQohjyDz0nEBz7bW3xPvgZ4faJYhJH7YI4ha2Oz0q6kXJ4umBMM9OyPyKUola3BBEQJg5
0G8cymOBLzeU4i6WvLy9MKPVdyCMGSMSF5lSJiMz8mm6pxyVFalq+Wcy3Qjt2jOFSC/KbfDEUgUg
sF378ZCizLQzv2Bs3jzOB0D3Kz2q99oefohrOP0Np2tdTC3+m/rYsNo9+1uZwcIWuKkhpwrhrw8u
U3lbFA2oHBYTBdladdpCvcXtMs2yOoZ+YGwz9cnAyX3i0bxL0nmGItzV8GGF16YR0kd1yGGmHWnr
1Ob+oHIELU7u6wK6u7BqzZ+kLofA2eqlt+A+9hFQI9pu6r0R5pPO125/wzlWs1hu7oGwR1tJJEZc
u1O1cTpMDHNmTdUXqklFEiUPuhhyk6fJQ0fNOIW3aeI3r0ILfjKEBUY7tJo7lM6jra+MpT/D/PpT
rVfB5IM7yUd2lK67DQ1/Nk9EJ/iuYCSgyIn2wwmc6naHC3IPw5RHM7tX+H1i9TrjxeiLEGwsKUeY
yZOx0EJcahxGCbsVb+oogYzyazTtOstkXALRoQ7T7UJXhmeeXFuBbrChKwQ5QbecIGgDBfiaj3WP
s7HPfZ/nuB00n8/H6iB1uNp1DxfQkFy85JJS9CtBQKdUL655ljtO03vJvYNSWeux0UApyb6+tuH2
pYRefWYqUC+s3aTIyITT9k+telD6kxUSt0vNYZNY0EWfln9lJL9S69w5z1J47RG39yybGi3OtxUY
04fDRwnAnqSgl2t8hnift0Dnef9rKVB3qvxFxUMvSxt90wJf4AIWtL7uEArAcyx3Dh+mf8wKk5VX
BbJHubfmVTMZsdlD/p9BFXIAyW4Wu4cMfH+e9aQju/798FcN2FDR4nPNVNQJqJ1APBDn1Aua7RaL
Tj9BYca0AwXflfd4dfH8z3ULH8DwDwYvCSpAHnD8U7COUx0q9JmVbco/phFprS6dE+ZLD81gAqyk
jUnutMBzbxlyGKNszGHjbwk0Wsk10jnPXFopMlkAjcR1exmQUfpWIYubma31IzLDYx2TwyCdf+Jr
6cdY5pP2xiSj8cE6T4iy7qyJaQYPx38LskRl/hR7jPaQnZ5eNOwGaBQF2NaHy6fWQpRkPkazz3Rg
AGrifxAvJcTsvNxkrdNNR6B5lny/Wy/YA1D4a9s+24a1Asj26GdjWLaSdrPe1bQw3Be9Mkj+aMFR
61/gnAiJwblzMXD/u7VNbX6iy4LRQE+YWV1ow9gIAjgy6bTsItWBZzYd6PZCScXELd4Z49y09xJ+
RCBqDCaV/xVDJh2qbZGHQf+Hxb8XkKMGw/WOnx4AttVSGW2xIz6v4Kqu5FTHpsg0I7W3P6WvBHik
QG9/rPq1SgjrCe32Uw+gyb0xFsbdibum/vxRxIjoGEwHCh3nRzWS6y2OfasiihBxEI8l0yr/Gbn2
M2uvg3GFvUNoEh5w5kcXIkxdLmvP1/w2dQqcuT1i5WHwabtsqpM3J9ldt10GPmbbzWZDthZjljT+
TbCorZf12M5lge6e+XbpJyRAzDKCD7DYZrncwC1kV8lIz1VqidODy2V/h1nS75bf7saQoFvkI9Kw
KY6rMamU0gBL/mjRZEGW6eoYrxQfH8PFRc04AXJFS3pITUQkUEc9gx7pRj/4Azy0camz1YsAm+YD
34Ef7kAKjfHAnxSsSGzGjiLRnSaeGhd6J5ei4Zjue3uVL0A+hrrcPtHzcTBbQxDvpbmqUSsoXXNq
cNBQ3lJU/vw/ptq5bI14fL034+9f8bZWoweGUqWjBwZjFb6Qu60CjBlRbHaZt6W4/p1JLqs63KAY
RhJUToGGkZW7sus7rFr3PVSwJgm6F+HLTCwPHazWebC6CAd7OrB2ZuecdRZ/EpQgXoTBsJPqPUPi
bd1OS2WLLVCkvW3bw1oUXXNB0GN8hjIyq6vA+EX5466aXcPJSy0Vseswdp4JArcGI1gfW7cEkz5H
y/xrVb1qqF+l3paHpGxNIBUagSkmdltAWEp5PfVQmJ0Lm4tdP19ntUpXBxfYpoylTDk3axUaP6F0
QFyE6EkS3yY+pdz9xCVmLwcR3HS/0LClPOoM4DLA1siN8itPdQf3fRtqGOPtNhFLH+9x/HWllhMR
+JJpai08k1gB8H0RYPD5lV9I8idG1izM9yTP90m9+ywX8/ve/eGmkalD3UwWQHlVLwxU9nySo8MR
kfEBTBKM92fRBoJa1m/hNwG9ADp6oI3Emm9u/Dqs775PC8UquHdeJIqvlSiifP4HE7LcStlWjOI+
vJTjqlKcujptkhaOGCTUmKo6wkvG9+MIyRkKIzpR/AL+6jfW548x1aIgvS9XAm0SV4wnx0Bv6QVi
WMzRCYCjQG8bWHjdg/kVyqMx2veOs9cFUnp6JDgK0qJryEiI2/1UNoij82+xfV7MEheZqAXvdy0M
5L61i4wi0Gm3/2bxFiyEiY+p32jOrM+CRLpJOY4FgwNLHrwTU/eeIe4jLQxZiw3B1I2QnTK4/Pje
KF6j33wEeoSQGST5YNKFL266SVuO2YHGnUhWUOpkiPLnS0BjIKHMf2VHEHwvaoMUzmiEGY0kC6YQ
Pe7OaK6C9XdV1gmoIY8Vd9QFtyz/axOZSkUCdl0nPLkTPdkUh33VY0znex4Vz5rpoGymj8hby2A0
gZ6ywnfWM4BZ8CaPFaiAgMEy35jGn/k4qLP/LY5vSVa1Nln3O0nCo387lCa60NU+xVbRwJy+iSH8
wlDaYdRHUbtVBUSPBbisH/7j678gIH4kfC0KqtOKqT7g2NS3Lk83XElkFq3oZwlxGiykJqVEKauh
iyzlQBnGW68do5JyUXSbf2U9GoyoDOY5IgGrCKES1KD0s2C+oenp0XHTY5LAx45n2+I6WgIGm/cx
LohlhR2zK010lMae/lvx+KkjgTR+oVq+7WL6s78ojL1xQIKbEoMzaAobnkQRWtxmZccMDaBBeNSb
BLp+3S10oTNK+Tdat3ylEcS4NSl4JqOZjGOeGcFV939WqVJYx1+mlhTtlAOz4cfKoICVAIZZusab
alTSSKQ6GUvpNQcpsjM2F75CwzpXNyYuwcANtued2xpM4pNda8HY4rtYpyj8uiv/pThXP/SMqPKb
lRwscCNqa0+shKguDZdKaB/4QR+YN1/nisd6n1xSYNLM0JfDuhZ/1AlsyG4ujj1FuEeu7X1xfMx0
93QmMOUZOcQm6hVHbfxEft/iCu9bIJaZJ7YBTH4mrTbxBsd9B4mOMAcLgDiqtesjwZWBH4OHwFqK
o6u/9DMEwhAH61hAmlGGRQzatzhYaug98+0iGKSnZ602qMEbcyVJ/K8z9Fd0Pef3mrg/6z14HI28
tbPBzkn7qALLwmPGlqYnFA+qxNxHT6mIVrNoGIe7tVvDTRDHIs4ceES3qikQ75rWSCMxJ1Nvv2Jx
kcgi+KlEqkuxjvBNcxVcluVemegc9GCZmCtBrb6ILs15QocAw3OTmh3idxd5yYP/tgMm7DFYpwUw
EhekQxBf9iELPTSDpmYvGEC5ePMrq/Nd9NBIozA1URPOeMQYkDSvTNAwUqusqqGuIrVWNwrFAQn2
PmgL0A6kOVXMVlAu0cV7Y0SqZIzTbohZvHpgf+hkOxUodb+BCugl+QRMILw9THZmnhJ4XzCwWWl0
F34+iFdsd2AvqUpbnWXPb+/YCMr2HEae8pLJuBqwaYc5RQqsE5I/jIm2o0q03H7oId40UMbKqw+D
4FGI70YlS4jx9QsYrdWsg92Yum4q946cKn4U/LLYuDPcCuz88oaIyYPMuwuaQtoLXJrDXXbnH31I
RnX75jd+Eh2SciV3pHatgDifDsBe3OmUDUVNLrThmaLpOsZpktbsi1z2T6fD6Bf/FVUuUDlJ+9SE
rC9z6H3IcATTsk5idnbZZXE+FQc6WCOCTY1jz5P+CAfL+LJpPY4pBrtQze8DiU4wxB5jJst1AM0N
GkfmFu3XROwCMCXRPiIx5sZBnHgpDhaA0Lzh0PwZN8LUOIiO8sU+0Go4n2BOTLkd4ZljhP/aIW2r
4HsdubLwEqZ7jn3hDxRLWZHefAK1xtsQHYIgTnbl7muKm7ZGYGOldu6H/gUfcg/uRNzwJrxbqSix
UfuV9efT3qvVy/dfIbpNWhumDTEGoSsfefnOCiafIZkQc7O8E9VR3GXhAfFpHP1OusVQH8tPf/2l
bmb/f1ne85+0QcHp5atLN4CZHD1+B35VpoloX+PTEiOo9K1FcSYldWOCRmo+cd3qCpzvV/hNvnm1
Ru4Ba5TiaganMSlIhpbYyYvEdgYljVYL+I0PhT0njhqubZeROxK84KZP3cu1fvDbdwl9vJjvcp1v
BQ7uzh00zBjGz9Djj1WokXv+dHVkL5w1MwXG7ptGIE4l94krK6K5WIPE49g/nHH3bVrEye055YK+
TNXmeUTM+7SAA97sv6iFncWjb/tAhZrzy6BHTffaOnNl1igQnz9DBNC7E74dQTY0jfs5RPArhE+S
vvS4kg8Jt2Bv6paH+Xq8KYAxpXeixc6SBW8XB+KIPe78xvQICS2AQ6fYSwvLw04T1hcVckuKQLcq
omJfRsSQSVRRBzM9yqPTZ3jqeUXj8fiI4fcEvoXFrtHNXpRadUpBk7lMC8ZTLgVDJfksgbdiy62q
d1xXTADP+9sl4nlng1eE1LZxU/QATIQ2mgqFvQZ5C4v2n3WKrjg7DO+2QCgZvd4ZIodVFQMeNCvc
I9vr3ww1+6GDi4w740Gg/5rXD0tYXyGFND2yH2zyBIJ7wFpqGZNh6PNNn8ONYscYbvQprPGV5OiJ
y//gMIcFsKbniVEPTSJs5q2EsmVzPPI7X8rPO2QuQmNOkS60tJQXpQKjMKH7/Btj3lWSCfh/+mNi
1aZ8HNUJAe4UrzAjyCcM6etEQE7oYfMvD0RhB3K7aSguZqCSWTo4TPkcyVWxANi/8bmtORRebxxD
+ng2keJ9C7DGUkCGdXYD0xH/dAnRxqMrszHRsaGwJwjUfPkBdQusfxPOxdTOhIvPOpb4RDmNmcdt
e0Jm0ZNiOnPzZcjTEw1rt+aQT5RI1RRf5ZOFWg2/sZJQdx/LN3WkOh2/3MbmRAm3SW6GqgiKm0EB
0G3gwtu1f+q1eje6sie57GZ1IpWaAEOchH8L66osVntV5uX2IcuOSuse5XJx4rAFb2lPHZ6SS0mH
hykR5aI5jtgcWrVGaxZi2kHfQB94DuKGEwwv32ky6kt7YLdbclJFyO51EWfeRfNUnlGhwPGjPEni
YFq8Fn855MgHTtrLQQVumhHuJKlGS/LoyDr59RA1XOU9ofyE5FXqCO06sMV4cuZMYYDiLPqU6L7j
bHd975WKNIb/xH3XnYLymmBB3WKy5gMz+EN0azuL4em0DMOLnyk4F8/KHYGFG4RiQcSfmN4C5Ijq
hrwAF9fgYs2HOON3be7tn7RtrPEUmShhDI97fFE1XmnRb7AYX0jUXdEiEA0Wm3VTcGy5pmp8Clty
qKzmQJHALjPSW438VQps7eVESyUMEhbArTAaolXyWegkg+UaVN42/WBDTo4vt0prEa+xyT8ST0uN
FVpCHHCo55DoYok9pTuEBjXA+UoN5vthUCAhqGvU9OsetNh0Sqino1j6qqxipg8KZvw8jJasEyMY
V0bKmRd2votQZlDVdGlcrp7pFjjayl1NjnOlave6IvR1Bm22CwmCivUPeIugQpFjjLjN6zKu+NRr
xKzaflLg6OjcMMFLPgVUVYE0asC2bjOSt8deeoc4TKIQupjFg9r1q5X5G47HMA1m4ku304LekhjO
OEE31ROrzJNANV28sLOze4cCCZ5SiOg1A5w1DKTIHy7EdSKvyNmzktgOSz0TcE07AlHhc5yH839B
o+EjVpg9hldNJU4BXTRo6yj5g55fmHAIcljM+y94PzIwkwBaj6MItrigXBhdze6zFPa/WFhT6/5C
Ggr8mEEvnPic6qZZTa/vELV4kJ4gOuka9BYVVMlwjYi6LcgO29TfIWaqNU+dbYasFX9HH77FimO0
vhNnbGJ+3bG1C3lNoqL+lPJdOXGxXDz8HQYl9Es3klYS79JGWJfWJBxzSB3y4TAdfzaPSTod0H0/
449DtIF5uMZ74YVF3O1tA/qWDJ+5dtjFTaX3PW/tZPhrEnhZcssj8uWAsmguPUSuL++TS8/2r9yr
u7UgKsDVdktIcWXAekMKTHwM54FwnV+wdgCJpcVvQ/nx3SZ4zFjux8D+G2CcXBujX16K8+N6Fzoa
/xxjY/8+Baw58ZXziYlJ+0nLfHAsop+dD6e75OYac5NBWaIYeXFD3s8D2pyFbVflwSxurzDEeYyd
TPTp7vSHQiBOBHjD5gCcmqD4M3G2YLj+Y71b49IJx+Zzf7Uwjl8UUEFoLp5P4FtfKWEFm/XHO7lT
ulqcMRmDpxS2w2d4haRf2Iz4bYIe85HBhbsvFDzYKbMbZbI3CDtmBhBSSfmcGLj5puO0wOCTDOCM
cmCTVAUZq/+ZAyExOb2eDMsAgwL81JT7mqnNIiEwn2+EhcpMvsR2QLG1O5IFHyBdXAndhOycXFQf
akEspKrk7314q7liZoBlHlcUqZd9vh+vDedrWmKeAO2D75SA+5jcUkoM0wm/MX7RC6qwLDQOYeyD
Pt1FSkWK3Du1c/vdCOGuYUztPNs5XNgph1LZauK7hkW19XSrN4D5VtmFeB+XaZjOFFE4ocjUD/3o
rK+VbtxztJkT6o5WDOIuwywpKYLD6KtA8bkGO70WQ44U9nO94i8KPvF9Rn+WeR/pwBqZagjccAA/
RIHqfbtvCJdyQ7bnWpQuIZGW9n0Vr6gAth3mlRVWqyqZuBib7WKeJ7s1dS2/jsZQTh0WJNx2hNMu
Ghw0bqaYp9Dn15ajBTYNxHOVfNs6byrvGRLLjI56B2zLyf2x/RLkryIJG6EXsolXB3j1Qs1i1FmQ
RCi0CkVqAxge7kwTV/dLzA+wxX26Netdt3kpxkDM7qN78XqqtDS93og89y/YTJhUET3rbrHWd+QW
R3BUszgOgcXVugCbMOZZUwY7O+055PlZ4M0KFXNWYxxnS8qk4aD8rncjhQwpLodvermvdlBiJWWz
Likktuw+xlpsavLVDeKm4qxSpCrmbrqrCmnDuJTRlqjLOvFZVsr8HXfH+waGe5Rf/1Kff6hfDZJQ
bcUCfwHhpXxYthxdwdPE0OdB1Xad5s9fJ4h2LhR0swdirZC+Fb6eZYo53boh5Dr4brhuhcPAJ4my
5PQfw6TzZSH6SXCf01MCsC7TYOsoxn7PyF6GbUlm2vpLUka3HvXMg58ncjWqi5x8XCvdGWyzS/i0
IkQUJsmuJ5f1t8iN2vWBDtr0MQ4O9Y4TC/MqUjsPzm7cZwqgokupBAb5IaS+jG+761BvFY1ht2hi
XjUebUhhPHlzNkoyOdWo6R+CwC8HZ6N59LifXEtWXA0xU3kWASkGGS1cbVxeAUzvvfU9OksGw0mN
lERWNL4oUZqxWwFdoNWV8OTpwXLxT4DTZNGRgTW0LHpLTGJ3yZwnMu02JGudaP6rUKPYMErpEnxy
Lmulrg4QHwixq3Q3vOa1zj/55hQ2UYG8z1owLS4++Q2QTSEo6Wolz0hVaN9iJ0SyygzTyzwmvCyi
FE1qokPcXbRwrrgTJLaNZEGKy9Z4wpyk48iuiq0fdfqSJUCXSYBXf1zzJjf46dQ5kYI0tkFCr0AS
q7MEqeR7N1D7+bNicQSFc0luAuUz3rJmRu7Mfq99Ath4QH05Mm7Fl6K2/fj6llcUt3FhomU4StfU
vCoPZ4CPbANbaQCjd655U5rge3zKyn3x/WjddmtE+gjuCsxywW6N5A6mPPYXWhkaF6pLtJyydtB/
uVKEVW5FNkGgI6zfTgs10e70JvTQTwwkJKeYTFlL+O3KpTZlC1QRYPo1SgETrvaF1rV4/DS74ukj
nWeT0+cSA54l1kySCA0mR6HMMD7B4tyZEmlLMdLbguCCfRg1beecABuAvTENPgCx1v5/ToX6xBER
nkdAVlbTB65kMB2lkoDEfclRT+o8LRT7VO2BDp5xYZ61pRFcA9NN+PGzHgLAC4tCAkfffd2x2zmd
Coj11Xu8pDtaWraFMAuP8vi0EmrLlN66e6QTnGdEiFpckWu7bwziOzGTiEMZUlFddBWHaJrJP52W
sJuWotf1clnwU1ZjY5HGIWno3FXbTmqbMlwv6//vIEB2BZu/Gjy1Lng2XObgM2BYo4eHhfSHhWv1
v1CJp+WyyquR2x6Gig7OGC90gRZLJxMYVqgi/Y1D2vl/mak1k38VUl8X3HirpPjBfwsaFyTUiO2E
65DdaR5I5euq7yQY+HRhw+3Tvw2OEzdd1YMwfNc9SdqFSaXW9MYlVRsFFYr2BKEwDjoQ76CecL4A
D1RddxJHpZZKUwJ5HXkJ5KnAIIbr/njeIOVbyVcHvLDcK2DoLWlQFSvlAzTTqwqf1+UwKRdXIqa6
kFPJ01kctzkXJZV/jt0wHo0e6Qeh8gjWMXGBhyEjANPZPr84R0HTT7GTtyO5MLcJgqb3M6UfXERW
QamVAyYMSACi+4NRsd3qiX7haG+1gmPv/MRy578/eTyumeUyi9hAex8pHTMc7haaCY8+Mw3T8Gfg
+lMisQ/P3sYC0F370HZBW3u+oG1chLHK3f7TWpwBKU2O5RCvaKsuo5kup9uEGo4lT8S2sfqYUbQf
yvW7bhRhBGRDIAEf8bOFS7Qd8adYYAyUHx8CJkks+fvyWZP4wiTu1BblXW/SQkfqB4CM87MTiOfB
4eGu4wu/WEJwX0VvldIWPafBCFbp8h7x0xjgDELQK9qJYnnR6kvpBrwHiLDbq9sG65/bwgjFITH0
NCj9CJ/HFKpNNJ3wAzMg41o5kY/jUpnSOGk11Vq42mv8uvT38CBtpQV9bzNTraLa+ANT3BfwZCLX
TERmh3NRhuT+uNgWV/tGh2owscT4Z9v9C4VkR907P8789gBiPXvu3tVFaYnQ/FPUL8SRhguCXQaV
iMLlEp+JAd1zVw7dICnGGesDCRxyT8lLYFjJUanW4mVXu5HFqjdVvj0uujzZh/TpF3bINFAkwTuc
pIa+ADVo6R+g8mTMhiKPI28NnMYo81dg9VYnNZQ/7oSFCjT6OzKOL4habydJFL0bHHKGSDEwJJLx
tU0WSrDXQs8RhIfzknVkXHrNK5fsk2FtLfrBTnuC+FidBWNiXU5wDvmJ3JBMqMxUbVwBrArLGVfA
U1/tRX+J5ZGu8NIYfp1Tg21ODgTGEFuoKYM8+jPDR+FCFL9jGaYBjVH11C004DfBpWd11XSQG009
Lz3XYgllZwWBS5yNIB5FW2ajrKHizExM2B9v7rMey7LrmwzbTdeNvoZcrwWiiOIwWTJRNemilZiM
IICJyQhgcwHmCCCfjwmo3qgwLKneiurhHdmhK+KogGOiJKsvFNDJS0sBjaJNz2KlGXbkkdEoJ2Sa
5xIRPT6oZ1MjZxho0jLtzwqUJyk4YAuqkMhNUjpcHWHOSgqWTjUAnz6AXqPQUn8K9+Q0J5FNvBab
jZ9VmibN7xx54nRMEM+Fim5W1fhG+5jgTQzvGSi10gIjMM/R9SJ5Hq0WXewi7bBpNiQL3G4gFIaE
guJjxWdhr61bSiMDGPx0vlbsN/yExSZTRtxjuQiw7HpFseXEckZ1QU25Szs0BQ4R+yewqynLmiDm
izCdhLpCaAqfZzmULsmeSKFhcPIj09kwdZoNZzL4Mijpuajn4aBnCd5R75Q82Lo/KBaeuQHsdhh8
6/R4dubE0izNbte77OM1UC5OoVMDHpC4DlvT70b6Bjvy1pgtHSm0g1+w2R841GPIIB/+FvLnl5IQ
kZy8XEI+DU3Huocc92+beHHbNsUO1f33xMj9qXaFgYbNUjWU7Es5OK+j05jovfGF32SPcrfrvKQd
HHafndDJtSGVZtaaaz0AmEqzYOHnvajnAWrRoZHgdY51aWonEIn4GYMoY4YXFfA69MIv+2DuVzjg
I17UPkmK39PJAapafPMQojVSVqvhOmH8uqYxYJ0ICDSwWXy3bOB2J5N3qSjeEj7T0p6FG5gw7C4U
f43UjluZ2syNIMFn86cE3YaW/UrUI3ibOYkEvY/Haf3EFg5m1ZdyKPTNIHiwGky4xHGVmkz0HNIk
/kh8RQIs2q5FD9KLW0G1BOj5TGtMv6GVgJOUzFjxy+byA9vfa+3gaW6WXKlqwRlI9ycMvZ/gkk1l
Bu++8CAYG/7YfHA6NZdXYR6Wnmif2XPb19obKy3tRu1PXwJphXoHk6jRI+1w03pu9Aqvks2W0+68
e6lowDz/A1Cg5p35nyufsER668y5iHhOyYcYv1g0mJoREPD3H5SRDiiogMHa4nUi6f9euBEX/+KY
yGbtNwyqCCgCDUfv5BkK1nfq+XCkjEwv3hkkzHCXZcxkxs7Z95PREnu45FW0invQDluhEHiX2syZ
Uj4+WnlstGWArL/gd2fAMp6VSZFUZ71VsJMfEJ5w9Ul8sJxdl/C1ndqrjMqK7w3Q9JkOG8qV75gq
NYoELTju87d8wqgI+BKlxsJthdCj7qFzeRhffPsBbFwC9wTx3PoDbJTdxTjUsb7dxWpn0RR9UJf1
qwo5VFaCzqljaI0dQ0URhivwD8c7lQa203VKX4IiQSq4nNNzpH8GnfQ/PjbeigrOpButxV6FCAgD
CBV5nJtu9pUzWOOxWjBHhf5J6keES7sxDYjY66jCe2ZOr5vIx1G4ip7zZUD3xkf/uITuOYFWhWop
fUtNg1L2Clu1+spV+0hAkC2+zcpYcPbuU5az91GnWemgweQtRR8J8HMY66s9yGKtuTxP3HUtdYyE
r4XScqn3vWOmLNhSFCVIUem/L8qWwWEf7mSyCGvt1SGlpPvDPxION2NZnsefPlQTkpgcakWggFpO
vG4OX2Uj3TmTb9UAT4foJXy50XwDnEenpzq1Ya/A69dQA4WSqlSkB9axjAE4jpXBq/VWhllw90z5
crD3/BTHlEo9ktYUNEJDuyFLfEtBP2tkIaQDeElLb84/m08ubfHlcU90J4QQLtlczKX9ipPDIR1L
uuyfw1zzlcYfGd6OAab+iNmN+y/IOfjhFVZwNE9A/S0ikmqQzcIuduniamHDxO3FfiktJZRV1EGh
Xe9Du27lvPNEy0IF/kZ1UtOiR3DwCIFaX8jMQI7vaSebD7l+S40lB5LFHePPqxGE8D7ghfLR3lTR
hMicB5YKeo0UpqFtC6g8rCg/DDir0zBB7aq9hVx/gX4uPVwJ3Yyf3StrEbBkuY5loqvgh/JslkgV
io309fXRd+BYmGjiQm/wSL1ufM9VdHyhZwzkibfSMblSqYmtY7zHedSF4Hg0mXXfB5CFE+VMyU0R
lkAJeNHSFpYDAhV/aAlIvsvC5QtPIWqPBcMUfXkryOC7a+kyW+maa87sM0JWRFHR69yDzvQ9vH3s
blVkZwrg2FDaQtdprxqSoHpZgrYCp6O2f8BEsAwafkg/kONmEIv3G3UqULwsAuC/QK2kIWTrfZbA
T97WshibBi2Z/Uu57bii/9O85gxuvDtNjfma8rSHDlO+z63wodVy+wrk9bPvxnCzTPuUxGqfLr/g
fs8peo+aUq7uavRw3J06XJ3k73uRgmEDPHQs/tu3Hg23rnPQyYKBmpFgqy/KjclOikUrGcSJqTzc
CktpXTX2SiSdhazOH6OLwRZpeyWqfMvPeDtyVN/+A/hx71F3Clej8X0f1tIp0S1Bd07hyhBAeGZ1
7vWOnTGEjVHc95QeVHg2z4IpPfhzbfbw9KrdZnJPpITbzZy+o3Rd4VrS6vAB/vJTaOTohzxhl5rF
cBpx0CiWuBKdSVLYYeF9eFBI4j9kIYY/Ye3eShfVlJ7/rN0diB33AxxobD2p25JVleYE97eLtyms
vgdj07q8wrFh2f9FXu+AaarZF/9DboUm9+RndBoOiFhsu2tjbYgavCcuiTuVFUZLv87Ef8BVIGYQ
aYvAAXEvo5KfPB7Zn2j4b68UeM/94o7i1jMnUm2r/J5whOHA3427RjdbGi74Ib4qX8iSegWsxao/
ypyWvvxodPDcmvmdrUHzDOh6okeWYA7pel3cIlwCDxqhFkMnk3bMRwnRPhb0isCJsgNul4SDFGyl
muVRfqwx1lDl8OBQY6za/NcMQFqszm+F97Dp35cE4ps0/3wYg1CFyNy+3vz7nb6q5l2GBdiMxIMe
upqT9rKfIcp6GdAOSnW8X8U2EZJ6wRmBVa4JfLeVmAq25y3BbKYuquBtQGmNyYObxCKRJJXO4V0A
Ddk52qy0FrtV6KkGvrFouxnNMuAiym8OOd4KbwC0DyVORIIjKhdG9lfyr7MfhYPDilXtSy9tYZkg
IYONwTFuLqGL/v3DF+FHmXAFqjrP08f5G8MAk1fUBOvq0cOujBr5Kl8lgzfcE+bDtkvwKkmrrJBi
0+WmwAX+meeRpp/3ql1A2CLLUNu7jjjvTZ0fxr1MwXFc7E+s7ZL7hyi6FQRvy0zTFmEANmqF8LpC
Dn2cWwD9JesGsJkBM90wO3njO+i//Kgz8mYwpCa1AYbm4RtkVOxzbtkteJe3EE7f4X+9HFBTYnpy
JYtyIb7a+Ad+X8/WcFqy7v++FFJiLY4Kp5aJglfp7sLCebbQNUGTNoD17URv7Y8wdKLji61/2230
sMpuU/McEmdLM+ogsCqfk7srzH3pvwR8E3FYZs3qh7xYpIxTrC6bH/44Msr34f3nybMRckW8xmRU
A5DVhcnZFNEjIs8qHkD3KQaAtW0w9Gi2K0+JNpaCKPQ8dccI8kWoptJpcSTXyd0+cBYbEJVlkmzE
bAmD6tjYyr3hEGfe9wYj4+ZdfHbrqeUtc9v0/J/6yegkY8X5JbD5JIgSl4Y0w4W3Mn41Is+Lzx62
lPhfWmMNr+3ZvEL3RZdu6KXtJm0vFRHO0kXA6qoEIJZq04+2qCb0Dzq9PGSC1l75TJ4MJ/oKtxGA
7Pdn1erzWiFkyc75nsMqwYY+QrHaO5tJjPQmguNxw1NyqonAUFjOwHojpzx0nM0n08KZ7MUGP/Io
8wt5xpjldEfetpYbr/p/w1C1LZD+wZ9CTVwWuB1oImXeltf2tVvmmZF/zS36N/kzVO5+tLZ3HqRe
MQCwBBJmqlhYA2zoaZV/HyNR8oeXdXXkX1YedsSe/VT5IA4VHGHk2vSaZz1qiFeR/unmHtBIFbfS
noI6HeEMU8tVGFICKkFda3L2F1bBVgeJlhKiVgfvY+xtr0jO3RtnBeG538FB1e/6XpIwkPVk+N/4
9UUZ6iBr8cZemV4NgBe0I+oFR/o5Xodg8+W42iFf7QaKhnhp9EMlXcRJKx9QWpZGDoplTXJ7svr+
/dbYgYNmau5divy2wi89gr/1SewoysI1FcIR3KV9NWjy5DuCDI45Olb46gmt1c1BzsnIvBwRyikN
5bCaJhhHYlKSsubJnVEQrBHcPcUoRymVZSToDJ0L1/4EACNQkWtaURS9Lu9O/X/Z8getBMT4/S/w
sNuXIVUJ8gC0GPW3EJuG3kKhRQXEGEDhpy4nhx6xrfjQ65dW6jGeEEkBesXOpabXtBiXP+nrqVd7
iyXFzM0XxgUCMdczev5qjUFfnv+KZtPhla/S5rtYLtAO2mw3RTtGGl9RagAsSrJBmKZA0/o/OcKv
5eLUi9z9L7zV/zqL/NtIm67KbgRHKU9tzY0Q6v/sPow28BVj1gUTM+xKMSvZKc2oKJzvGzLJhDI8
QKHGmeQS8tq//64mdJ6lhI//VVqx7SnDC0oLdsJs4Hj9ZPVYsM9I1aLVqUmtglAi6KRt+c0fWkR0
atmQ78hBqh90uGJR9cDzsyjv/9UdnfeZksTNEKzpJTVgpjxzJGCS1FtWTMsNs7bBrPKEND+aD8GM
ztSn1kDjGJXsPUPRHEGp1kJPnRA8tCEbyPxB7/MYDEFJb/MRSQJLYL3TV8b9eUYy2G/UjhQmTmyC
zKbp1ottcFKU2OJ67Qb3P1fQ2mU02s9pfKrYzvC7go/iXF/PuYw5+dgTyHqoJAnDNcjszSg3cvhK
uMsMrEYqYel+pXe9L3Uyi9nLZ5qBohap0pEK1m+J+1DcYFh06OJei9cSOoScmCurz8p/9eEIL72S
sAx/QjBAyLyGMMP0BRT4DQ8bH611yY2q2kK/3ABEdUcWr1qy4vTpRKo4eB7BEvXoej8Z3JL5Eo2i
0FfinKopqBxyOuiEidHMz2A0/VNlRlqRO9kcqpcCvzJ86PcMSnYsq9EzzuL1HWh71O0b/B5fCDfd
4HdBCGIzkvtMkf7KLFgntuVBKprDLF8oXpNh1PmA8/AN4VDpolbIMIZBZVl2nYWPhEp9qIAJjsG2
jkr7OHlHTVRyaie+BxdFkioCWHT4+DEvidiLBDG/A1hOMGM5jrWh3bWBk43cLxfOhFsQeHa78SJU
1OJuoBiR3IroH/QOCNTPp1pHRY7j8QxUV9JEOLW3w1M+EwMPCls1FzoD2Jgpl2GMSXhqlDBsM6zW
eUgiNCV9LiNfAWK3U+JbYeP0mbRmBd2B6C9B7EaROpwJrAxbDHjgZaH3iMSpmNw0dmy/zXACXTbH
EouhvFWj5mcI2WoztBAYsapDMBzWJpOyOR/sNTHIwNt4IWWr80hBRT/UkqFP8pzOaXAtiyJVE8BG
jVqBc5wI7psj3aoM8AggZ7XCLIYZ1vrfd+DwgN3hfosOUvOqsXrSbQBj1/Cipmd2EWiWGVwWjDSP
6V6kWHPNyNrA1Ow9AuhromxIU+LgxeaP4xufBHAzZYBp4Ca//wdF8arBYUULH4JXxxIbVPqZV8gk
wSnuU1laCN7S/TJCFtMKnJAd/lJPuL7CkVprDhJcUPP8W5mT2rmkVisT+AtB5bN7OnIPCfjClalb
l0c5rE96onZT/CAaDh2UD+jTzzpJJyHBc4r964WANilfV7UqZDkjp53P7exaGma/nrqH/GCjHPf3
s4FcecqOzBmJJUyXfHPADaAKyNggr3TitlQcu92YdulJT+FDR21g/BAb47RuHegGQVLrgbFX2JR/
dsQvyO5Xy+X/vv6/cUtRYiOJDy4IcbPan9yv+VVYdqHdQq+3uy1TyyUOA9nti5OzmKqCsAVv9Lnz
2lbUfdfUP1FeuHHkQE/q+1O+vgLnJQjnQ8sk2ir9tS+l/qx3aN1N9v40IK9NjoeARutsrBsHQ2sX
xHtqv7GgIxKhIGnfL6ZSTXi8HHnR44FxG9nKOYKK5QWBFcs+oevZVzTxgQdTiZwXP81Y7RQviTml
FjNzAEfGh0ceRe5byalxCbd7f3uTyhBHnO+Arcpd8DOy7Qx6Xgt0dnIo0W48iitjnQKDbrNXfTrJ
Ijgv4nR4xIoWNjz1Xe1SPBersK5RScxLQ+7zCgaKOehehuIzo+ecKa14fsgptKuDg6ZGWrM8l7r+
eF+kxhUmmraf/7Q3GjKOQ7+Gxf0r+qnYMvaAqJKBCZRELIPgZiO58htO1V8Vzm96PxTa3BPegF5j
kuBrIp6pUgBiXnM3QcJL+PwkDfdFv8y8HrkOLd2z8KhPk0XWLFEK7LuUwlGtJVzrz9aAVPbuVQRb
KnVj+1sE2lLpOYajABEfBFduTtH3tmJarcH/EEt6ffbpD5wLv8K1yz6mnjHqlEm81J1xwYz0QXBA
bqsPzJsKbf51N0sxBBkTW/nABpkx4n95eMGvwG6+/tUGWOqoGhfZieG6XJIbwu78chUimxTivRbK
/FOAzjWtJyPush7vCipbNB307uW8uDcMXxCqKxTof/cOPPPA+y28Yf2Ey7GoY1MjAJ6NPEy2CR6Q
RoFRIfnvnAwyIevJ3xtt147/deyP5DTuBVP69HcWL7VViv5gxbW2MDwKacOFKKW0RaR1OMZ339vL
xn4+1CslxWA2sgJa8CDqk6xUPeQD+KY5pGGC7y86rI2SJ15qgfGbW5fWVQQyjBOtcGvJ9/5eUqln
B1cSf7QSJuYIaoZE7Hirxag/wuYL8UMkvAuc+biublSuMEyQXnuyQ3vPFlVWsFz+2s7MjhpNbhmA
qHwCXj5EcOyXSrnTHCNF/+iZv33WtebW07mcpNv3T+gqtL1B29ZKQ06u9tqnV3w9thck7m2ojxup
/8PdekeHSENNWQexUV6Oem0r5FbPnf0Q/B6sdEk6ZKZKUgkdToZRCgDQo9+JtkIjD7Ysb3ZTPSdr
wVooBZB0LP0l2catw547gURybgnYwLFd0S+b34sMFvBoj/aENEqeLK0QHF6E7s9rJ8N2EGBGmyWs
tQ5hBqI0NUpFoEuUXLi/O9zBZEmkq3KeMN2vkqpzGtRHst9Q2YvWRIV9BEZZrC09O+2ff9e8jvmJ
cWpnhv1gu/LM8Q/skxyJGtGGKa66jaEkqx4eRyGHGzrv0uQTMnmofjtNbCALeV8Y4DMs/qQsm3Ia
QL2TIQ9EFZn9X4196vYPlbTy7749kXTJkPhfa4+jFOHeqtkXRpZLSha5PeprSjPPoNsNjpFt9XJA
HkaWg7RdzQklA1sM7wsnKId0El7/ysNXJmbLLC4S1F8tCGmN3ZgBnV9juPvP+qMmeJ1jCbrn1KxJ
dT58g/co17WhBDAQmNWhmiv+jtl881ZvmSNCIDaeh0QuRf9+rjD88MLHXdu8K/Ut+nfVbQbwHDCu
zMvPyk6v2DIbOJWKrFzurG67GEc4pWjPZd9f5VhVoIpsR6XBX41exMpNcgu1X14mDQZQpv0GLvq1
zcrOXGlZ6IC9HKBjDTMJKOzDAl2l5+b35emJuMjp6bbysgkXBvwXAl+aFAX9ulWRNVyf97UPf1TC
N2c5ZJWm2/oo5BgFxv7mkbYE/FzstGqL/45QLFlK41DEfcaI9D6gdC+Q9SBF2f6ije2xY/IYFjW8
Rf4gS/SUA+b7ATsNPIHpnKax/SQJfP3+uAA2hkys1iQpdXBaD1kFqER5/1vnGlcM2WE+NDUEuR99
DoGox/u3y7yzvNJVtH3efdEp+Hi/+yA1kj+DkiTHUsMtWgOwOKbf35MLpNyymx3ibYmGXd3QJsOe
+XxRuqcktqM9AUULY+zCVmlh7nVmDodlkgBEMKZp0/OeZn7gufqnwSeE33a1XaByhKRhwVCpOYGm
x5yDNr+zIq5pg0/Z9XrvuMkGYcTrSwS7YOLoSJjDT6+lhDuivKspQLH8tvNwTQlWlCSmzEYcIOSc
IKnjbrBJq3quhHdYJbqA94bBkTIre7ACFRmYtn9V++puv0Y3EAuSI5DNC5pzvg6jibJQG6TcRxs1
J/bji4zSmZVQnGDeXux/uR43oaLRCHXmGrdmNRoPPgBQn6ecYhuh+ljJiejtj8auMPNm9RN8SacA
ds4vlz962rIkc6OAFVwJiMHzlBmA2JIYBfQZC3JrZp3/wEsEMlkOR6Zdy8d6yrofjLlKFYwVi6B0
wdmu1pWrR1m0WuBBq0+jD1ZH8D17AfegGfsTKZSz1LHQiDI+WcAmmsudC4k4WbfZfqf4Yj1B7y7W
WdxOP+svPjSYtuLvz6ghuc8MredZx2cYC3ZVuNZsLSiwY2z5O6Uui8lZw1ZcxQIADJlKAyRqsLAY
m4dGNotkHrMPkiGhXx8fjbOR/LP1mwP463Hh/1EdIqn5el48R0R/8Dwl3nqxLsT+R/Zcq8s2P2MP
hyP8CazKEHjUt0cS8Q9PNfrTFpuIzQXDbFvLpxtwejyEKYOLGIzjFgXU3AqGU9IclIeIZ0n+po1k
jowWcMdRCnK4i/NptN2pvigqaSqFZHOrN45ysTTgjyJTnCzKUCnACJPYC/Rt/jvFZFN7EcKWjnOI
8hwbdKX943TaHv1TfA87typFpoYFkno01g19fZ2AuXTNQQwDN3hZEd4kuE6sGbPrs4rTRMx4kX8r
I9MfF9Z/DOV7m0FlBnC8vV4+pI6rIvuA5Qe9zJwdNMXl4GI5Kk3JAomRVFXq5W3c7PwxcWB67jZA
6wUIqSrsSAG0+rAOS5oUhaFLTLb4lEV9inrVC6G8FYnJbV0zGxoWPqaqjbA+XJnBNiR3nPMsozG9
1myRXC2XSkWD2RLdHAuoKOc2GaOHyvoVRSIy32MpokQ+akr+1zgMbVQgpRRPeJ1i1SH2weMP0rsR
KmufHzSfH7X22vMTCwYtjZL4bDut07VPdopc6qfq7R85Eym5reTjvGAEjY5UfKdt0nTnGLl4jNsy
Bxe8fvxae+lR655UEMbXrHAUrAECUy8lpsJw5lrn4tUWiwb0Lx53BreF7Rzv1qjv6DDJYyPUH45j
uoI5YUEEiLNhMjS7rQTb3PTQ4MILjcTCx4SnlwhXcEAGDyWK7nat+Ryc+Z7s/ZIjIWdBhBWbBcOR
/cFjB1D9VHzFEjXNq0Z5052c7exGSWeBLsmfL17KmnTIAFyIlkwWlEnz5LJxWWVp+2zwUuJr+AKL
AuiV7wELlA82yA7XbVYLpwvvz05yI8HxAb7IkVk1lq7I2Pbu21DRCK3by7fB4u5Ei6ku1rwPNgbu
WoJuegqSzsMaDXr/hCK3ISoE/5M3f5LzjEs86ElzR6EZ+kIARCdMEjC0EWFbTfQbHtakTQPR411r
ig6ah2KBn88odTkDsCC/lqX7Z7OGlenECcSqD/5PYKxOWpXo8JRVwzEi4JYMqBET5jtRa4UDTiep
pCBB/3kjvt1lir9B1BYPUXRE0nP1MNOCW+t+1BTKoyXWFQvHHACwq2T2Cn0j5V+CJ0IlQ2rsHxW9
eyhtqEBaGAeS7uv6KrTR2thgKxJiUT3gfRqhqDuWBMpWkeV/u94GScubwp0nRdo2GobHFSjbw5gd
fFr+4NYkhy5Dhds1gQ5Z2B5eGgrvxX1Z+Htt7ifDlo2CfIAWZcyXCk5yLHDT36B8dxs2As7YMS1L
EOKlt4q18kDbemRdXll2KFA3g+Tgd9aHH1TN4PYBCW7BGeChjgGzbSrAH+UFRb4Nq0YxRoJT4jfq
1DaUx2QMLNZeTVsARRX4jUS0vxeWUUOG89WOF54zSPCoQlObIInq9T8BZ1kYE/yoPNL7ysvHgByj
juphSs4xVv2JEGdEs582wMxR6i9Ym28akU/On63ebUtMZ47Q+TkOdBIinisY0HgJJwqImWUTAGUu
bv878+DA50Czu4TZCNyIqpVt/rAt8AB9wZ9nz9OnkltomeUk2/Avo63TsWCfpEwoqDsTa2B3Kcav
pxtHU8zfyqGbIFG6bi0qcuQqEJAyHJJy16fgGz10fEMkiyyEKWvjn/lmvQUR0uW/nFHq3N/48Rbv
0SX9wmauXFGB03rS9OA8nT19IeBevI1HVqJRcxCop//dObceX2oY6stAy9XS5tIHFq8bbd4o0UX0
PEwlmRU/U1rGDdBzImaY3Fq/q1zeM3URhSTlTdehtxtwGG4mVLDyqYeY+4nGVI7u5IzZ4+jB8Vpk
EScLdSBJ262m77DSLNrK5LLawG6qVkToh7wi6HD3CX2VBYOm1D0uWBLTZbDOGAJm+WSmBN9rFs11
wqX4FLfCUoVstO99o18hmpMBwLDvp2u8A2GPMGteYPLUXAPCiw8vH7YpsfH44UUTPhH+0HcGg9cg
JwhRN9OXfgWyJl05cBmVRN4k37H2z4hJwp/wj/sCqIEG7BZzCYzG0JGwJYFZaz/SREls1rlbOh1Z
lHHPTYNWKFWeEVZrAIPS/pou1jlH6Z6TWQttGns320fE4VBQa91Hdu0Ll0+n8aTd/BpS7/sTemNB
Ew1QxkW4vZYCNJ5MVpbG1+Rd4n5mDvMykBxmPZccUBhf6d7RP65NX847tC3RkOSWjb8jILHigr7e
pkrHeTP3bS6MOWCeLqXW6qMmOHscEKsENgfy0zBD9gcPTI5L2BzHZz/W/1HgLsdN/mS5OtVIbkUh
Slwt2iXRpIVxGQ3tN5twYLF38QgTgJ3S7lwZ9Oopu+roz4RJfqT/6lDH78OwMRD+JhrZV+czIzpT
hGaXuPlit6Z4C/xeGunUdjd7Z0ifDsL1Q7IBOgcvxF5pp4/bDQBJzu6zBuX1sbLpAfTRhs9wQjBP
FKDaFbq9wqmJ3CAKZ+++E0xhQUAZcegReTzFKkuEWNpNygMxwQyagtD8dTzXyBBh9ZmfpLp1julC
2lcakytgbBSY3HFCgqdfEBOT6mx3tZO1D9Wz91CJkeglSIqdnMAbO7fC36Ca65KLQkXccIx3VbU1
Nk/MZcE7Rb/Te6E5OmKRzQ18LIa7VmM+NPh9y/MZ3P6DUQ2rFozgXwYbF62IzqPgRmRGIo/NyGBC
NSY8Sp5Dg8hcsWAiix/52+PMzErrkuP8gJ5NHYbhFrDt6b61RVufy720Mh+EGfV43euUcUaCtEiR
ZIMSZiAsnz0WYz5JElTlrCqvJ4mPBwOKKmMRVBWm/Ey5vf1wUC8TFOihjfmFmlfqLpFgTmVwm6pV
d+GKCZDmKRcS1jHbgCO99czjUzvHv8gm19cEBC0bTZckz9teBo5dlAsoaAgANsuqLZ4wGG/BnbZn
dsHXC3FSPERW208rSR1P++80pMPgNHruxxB4q+mxdZe5dzSyWNcqWFOmyxJ0z+2TnimCW14BDdT0
6dl8XcBDaN1kmBSXyk2VIstw+ya7rxSJnfrg42YPT5K/nM6aurrTKU3qzXfrYCmQ3886hcaTZ8ba
WmGgPZ62AOw3BAQHAvK3ydBJXb5+yqx2HKtWBvdALqUQxWzsTIZlMnlOD75pGcNrG8rVqnw8Q34U
O/yhDI6UwKoLo/7gzbcq4FYiQGF0rMgseCzGkjqTH+hrxOHIjKX6K8Pfl+48TyNDlXzHZ99QGrlY
pu6W19QpSPhZLh7don0gjbnUeoLx6WG16904yr6jscE8bJzTHo31O1Ew0SEfpLKoxyOIBGi+ciaw
nNTPm7KJBY7Ekloq37M8T0WHLAo21aHmW/IxHcrUSLHj+Psi0VzURNN7d/YrCIGXjlGohWZZGt4v
UPrFHI9AY/ZJanBsQ9l2k3uV4cpX6erkW1rL/VvGIfy3AUAIbY4Rp0C+XIdYcG/GPikz4IFk9H7E
mqoz9CTYA0PQ+tBDinPEn5somYF/sABHaYXcl+FIdG/zNbhHsNVPJeqV7h/V1t/Do8rlIT3nEYgM
MM1W/j+aiezXd4xxqBGc9bvGxLmTcxdYbbCyRQexvL1CYdSWXb2eoQSY/4NMyX+Zf6OVd1Xgbe5o
uXmaO212AouXwh0h0hLiuQBF7v4CWVWUpQp1ioo9HfsEzOjA6J3f16F8sath+0VJyOxhVsIdIEhi
dEFSN42jJxW4a3F9nnpjdMfoesi5PLtPzCJVazkcG6hiLYKvn+qNsiJaGHtkEuBxDt31w+/S2YSw
SORQgqwLSvIk040KsagAbnAnYGJ5j6sIb3tLThXiV1M/BVNa2TeVIQDlPip5nEjpMqVXNgtwQWi0
/kkBHves/+VTdjqBIrw3fL+XLVpB/E17xXKXTftymVbFzQ6Ghk+iz/+J50ttwk+jNX9/vm8PMaqi
0Miv6na309L+hOtnPGv+v0pzYSDjUzT5vLZPuOZAI6ibAgpSDC0Sz8ZHMuVm6E19OjXmIt+MRKRv
yNlvWwKkZrlDDBaiYhWazv9O1eRiqbURSr0eOcyVhkdvbph9tLMj/qOgB5uGiyRNebU+REaCFrPt
JpoXdVM6jgnZBiAeTwaHBve9aWlLo92dDYQ4Uz9I/DQ3M5sS99m1D4Xsctkn+CUzr7CrPmlZL+mO
eMO7AaXGLJKpa+QDVlyxo2TnyoMJhI/CKwk4LW4C0jILqioyOEYxIG08RUm9vjbvTzkTOq6ERPsE
0ZWtmhzB+WNPyFY6FTT/Q9l1HxmuC8HzUSPMHurn6D5Q8pkOMrNL4vKdo5p0cormsuVMQ43lwpJX
WeRZzGS66p0JF8jx258emBMvQMGzO40KGtjHTicOVcUkSQ62Ea9c5shTwdrBGnqoOPpE62ZVlTAx
ybR4RqlUZLl72Gy7FRM1h9OFhuDvg4bVVXjT9YDhwgq4c4vDpk3x3cnRmoY6UiKOXNa5vVMC0GuP
LhMxlBmS/6plim6NxyEhsLr64ZsI1ntelrSCPFA11u/Ac1d0Z2JvfFX5AwkqFDjqAAIRcV74CmNS
gJI1Ve58DOT4CHXRYeYJJXMIHbT6/QnCZCTCuEN13R4t5qh0POxnI6+2vXo/RgSE5PpaSAw6H2pT
5vg0IM0ASumjxQxUI4Vf87m70Bm0WWEK5yq96DWRUPZjJaFU9VjUAsuh9a2Ft72053WR5hcHO7a7
xUibL+CcgY9rfhYHKkUVrXTwTg3Js63yPOj+EohVj0gzVoJmCxcPfVm/KIfSSSNwPMNeqkGwSh84
iLRvAKPYsirX/kDNkuzWilNYfWO8hFk0iAwcRTkihTNRik3VIgIoC+xQfBNEyaZ/KHwcS00U0ya0
xbXtujUp2/bmXReUQcY7Xu99ITozyZte6lYi6bdZgg8EQkEjTulcenJiOn/CoBgwcs3Ob+48gtVv
oLjZQ5E3NlWxvOwXDFxzTg45RIn0wWL5QM1dmNNYqWKqtl9A1RzmzVVQoZ96NZ+84N6Jv5xOU+HL
onUJZI+f+UYDIZxYRmSk0rGJMD4qKVOZsgpSZTBUn1GKz4dwsRGcGlIC0bJTchALd3jPGUVX1Gib
RlEhUQRs8nrRVQL3DHxKOlbZQdwemPLB3woPIIbH09hfLSaSfOJln9Ik8ek29egE8rKsr/OW/mi8
kaSJJuZKErUmLfmCvrxxFtezdImmyDftikErMrSrt5hNEJmlGzjHj5IEqTl7WU89zTaGC70JQc8w
GDnsa4wNNmLzv7a2wTeI1DAKn2swaO0nANMEfXf6AkzZzREW4dWOuWVa986pBQ35kEaXCgff2CFD
6lI6/MKkU7zH/Fc4qTTU54UqXpt7BrKAMhksPeg767qbaVN3cLywrJbgyp1DMwaSDd2ZAmWfn4AR
K3Knv3Jyn2jVyaubByz53LX4GxrEZHo1uCH4i6CFzOapG793Vuati9gh14dD16Va0xzMJU/XXpso
4X5a61TH5B29M+l6Nd9kdjRLBp6WmTfVOetaVajuC652yQlz/78xmMOA96PYb3JKK+Xk9iUafoi5
AsVT4lUQW6WR2dUhWOQl2vmYsJnaWJqybxxwsgiJ8VYIOc7uiowApDI6znkpodR4TMhGRXHsRmzB
sPEHvr03NucT5U994n4NJ0la1k/XEorI/WOvTibtnsJakpfvyRZccHW5ZDYEI/PAEp+/JbSUEx16
LCYNBWxaDlikmsr8JlM+CdZUggD0U53l3I6ZDu96vYYOCGV7I4GUaIf+SOw2DkGPKH4ocq9CM2yG
cC1L0AtFA7ZtaHXG5TpQhM9JVan6UKlDNXsEIMgX2kRp7eOaY6iWn6CsTR/MksBOtDTR4v6Y17Xe
L2Ij5B1tDhfyFlLRHHSuf3uMpw/L3URt9r09NGji5AjkS/ZUwEWYcF21svcuzhru3NkkW92qY/xs
1/3CO9Lfr4uFU7OCUYGAL1+WRmFno2TeDM3+W5ORF74Gee14+l7TFvshi/3v40Uv9Uj/Z4GsqEBj
A9cwXfSLqCYomGis3prhL1VdRTmMv5VwbFseLyqzIkP4b04kyT2C3+J8+N3ZW0exvjbm5hzu1BJZ
CIwuK9Nd7mpboqxhUwsYag97lUY2A4RK9rjR/jlj+Sl8bhQNxL96aTmkXSC1eT3pwqxUWXOVzzlI
WeR69QBGZyUtki6fSWIPU/aHCdzV5o187c3gCS5SvmggWXPtywI6bm2A6DbR887knWk7r6pQa9Z8
3c4o0Q62DttxG7ekUPunVhJ+oioxqwFxzhPCQCEK4RoppvRsKLUfwCHT3Ux1I0ZgeYsuIvCg55WG
4t8TtDZyDrKseGyp38S8n1Dj3xceMbIGi67FCfM0tIQOteUn4XSiC/M1Er1hv484AmbxA4Qv1oM1
7P6t9HuqqMfXhWufl6gqYAJEvsFlgiBYo0Ki43KwEt6Ztn+4zzZz2m9dsgNRqmFrC5IGp01R1Gl2
sYHFaW3mYjgeVgiBwUoajqxC+7VGAZ7820FwxT47tGodDssii1BqtqZvD5EdmJcYi1RU5lSjSeLQ
3V0k3hBiLwXxyrNjm+44U5YvMkUbMNMbLTxk4S8I8qTfgvkEOZBibHkz5ShQZATR0QoMhS7J8wGQ
iGtbArOCL2/+CX3Y5kfeV/2fYHQkzSrxzbqKOWZm+Z3YWInUeMKxnR5w6Tjsf+QkGeTu6bGKDW8V
ez6iT17s4HgQ/oszTX4WH6GgUv75aC6TJ1d8/dA8DKjIXrTRsksp7BMhS/RVz06Rat0YLq1rO8x9
wH0HHvyiG/mwVXO7c/HQNYXNDAIOdsxJY08HeA111RzQwzQ1Y795qJAPfXkBhl5arq6BztH6AYcz
IvXhN9pA5u3kNjJ5AhFGH8A78lZFLdiQz8Uf0HZ4Cl2Z+70B4a9v2Q+7JOQqtuVpxDIJnN3E9jy9
X51mrK6NeopQ676tKwDTpWnxFEVb4eviOLXqarHpu+6JnPxV63uW+/DktosPSgnUxams1VjWjd60
gz8JSvvd/Ul8FWsUvxek5iQvXZQsbhsMWshXj0Y4LOP75HYIy9wZp4IPuJZQUSUa8z7+x5UkNjcP
ZTGCBb7zIJz+rMTJOhRCJKC9WiAEweiVJ+8ApuACsyPtlWmwdZ477lbmxolRLJNACPIqcqqpqMC0
84gddQexWbTzc/9WtcsE+kDJ5Hpu2YWLwPuMLHieT6S0YQjxnYczJtIx9h8gm3nzy8L+MwMnrULw
NRaH/QAZoGmly9bIEbjyZLnqDYQ0gxj2Vqv1CNZO++ZTkDS7xavs58crZG2jtlpr4F9WoFpOP2DR
FCAjnkGJidDLI3GqsPalxYABimLXv0Axn1Agl2nk/NmqFxP6jAb0USxu5Ng5dvdlkD1zwPqaxbKJ
rsRlVx0xNTyfZwq7rvcFRVuD96dx4PVkHX3dMQd3CaVfbgActjrJp7xhBHrFnr+3gIu6AV/O5tQW
aCAxS3QSPOdihrtonXTyvTNO7VLfjfpjy3FmTGqoYb9dtzsMhpZE1TiYvhCebpf91U8HrztMxrAg
8XK/6EgnRnmQTuiewG22bj1gpV57yE/aCLG/UD/mNEoWKjJOvumnmJCDvQP/3jiAEfsZ52yq7pqL
xduvYxKdUwNm0U0f0VzXW3BPWUckTX74tsjqGyaL1r2Y5oF+I7N8gvd2hF08m+oLm4Sbs77wS0p8
MIq9Aaw/lHfe9ahVrof/dcicrY+uSVM6N6oBCnNvLvXAkOFPRgG5HGqC46VWxs+elPJGdbypcDLX
MAycSPPJgAtztnBPwuM+56LiVH4z5FIkXwMrqPxm8O0qDKlDCXshtgfP195Cu2WlX93Rkmm6jMXR
w87M6de/m6EGVJtHK5anuiK0RCOD6gkp3c/q2x6VBGOOHIDG7fBrajmYFgBqqka41rOQZibe9KQ0
s1N/ENPgr33jMDePk3ouJxxTyeysfK1m0OJ0d7uiBm0DOm9eoRmXoiN9gakw3zSH4kRnm44I3e6K
tiQtcqq0dS9kTzdSFOy5xYzjqoADA7OoLzlt18r/LSznXbwovGub6egpHEXeG+Hev99X2Gwx21OK
Mt1IsDXh/ok/7iOYu0NPvosleHgJH1B4n8YIAKJfRAvTz5WbD+l7NDxNeRYXOQpUsujNIaV35YjQ
qGYolhI3N28PBDrl1fqGYqqPWAToMFPo13uawEuQ9wApf8wcEQ9Dx5SS/Ho0U6FfgdKDrNz9iHrC
4qPLWn7a4/Q4pmMsd2I2kBp9iQMygIWj8dty20dHG6NVFLA6bk0dWssZXkK2NCkaaEjQzR3rMMgm
zjGLWN4SThqKwgaOKPvED0TnN6gSfaRJjKuMtKLh1qbYxavQoAsUMz/A0rDYVPnF58BTt61jAJ6q
7sSSTe4baLxqI9qUD4YaDv+F5PdQnMe9rHQRES5ip7EgpMEeCJc8UfsCCH8SxUSaesKqYhaSwC4D
c0kVo1od42SPotpanTDFc7di6gPgLPSLIMk4xYlzkBtmcfsRmjr3vkBcA9Jql4h/lZFnXvorbRYR
pHzSfl/Oy05Q8fOGimf55H0GeCE/fbR29ZgL/20BwqgN9I2SVEwLyKJ7jmcWwfUM0KsbfGe8+jOK
gn+oShaoFODThdcBhhoTKl+qephx29dlF3zIL0qDDDUVJhneiclgXOGuiNTawPfHThnC9UFbRxrt
GgADiXfFppv+GKasgIkfHO4J3oih07Lh9wxOF8KZL6XtkqpZKTRSSrElviA50Dw8mPKrdjI4gKU0
X/RZsWQuJwog6BK8w9E7eNtMiNRZczPPBhlGj7g9XFS+rjV6z6iI+MB6ek1CeLTHpr/GmG50tT/L
rwFwlipE/oSC/PnF/YynA8iBvpoLJRz075f3H4RYiSuS3Dg53rX8Fpr4W+l1nzVI6p7miM9K1MZS
KeVzq5o4SPONuYfNOxqAnwuhnqxotbdpxLrMyUaCNM1tAtg1rqG8OC2EpMFOMQ3as2UbzHd+byaa
B5Zbb+AtAK3hVogRbZ3wIiHxNPse+9CeJhNfXB3mLs+sW/ygjI3UJKHfsLmkKYjYYCDiM+DQC/CS
l+wQyRPT8bASnqtCyDzwifUJs+S2KEUfNVGH5/gstKPhxcV8GLFjrgE93FopVJDQHJIScUnUGu2r
hFN6RR+T13Q1hDsarBvT6b083Km+9CBh0cB/P8yOY/E98qMyPWPe20/0nTfEiI9V09E8KQjB36o/
J3zRr4eibo50VLv3fjkNPwr3hVLYuQBZqj55wKzXJQL53saDZ+hsgxQ7fae04mYndKaLefKf9pxW
IoLO5FA+o9LZmibOfu9hq47BnDpus83woYT4G6qpDjmb84x/2dvr+1OQpkOL3AQP6WSMt07qICso
8izEmmR5M4gSxmOW/7aPDAZyzamAN1KgXGxOdNH8diaeVzZf6ogJriy3KN6f2ZZCnqIr1qrKFo8i
yheH4UJyIeA0u2AEKMl17egvaXVzn50keMw/+eQqhMeaYC8I43dEf0cgtmbUxf4imWqkmh5Upy8T
vGyYXM3sf/CRBUKjtAkaLl8GB9g8A3ClMkv5jgniC71ISEqfsKYBiImDA5WQQsGM3A0J0x7r/9Wq
dKJWGmG1Y/BM3VpEjmjY8+K+TTFFuuvJ21k9XfnodW/lw40d//P68AJWZFCVWHyC+1l+4CHGTUFC
LHO4x9p4lCnpwioK6JvCThJwl5ut4EKs9VFT2t6hBJT5QBlfmIg/m7oO/4e+m2Jsi8tC37LYFtuG
Ha1fMcZW1vctoKJrSnYuKL5EY9TQ1pCAO4gFRm6wnqgqNJi67lfUxbuZuL+Xitf10AI4qN6U5RXj
gftPhXGnFeIQO/ERMJgRcBJUsCxNQCSAkTP6h+keGama2aJ6vVxFskNXRmG+LinfZU51cZueRUvF
gf3/Fd8aF9Uozk2WhJTgM7HFj35HFuWbjtTrnX4EGLgFJZHRQfc6COcqnQD/+m8f/CVQ95HV7XD2
nMN3RXKg/vXRF0BYzUftPoKmxA1OsujlXZj71LM0sEUeXWZZS7j64VAY+uslzHgANO0S3iLXiKO0
MhlNNYkgBGuXy0bC6uG7BhUS+FDbT43p0cx0WJjfGUATvs3Ypw1OGmm/KkB2jQ3YNyEY+vE+2YnY
x1FiQqc4Bm3Su2Q9CKA3ra10Q1WgNnyJG1veZdr/gGLkC1JWWpAZilzfImh5xAbHdDxKYWMD0BXd
my6FTukOCN+jgTcHexMpDoQVZvsnVAZZsmoNW7flGMiYOqANFlUYBYDirEJqk1S0V+dJD5lUCPlF
olj6aoytZ9j8iDIlS5uXL1dV+6HyG8CnMuB4EmJd3Zq69qPGUmMEi2HBH0uARUKEALIPZondqlOG
kG7Pmqgdc7V+0fbfqRORJ3yT9UDsAWr0/GGuV/e/jz5cTDNvljXA75Buwxb7gDI0vjjduIMn5j+k
B/yBM2GtBLTc5wMaUPhob3+qkgFPx5tL/Vb8ZRHNJgmHN1xmgle7nFFejGgwdvMAvL2+uagGeeqv
MWKWsRs53e866bnqxpiEWxmXqIg7G1v9apXi5BfA6noIYocpVG4ildBK4M2wBOfZqYJW71IVVP4x
WOs85OAeBOaeWfUtvgs+7NoY/v5hK013jlWSVen47HDZ8N92OfuqvqokFm+thl2aTPdb4Tgnj8vN
+MFXjabYb0uQb//DQnsuAAxmh6n+VW3htlpiJCBuGvaxXYBndZ3ZWM7Q21RS2p33wyCPc98h0dv3
ynwfmk9bBxoug3IC3AJzPUmxArAfNLSs49IUSNMy0d4k5H3v1gqNaGn2AWDe1zUTaL2nvPwJx5bB
llR/AJRcXSBs3ypGMZiks7kkwZGGs9//SHm+6CT7J0xAGv2K05Wf2WUN7R/1ld22lZcPg8Tnsipi
1QcbKwnmpEs3wg46CyzH9AjRWVIwpdNqM14QkBuOtkFj729hx2wBmmDBpjde375OdqPDQkKHQG+n
B+l8hcq6F/VbcT+fcPcxI2N8BbqOm0cByz1wijwXG0B4gFtn3VMCpVf4GQMzVUWOct/nzZGRcNkF
6i/uRH9UCf5PNUvOki7xH2YdwVgLG4ezYxUAik5VpMpTuTz7XsjBDfCHga4sExqeDEaNMr8P6gb0
EUQfT2/NOh3NfxnUVHulOeeWRHOOeJXz7Jr3IVXiGIIpaA+zscnjHC25BOnJlh5JLh2619Fco3sg
rM46pyHdUd8pw8pwVx77SszDYcHg7wpzVvg4+I8YHw1ESSRj2krXi/VPKsvPQnnUgUyFSgYUc16b
FkiavE7RIP0LoSTcQCDyozMAtmpXxo5FlY7YuJ2iBrviIxjIQwB/50pyKb8g5qMLIqqIxebWtA6b
n5Fm3KNKZgfvXi+MS0nbew8B1Ev9sScLFaKBLCa3HcPSgJluwrpv1xSBEvmbuZcEGsyMg+8lNTKz
r6IQyb73Niu+z3RYAtdl5jIEOP5OvIMOAqBtJWHzTkeZKjsZc6RYkNEWijrrYLD1h5ASGvv6uQ+W
DUP3xhN8TIeQ07BKHlELJi3odSRrdOR51p7/QgDxkyISi84YMqVnVgMpYYDzG8k8iux5Qf1HZI6w
e4MSmx9V66kAym4/Dsien4s/wru7Zp42dUxPGQw0fWQxxtlheb390nDm+n34yP/XV4gfbEc4uosw
Pc4uX1WiCxCErT3dZNgN5fwlhXehhxqKhf2QIxpseExC7Xqudwek+A7QO1IqkIQD5K8o0ctQHn3m
BnzkZxmIcZT6A4fq3mFxJMbaEpb5oh+P8tDSVTyx25ow1iBxryS5ZxiH0M4uHPjoEug813My46fz
2lCNxXkIOjy4cz96vR+8Ht9HKDjQdwTOMNrbxMXXt9ZEpS+hfocOWQUOVt+3Zg99jjbUqnVYSXP9
42rGSeZdpt3rcusG3bqPCLjMEta1WvWCPY6OKGjD3GmRL3TPAX1qblGmsyGjTxlRrHMh5Hm4OWoi
2YFRG3UPp0lv8HOIFrhHRIOVet4/aKlWBFn7hUGEBfq4U+R07uI4ui+L/p+fPCkenyW5E3tHDvaN
4HkEEWFql1XWBM3f20b2lBy9DX4rrGbQR5hLyqZEd+1vyXASx311SLwoe4vtk/gXSH5MBXzo0qqV
2mFFbzJaleW+XtMGyb9sVhEwM0NtVYnyV36rX3bMOZt2kLqdRo5w7NRUw6XAmyq2k08beHQU62PE
AybEnukVyawhOCy5XufHwDlZmaeN3Z1DIov57JG0xPk4RfXXXMCK4K2XunveUEKRap25zpkQuIhH
cA7T8t9Tc2CZaD+Luf1Qobzzovr7rnfnqFQEVC7y45pNeRElpGHoz99eGZuOg8rIPVRKYZi6Ijuq
ju/TOnkNrgmQPXi+25ssgCOJLVI8+2ZmRzDwVp14QWdIhTcxsb4xik6gsYgCyJOeWqf3Q8zoRomR
Z0SEN6tFUB5P87jfoYv1eo66X7t18WwgKdw0ZIv72StAFHtoAMwhfnu4DF9qReYvST890AOgURsh
8hypfKBB7GeVjP2EFJNIxXzQkfi0v8HmhXhlrRxeV6+Oob/KZ2Z8jn8zTBKpAFul4XxL5HCDSHqh
qYGkFOe0wplpgN8JoKXS7xzmFiaJSOv7VFej7H92bUS2m+jsiJ2mBw/9+w+CIxOfMVzfI0pfHTt3
mZOGDlwgZ2nOJj7rFgSc/mqWfsk2PFuXIDej0wTFmh9jLHZn70FBsXIuvuwSFrPBY1ruE0iapNy4
kC/NtKoa9sHtDVgIw2hETo40cViRfeec6ZfFJw+42B2avf5i80LhjX1/VQB7WceyB+x0lWSkA4/d
zLg8biK9fExONDapmaUB+hQ7IH/LsyRkYaQF0ea8GSVpICCjOb2HxcvO6WY7t9RlKElt/5lTT+MN
vMyZtZ9V5FTXXLhq+41fI3kQAUcMqtTuh0iMKtlQLI+HV5cvXZWtu3A/Re4MQsfmL32RlLD9ODkt
dERM+gmwTkSiLH6AG6YvSvGdEHZ5jt7yGXSQ8dgTMMG1S+zDj9pSHHCFg1/tmx/oajj5vR9Am5jt
ZzzNTh5Bv9nU01aKSi9n1t956VB+MWWgyo9HkY0yMS7tZzfBMGZ+39SpsthXewQxZGoOXyBGz4ZN
+Ptdtg2OEHCauwjQxR+/PjvfdF8P+auEYeFcZfa3MwRSIYgl1W2t7A6++EQ/yW+D+32jolJBH9pN
PYlmMqX/Jr+P6jhg2UNGHubFkTMrnaK4h83CKwHsfBqsmv6r10NS/ZauOFvZLYkbWhWk65IF6nYG
pA7d+lUqSLUM5xJW8XSp6N05S6M/OyDo1zaMLSyg8nu9TY5vWLl7RWNJZsVLHQDOqjn70c8yBZ+K
mXEbeNP/oAQl9cLo1BTlFmtwDzZ6PBbhuqcgjT1Dq2F0nPG1TnxV80cYAkGxIOMBX+96hBFsWMer
O1Lzn/WYy715eRdDmkb8J/TN4Z3SaohvNz7tIaCRSCrO3a61apfYCMQqvCgEiNR05Q5jCwicj8/M
gv0+4txuA1JMK8Ao24Z4DLg4maPg5gqROq3XWE5EHNGYlmZ7JErmXwW/qNnsoO9eznxi1GdbnZX4
ebS2u7Z4pc88svl6BY6gavrbTOrn3DSRu8sYg3NKAxs9OeHp6vL1VXy36VhLg4gEOGjvjVyR2g50
593CQ6WzVKHS45skzownVa/wuJAZysaAfnJxxAKZMInDNk9KbvMhXOJg20dFADKLo0FHXv5IDv3q
GuT4Ju603lJoPt9LoGtmofbIjSAMPeQB7rYrtFwwvgK7Kjtw2XEnchf9mSqYuxBFoWWL7n6gm6fA
8e8Ey6kTy9ORS/5r0wQi1f6Z0z4PKfFY8jazXXsUfcXfPiFyG7uYAar9wm8lTAJ17YsGplhm+GNg
KQheIwzwRTEoxO+70EZoqnRytZNlPibP/r0rF4e0UhV0fHgTpegU71qbLjXMZoo6rgBwOW3lK3DT
r9CRBilARNkwg/JwV/ssTQpVUSoHvPSC2yJUEptCnL6bPOQjQj6MQpPDGZlnxCX2jtkyF2eMne7F
vRbBJF2ryqfeZ4J2f2PERU9cuwhUDprKGFnguna1NicJri7DSuAG1EHqbP19K+lYbNMqtsudWO8g
OMFevClBaTAn86CbVNAnIj1F1F7Gt1r/qU6d7Cg1CUajBZOpd03TxYPIfJlbh+nvDC7WGLbZE9dA
KN4r0yEaBsBvIWR6sn5he9tvAaGZ6YiV/v5zTT7h4qEhV198fW1RpQ8rqGI+NvSyt0Tzov0l9+iu
iN9PmQovxf40u2x0ZzjHZ7zt0y0VHSoq5vvYUfXlmJcx40t1REzg77go4LuI1RIIIdQ0PYWBX97D
qDdD6/vsExRcbusvqF1g9kdLMNIYzN1AHEUeE1C7mtBcMGkwl+tapjEZBdwpMOtxhTRm6xl+RNaA
aOdImpLPh1j/pgqPWBPtKciu07AHeexYdolUF9iDBXHctWdZcMeCktcMGlVz6qjOj4HfgIC11Kv5
dcZBh6d97uoVkVPtvcr4mDFRg5whLA2DROLedh/kVZjsNYxkeWcIQpbOU76Zdm9sr1BIzyRFNYVO
Ff/zKF//PbwZfi3rFFMDi4GdfzP6pjRVhgB85z/H7B7NPD/SRCrc8H1qAR16aDhwRMR9V30KnaH1
JMf2iBnLaeWEC7/xOTUeSXQIx9uuS/EpJ/rSwRfGVJ8EEx0fBknYqcHO3Lv5kLvJX613RS8NrEhr
v15fBM5KRogrCfbAVV52fPKUCrVMEYkz6G8Cu90jlPCS3Le16NqJJFjDrO+iNiBVYBtOyE/C2y83
/0ez8o+HNZVRwj3ZV0uT9OPtzAYOxaj5Mhg4oOvMxcMOY3d6mZ1dSJiIcNRj99TJj/SJPPqep0RQ
7kQpoAB57ePfEz7Jj5RZ2q6fEMeR7b1jn3JJ+xkb24vdD3mhrsgxZ49g+erCuD5Dxc9Ds+UrpSuu
NsqEZi9yhjISCjjya7c67Hs+fmcztvf/xcWV3DwXP7nSjB2MVRalfqcjNZHZZJqkJ/Dcldfp5oDM
HS5JlbpjhkKucv4rDsbQNvV1Ds18JUCB44tNmR+PJ5BO00tvCmMkEsg05GzAIluYsmcXf7BoZbwD
L0RVGWaG3PW+PlbpjzMvGVPjkcomwqZReKZrfBH8vzWZQzcg8GkWcRPrxLVHKtuhEnNGrkmqFN2O
ItCzeMB7lnWz/Lknr4/0wlyHsYlWzQBNPNNuuwMMTY6n7jklirHFUFupGc60W+uParZcOksAxIig
xgKyOpVKhI/+CvSeTTyZ+58YtFojsG5/8P/bw4RV09ZCNZcxlMjWaS9PK3Fc9tbI9jUAJ/X6h4pX
eCqUHmvHbGRwyutl8eXTbJzbQ8N7Y0WQENrohqPwPwJju1xLTFn6a77946q0v9qKxFYsMHGy6/az
kEThupRbew5FXiy/mUkOI8d5wuR9H5TLZbpOYbcvr8c+ofo9d8q0mfDOmvtEVFCoCJ3STujJxz08
EVSu8U3dI3jqgenl4mVsqoqlIU0gtJvCBA9Vx+P30Ud8Zp11upeqjFHgC3rEuwvJNW39//IRYSmq
smUmz+TSC7K/V0KzRhJ0ykGiLwKTOZjZgajulTfCM3tCD7KCN413K11ULrRCbFxzfGOE6dUUWMQj
ujwWz5mSAax2olX4JsmWLJ53y9ET2PGxfcmABFYs0tHWtlSRsU3M57ULblz5CxEXESNmfgpCMgEL
uWbG1wSbg6Dc8FIm7HTKmj+l8nnHvxSTncAkz5TF1mFTQ83smddQIHV+e+GfTMMaeryZznzVkxJN
mXfW+LTlasU1bqHEEqapcghFEC8nlxnV7/oRyhOediQeWDaTRwKO3o3jmVi3oqOJrSEdureFv42U
rzurdClTQ2WK1NscOi791Q9KIXpTtD9mhml1DP+2w6uhwePra/Kd+lYdKUZiPCbfVoYKlJPIrZ4m
KF9NY6nQD1aXKye4l3f1ROEPsrBeQ4NJGXE4d7eUuqXbbTm2z2OShhvukkkJw55z8buSMXtSj2V+
gITFw3D8+Ce31KQPukw+yR674NrhpqFasIaYjjPDDvjVVaSvSFRVmJg3dgGCKYyWJQCKpBhpCQKL
fiJQfr/kNIgVHwXByCf9DEDQom2GpHCbdo3iYDAi9PboGDCzMwiVc+89xjB1REbYydwLGjfqwX6w
HBASly9BdH1npo0cL0xtogVVSrN3m3/vNNitzYLeaRrBzlQ0dLojl51E1h8CIYRqwedR+7cf3BGq
cLuteYFnvAyS6p2IAs1OcQHpsZ73NtjGDEI+IE0oh3kXhj6KGqj4i+6lowjx4BIAY5w1CWd4kyt3
J8RECrzm0E/kiHV5Nh9r74XUk1xx7cDD1GtGlNsR+99G+2ukqiBvCZ2PKp7k+b6N/wH6tF+hMZo4
bWvTN7eKj19qoeJLLv5BhyMpyUSxslfq/y47DAzHy1CMZ3pOa93hF7mp9weqTNrHP0B+tAX1IMth
T5aSJga2RGA5CnuX8jeSKTQi2umwyAy78GeyUbJNwAffeQGeNNTaUFsaNAyJQGaqbshe1T2bNX3Q
sC16M9B5FF1rhq4Ad0A6FeVaUbGmMr1uSNbm7juzKOco8X6Ni3PeozhRILvG9FmPQV19KeSgH8YL
j0VCLlgaSwdlHbHIG11WN/JWjIh/S2z50/5A9OQ+aBnuUVVrzZ0cf7tcNqaW0YrOAOQbiMvxKDFn
NaEO91DkM8MQBeE9V3aETPmlbBEBqq0NoMbQX4300twNwpMfNU9uCI+E/uX9CDGlPg3uMjGZBCW3
ouR1kliSv/BxdskbSJtAvNXVbdJv0POO95Zk3vc2I9lSMP5fjTMV9+dAOm6JOeT4fqvU5Gzm1W8j
K5K1xXD6GNocVGJT4vC9zEc43cpaKY/WCGgfZlmkVXrUB/MiR8mu46lJ1DTEV6SpVrsnxrDBUYQV
r4OzKdzmnnohKWNc9l8viqWu+EgKeGHi8uxAo/DOLimPeGCrVVX1I8jZinrWn0iVIoH7CKTXfI3G
lxgZCV2TbLh3s1miuyraZOvBA6m1TceyIs1rirY4JSAO5N09hPhRJfxVepy5glRJ3ZWKzhrob22E
trBmoAv+cbDE3Pj5n8QD9pG1EfI8Zq3RXb5v1RQ8fZVkLNh4jKZAa8iTtpSWqxV/ETGZQfH6wNv1
ESxyMwnLmULOE49/dcgVTtd1rboN31NNP0anZBHTTeG5xvyVMF4P37QpUhncx0Ow9ZmtTmiKx12J
ZEhhN8RUnHEervUgehvKJuqVeysEfORHdVQktgN2rynl03OgfMaZa19q6bXr4xtASaMdXVi7CE7h
kpifrIw9tkETwXSyd5lxLppdIbvDT9OK0vKdmWM3pBh+Ej8BMoHWvAGaj2UU67QEMQ4lJkthHahB
/GzBUb1stB/OcRH+MWdvzRmDxJJmLQbYO3vWnE1rOM3VWezePDcB5Q7MkXMUaSw1HK1mvq6QONmH
iIxFnuvvj9SQmehl1qZuDanmOUos8ZgeZMpZ2iOWorVKv4oxomwPaPEhcn5skcZj8LlGxDZqU2YI
jFBg3pgCw/D8SCYb7XjeeZTwHyu7SIFP2+wnQuQTaIhF+l7fMo5PpxMQHRKnOZCpxIbTIpkRoDHS
jjB5DKcZmZ9lnsjh6XzZaigz062zvF9yjjVDw33m8IcXfKOAaHM7g1erur77InaUOHw3L1JjntzL
xQBLELsjO8qRi4/Tm+BQMbikisEpoAvzux+ToVYxynd/VKXr3gkwn+BKa09X93+l3MzJS8RQcAU+
AsPQa169AUlCwIHbshL3S4ZcDqANWD8yTRGsFj78uO9utNRnunEUToNP+nb4Ztm+ZAiIYGuU2tDx
FMPIvLpxrBZ2bKI859W02DMJXZ/VIjDL8MNEnZ4WvCHqhHkLHu27tf38luY06SjSQ8TmP8iBchtE
AyshJYq91UFmG/ST7HHChq0A9D2Bt95oTzbJr3vkPuxkkfGDbOwgAofkwiGhVbDAg+b1SRveFbSB
dtI4RCz0MPgVn7Hz0jfa11PKss+E/rPJMdISol/b+qwwwEm+HwEKSgG7WQmh+J2iD5b6SWnTD8xC
e7iN8uhhZpgU2C7yUmtKBIX7ilJ4YSe551Q0DH4083nxz1NKPPEJvFsZUwnZ4W/JF3teOolpk+1i
XNOSZ3QUVXobUfuR1d+YPp7cqqobRVY6bNLsHaWeSmx8/ToIVeS7/CFZRTZoQ2Q92MkmGwI7D0rD
U+5do+rYBiDTi9scU9OvkNVkFDlaeCBS2BVchc0iIRqxkdPvASnFwff2HJ5OTq580jabBg0HlvRj
gNHlaHeLoECAUcqBhDAQ+f3ZoOs4VDT+3q6qvDFOwr1GVTe5UzxedBA4RhuBlylCc2hG7hTtMj+z
et3OQ6Ng3FKX7XI0v0ZZlSu2G2ZLq2byWJBLzkxvBgdIQLnYx60Ssy/VBT6rRq+IpWI5pB+UfWww
uV59S4df8aXTdmNec+IENJ/ef5xEaZ/iO4KkDC4DkuslLsTnJ061a+ijiDHSZBdYzCmk8XMwT5yB
glcq5/tdoXy2TE88ttcwR2w7r29yUWWARXFBDqHDozm+HRDwxQMI2Jfd1V/xH+zD9ylqPUG5N1/X
e1WOeJ7pndpR+Y5xmUd3KBWQ3lVrzgd6TRjLo/nA2Nij48m1pTelvgY7+Ns+K8LdgkfpE51Es2Po
6QvE1OhlSfFZwN5/RMd3NUYnkRLHWf2X2BYJ4MC//BDtLIzI/DB9dB09chzYn0q2zobyLef0h57x
//A9uqAZ4iqCILYvAoRsAZZ/xCY0+y5xpmE7CoGw6HmF5XEgWxOzKQt3RL07LMsjUMHG2rrRFOO4
ZGjY4DCi+lSQ6VNqQIk3Xwm6PPqKVx2U2ZZ6t4gHRFO5C7++idf1SZqq5aSINVv4hZMhX+SyVEPD
Gi8rz0Ay2Yve1eXZMzXhKeiB9EXqRQJETTe+bI6GgbGcB3bshD9A5mI/YY0itR1s8loQJw4USfvI
56lEFlK/DK94g8KPo5xDPBiGqYjxRIg37dNAurC0bk7Zuy6cjb1U80d+CtNUescY3qu0dUSOhpvF
JWn3o6jxVXuzymahcnoCWdf5bgcOGVs/LoWvtZvfiRJudBEU1meU6Dx9Y+zgUod1t8juRIh53mjM
jfgaaudsgdcY5jAv5sd6sWT0jPsgvI3p4nQ9UjE4y+snIFo0MtuM+iR3Kur8/8pUQ6MTEFtz6Cy2
IrgXrLV1p6WRP0Q2LiBhcy/qoGPsFHR+32MIwll6bosucW4AaRg7OmcZQU2i3EoY53liCZn7ADzS
TkGCCav+Fdr+AOnKLsIefaWqJLhrzpv4tXgEkGYC0kUYF9BslewqFxK2HyYTZoRkEcDzmKShVTJv
/BeEYgLUcUcYiF35BJ4kslDlyoD4m3NdBj5WjRTE2LR7q6/qPyWldAMzI0qEShlfkDTlxDA17cah
nyZZhEVRU+8nJSNMYVI9+yo/zK3HJiu42osQa+KE/aydJ769z3S4lADXm4jbEAUBVmVS8kJBOfL4
VG3DMP1y9L1hDbz5sHeb3l2m2uvLbIVqmj7rLV23zk3KCgSivxo9BZa5yMGtObHlsp8vFQeBJHpP
mQTbr3aODrneA3Ee/9QDyw22ee/N8t9q7gKZMvQkL5S8iX+K1PuRJ5Yex7HApOvHY0f7pgICi/mW
hrOX+wx8Ta2DpcusE192f5Jz9G4P14Ix7fwZ4Z7v55f54zr26Fq4Hx3bbkzbecR3rpMX7VDsjDda
fEeROMDAf6Pwbx3PLlwZFBsfBi7UhNZtLsyaHAerwSuwjnRjgEgjAYD8mBv2o2NHLE0G23XU8Eu7
V2/y+e8Gzt6Qh5Dimisna6aYBnQDu89qFi6nBnv0DGxZ/amaW2g1DDA7b6c6DgPl2wbIZwZ6A1gZ
RM6D+gxpbunQZ5mJ+lw8BPo/p7LFbm71id1adoCTps2wUyxpS0mnuEfXAMmw8s8g/YTJQ4z7YNdb
MAEVI5XNYLk7CTK6xItCffyYwt/JR+v2zkkxUS3SVF2x5WE/3uNuEQZo86DcflFaI2GpjOom7n50
SU2TE66mUqzEOs2Uxe46WPHHPTORW/tRAU76MChPKzJbtC3ipj+kO+yJRwTXfzX1j1J/6CqtDEh1
oYmxZhwB8NLBweKiTNVVXicQhrdR4a9PJJiNJ/VbdbuUwHoqaGe1o5h1oSCHfdcSrAb5Z3M7nMxI
URC9gzxVYCGK1JvSMH/tk1tZ1CzTlM591+9AGQ38F0gVNwl8s9N0meMBUo1zKt11Fzf1ssqwdOd/
SRobqjufdp9sX0Cnm1dvh09nmMTudNdrA5kkGFR+jbIw/gVymfWElmqhjqfWIuO3VHJL0tyxl2Xl
JBDeQXGhj/UC7TgfLnoDjDCSltlrVmK/UXmBmSMXSEpd5FplF3BTMpSRK9/ibzFJ93IVW+IPLO8o
Z8EGgk+7NxHp8MINbLaSUTC8kJBdtSF4iMOcCtbthgEAQBMdvI+GwkXPMD7+LPyrY4JAeN9mkDGa
OfDxBQikFlwqKHKKfFJHJj/xXctLvOfH1F62f9BMAk/tp+ISE5F5Z3y9b6u54Xyi/zSLMpQ7vyNA
fY69+Mmde0VksjhFJaaVo4kNVao5nN8bOkmVfTdvRnGWtAOPMvin2e4daEMpg2I6ctOBZMkDJPQm
B8+d+HjtQQ+R1Q6Zi90roeMj3UbWT/5smyNYdvRUK0/IGzm2EI4goGAdNk1Rv/7X8mhEXsBA+5wi
T2W22Ah4XReRWQkkcBUhhKgtW/m6A3RlX0QI5oaNbGoTj4Aa1uRoz2gOeR/YR7Jgndah0/teRG9i
Unc796xv9j1tc/RBARqUu4FrGFTgnnvqjnZaR+4tb8k3bIAJYTcF0m04gNEjDhcWyIT5e/WB4PpC
oV1dajnB9iEAWdTRBfgU2qDQmdInO8P8COdFN4uxkw+xFEUrXu/FqlQDaW34PbRZjAjFELWneFQ2
C434BFLqa9AgFZvucU9jvBMM01/QZfNPAO8aJ2nBG58V+SXGJLoQOCkn/xFV7tnz48yCG8vR5+xQ
1u4D+XwA4GBioLM5Z0Pg9frl+PDPbP/yyt2rEwWpE3DaKoPyTQsJRXEBONSLYw7eZQgeYZCkIxaP
leUqs8TcQeP3TsKvDRPgYp9D0hWdfcThws4mZHJz6H0QQxSU8SE9ApD4zllpH1gNRQQbQNwjtrxk
eMQbTGrAhG2WZqL7x3ABVv50byrFRDEHXcsxAHmUxzwq/E5R2e9UgqVvPMziYO0jGX4Urmlg9AZQ
vUlig2hviebfVJ6vqwvqVUcIYndZ+h8SF8HvymiODUoRTnlWJojHMZ2/SuPAeO+CSBj/xwRH4NbD
t6F2ArAAGchJ3XmCyDzrX7PHqjnvZ5tfMi+0D+154k64OTLh9/f1ZMaESoXgZbhnt75fMAsdZ10l
3PXsc9L4n1d2JdpVq0xnkOds+3O+wv6d76HUvMtapLtsSTuF3t9spPEUWJHGj85nmjxRTGHb6/mP
oNX+i757rvX6oyf/9HiT3jb4/VMuYRhY5Q3gULrvFvNJSBK2mRRdlOdsfvXS9RwPOOfPhfHIhTcA
Zr6yH0vpyKgraTvNVR97LWroF/SEBkxPlUMo9pqeYoGCdKAcVJ6vZ82M5OC3yXTPirBigdCNzDKv
mZg86nwusI3oBJ0kB1xrh9d6a7/Dkt5w4D5a4jMv3DxD39QA87opHC79YGVUH+1Sd8Fkh30E1Z3/
1wya7g++GuOppQmR4PmaLbMy453bExzlM3ow7cRBrG9HfoHSRZaCTI+zw3sMOAPYksvmYjWBRDYO
8918t0HcrvrE9uUoPnyIshnTEc5w9uKllKzdUnsAGcHug9lKbrFk3aNDxrH9WYg4/dKM59MPUJq3
tQZ9nNYl+w/GfCsdbL46mbNMkDXuMywmXDyLj6HZOzKQrut6mgf6EnuEktM0+y9oAebq5pG8/vLD
7COxq5oOhsQUcwmshhoG2MsaEgH/Y3DNnpyrrGEYqxlSId8C8BI8TtjShbhEmr/CWa2uS9f75cMK
4vYueAwSfaSdCVE+87ZsDRUvfSeVUPtWzFe6xK02hh2DibB6my8OGjhGmK9vvpd2knTg32JT/Vp1
f/3XjfPkrXTInrj7zzO3ceAnFTF56MI2/GIL7xXW1Jcf1eHEHC3KEko/72L++HclQgahunQQzJKj
mC4lNnhaCRIvjTibFxzPPYL2RInLl3fLuokQYNxj4HQn6Whep1ywFUw8kWDbwOK7Z1yoTFmWmJfD
5jN2DrGR4N91fwPmVTH5SymmYqGMU1vbpbHUG4iK3V1Z6QmPXG8CJ3n48AnklfexC1vkrBWYjvBY
HveF62S/NOpqPFbgR4aegF11cXVhqSWr2GwSEL1Nrr6WhZ0oPkzipMd11/eJjB6/O/hEl9U5/A1s
oRi5R3/77VOysdk7TGnw2IRVFI98NfOyKQukETVbx/DohQLS+B6L0RNIXj4Qu6psBjU3DOmStAGY
9arS+J4mXPgnxZ9eQmP336oK3nejEKaWCJtXX1QsTmQKSiFISQz17T7T3ueVCGQlxEWt1bPCcbQU
U+mS4vHyXIV929pTEV9+cLW2jrqs/o4vhbhp9g0Pqc7lUGTmtGFrHQZT0KX+BR/O4AKBl/YGoclO
O9KOuoV+1P1P36xOWcgtvz38N0jfwrdlZ04N/IglkX5FCUb2lbz1sXqxLdTVNgZr+Zizl3od85wU
qABw0TDLDTmCGj9R3oThr307sIhYmakW8AipqPNZEi4FetaKMgdXuCUraCdKIf8FmqCfbNNwuEIV
+/0rBj1c0E2EJ3BdOxm6l3ai7uedCoXi/tfwpankKf2F22Rnn62meoWTlp9R3IgIHUsf0QEpk1fK
Uq5/OGASV0G5UuwZjVtljoVlhWO0KsLnemrXWyll0rtq/6R/DzrM5PVr4aQRmxGKVEDFUGzO4Wu1
dp5qsV5Yrd7HMFECZ4JYsXbRkDBO/s3ApQmwN0DiHKLXBVtbhp2aGbxjNTrr2MyBrkTky95BmfPB
eaRwobSiiynJPd7Js/J8ADmihgW/0TV6V20UIQICWQTNzhSGkryTCQGhiFOryV5DmJMVZn969Fjq
18Z5baj81+VCU0d5RBRluvT7uo/FNvgsXzVsBJFvm8EwkTo1jWme9ANCdtzCLFGWFQDNPKf2GAXH
AgqRXDOCAn16qLvPAvzNFXKTCw/OLeFN6RP7d6rUm1QuhGAcTaArrcLzZdIaVUTMGt1aDWIp2p7Q
XAcQoyQRCPtaedHX4hxecXwYcsgpB/P0sBpOtUechduhA3d178Z7FqVO9q4Myes3aXVyjjmw6k81
+QDOq/E+3Hw7hFt8OIxP/0U1ygQZM68pGRP29vLwEp9Q4f1ZrMEwyOgfNtqDk9/lgCiKgx2hOK9z
qQXwopzQok65L+rBCZMmo4F06mVlObCrN0ywlyRjn/YzRpNnkIVk3k4rxRP3JdYLEnrXT+5Yd9ww
QFx2RAtEbmMPUzi7NpchTTkoDFjsftDWnD2EaoaYk7YvMH7SdT2JAydkberzwI8TahMh0Zb9pL47
3rTnI4Uffo2ruDdLWXRKvfoe5aeNNCULRhBKIDyxlVgekg9NKWE/G7zRPKodQXcybDlFPJ/AA0xz
cyGp0rTEsQJLawYn8+kOQJp2ovGA5RmHf5GMU9J8EZ01CBx/xRQyo197splbsULA9Ddzh3g+4bZL
XDZY2obaq6r6Eqxhq2VVdmNp8u0rBqBduLgceqZPPW4G9gthgknq1tcqwiGLB9CYEPF3F2HYBlNr
tJUS7Wxaww+8OCwrCvNq0V15GcKHP41bR6/rMwg4Kl39p7OfFBsXI3e2dpqTrD/I4w09/a5k/DXp
Ih7hZNhODUVAyb78Hv5Ip8o43A7s/XKsD5dv8La1Lx7TdCBpFu436WuJBmWIMpMEISrmtzb+/Ugo
cwnEJORBxP5bhRsVzZbfo2HSmBbaFM4McFkCRvW/o2fuNy3a73BEZcKz5rSJU1FfDCMdxEAAaqQO
JyTUb/hdWQBnPDDUc4CDswex6lcv0YhAex24q2fhYu82q+spG5oYx/rqufOKP/Sc0q5l6WemnkYF
c7A9WmliE6FTPMkTGZyk8e36GzAR9j9vXmrSggWuwurjkC67HMY0/FtObHnu2SzanOhhSCLWNYjd
JgCro0g3S5FLSZN0UqiIyF2vJlzapSjEAlJ7oh3xc5CjSWBdE2IZCYGhtT8ajBOdMyK3tgtGeiGL
ZV7JD+Cbg9yC66Wc+Fjsvz/oA9VwjRP9csn2RyhYm4bCFlYZqUM0zqzloZSjy59lmsD9ctpyoEt0
OSD/D7c9eE0WnEF7XETXHAPxIxvfC76hi8usDMGbzDDkw4t4S6vW57qj3LLs3+RZ1pOj4Y1opprq
NeHOORMBSjOOPXgvVY15V1ffbdKBqmtCN1mY50O0iii8ey0yNfyi4YRmOKQWJVhkl5dmWkb/2c4W
NYjkdRQfDoDoPxE5sKBrZaNx9grfGO9ODLJzHAtH2Q7H2iWm5Zl29AXDzjBuKhRHku8TqqVunO/x
WZeXiGoAH/6vX548Uo5exjpVWRIq9FOMmIuanr5OwkloPNRSupRSm3QmxA0VR8dgwdv3uUtK94sQ
Od4mlDRzAVSiDcby4Fklyf89Pn38lvAOrWLruR+7zstrwESYtWV6gLrUoIs7MBOxloDwkCtXIdZu
6uYHVMo6nXgkXbbLfE6jBKvC2qnr/XOP+pazaHX52YhiVmIniMvp18/juy2wIifUXSO8Gmt/+uo2
fY3P2fUIsgooBFa4x7KAQmz4os6if/R9ajim9DEznX7j5VrNt56qImlm/856GAMoHKG7aTlem3y1
/XWdcyJKhK7j6o7ctanKCdgBiI7r+3Gb3+bQjsd9tZPjv4P7WkIflpa1swGCjnLmMMR9I6ZXZRaE
POdgPGxv7Hfw+WJmibf9sDNsKhcrstg72+lt7BxFangMCLOzC1YE2UpZ7oi6mxan9u4o3R91rB4d
1QGbr6hQDs8nT7X9fXW9uIgOZNmOjhjXxbZPq1+vK4QW4HHLDZt7MIT+UwBgWpaeWBwptZaFmMZr
MNQ4JYX4EWSiKSbdm7IqJZ+tdY1Er3vwzC1gk0JGN7L13FaQ8MQctLurHUkPed7g/v/gRsznH5mv
0MsJ3g4s0IOW8XgN5c0bIFkXlYHhT1OCZvIdXS7+tVU1o1yISweePHDSTLJbpDPkr2BuPatZ3EHm
EJ7F5ve6gqg/6WrpnPJs+pJiA1b2n8WzpXtAN8xcz4Iu7IFzhYc7VubwgJ3Wc3SjPw0OiPuva/9N
2TcK3zzZyquP0zSk8x5lFGVJJKZC/J0fUL6no/3Xkz+PvGXjnRyuO7EVitQjtdGRNF/yPBniEePo
FybUYtB998gXfyY4pnbY650QVFCUYegFxO+17kpvozv1p3eFu28JsbFlJj3Em/+hMyzQJX6vIxKO
jfulyaNSgvX0F34w50NUvrXG4lO6QOMFoKnkfLnp8QP4uEV6ZaWTfg5oqHnUdZ3opky8IXi+37O2
lB19PvEj7Ax6n7iMKEEtFw4dIip0kyyVsxNSTXhGIyiZaaX8rvUY5U9hpLwGtj6T+1rRpYmmBcHw
EfWVdqsJ9RaD3vVrVTqJu7Wf/uiQsnyVJAjj3hspLwHe+rrWjKbB1NZYbc06n9srhi1GtiKcmlLD
/kmYNyqKIcsgBOt8FeJTmX2/HY3QTJGZiDQ8Oa5c6XVGEzqwSRlzog5WVpFsrLVYoJQxkuG9RHIX
7AT0K3js0dGMT8P5/VTRDzsAKyBRjdscwM60cV0JUg+sU7nceo1IuwQYGioHbgCiCclfaQ6kTKjF
XINqXKdJA2dprDFyYRBzZNGriQ8+OGwzh+bmBxtDibGkJL4TKKYKcgjCQGzfyZfFfUB8Xxi0W99J
Lyn7EKyr0Dpfxig5zHAPspNHe+pQaRV4CBJZJZggkAsoovVgwC3+eX1FQBE182Zn6G+W+cXRmYnK
OwKBbmY2AXTKZM+FW68QccSzn15NZKU/+hxDIJo9Q426Q9irHIXexda0BdIb/jhDpRBC06I5NkO8
vPLyxeWnvyqcRlSy8lpBBW+5XeIo6vJb8VdtpZE3zdv5heLP8rtmu7Yd9bIFH5CvWPAhfobTJX43
oJSQI8NS0ZymVeOrR8GZgb2oW0o2BjVwRgS1KAAj7rsRul2MeqRuAJvUsvs2JAnfDiEvJUGhI+1S
FMmMCNUoLJCWNDEpjMgT2xiowTLOprCNYr7fyJtFAA8mjNcS5KBSA1Ip6K1aG0/YNP2VBQJKgrIA
Zlzt4YRWLG5diq439k+a3e0UgSJ/bQhwv1HawR3INlUNm+ynfKQ9dBRubwh1/Uduc9RS3IWNqVeb
Sho060ANY66uflQD8JRiXLZe/87BtbkYwROcTb+E6aWy3KSv9aPb8J0xlE+n/hqkarE0VkC/LCQV
353QEnvBinZoQ2OPxs6WHbcQcbDCUtIZW0rLh2TqS07qZb+l9dem1OP1BqLenf9n86I0+B0C3FFT
GqWZv9FEFAoj4Vrp0pyOqaFEY3M3SCCcyw8+OkEdfr3DWspEsbbjV+Oi0p6JVJSa7i5BYVIWkF1A
QGLJ87D86hfnSAJY9yZFP754xLPYc+HNF1SfLZv7RQwh5AoojisBpWAUXdRaPyEso6dN0VY77H3/
gkAku/eXQ1ePn+tB2+gPPJru7WfXisXH5EDFFdzVrntOz55A1gHtYgwZoZXwBs3k8HtA1vILIRVP
Lg0wYhusETVgk5cN7idggHdSjHTd8OEoDCgROpoxgWVTuG0F6FPAq9lJv3LevO4+Wyqc565g/Dyk
gtIQ5VulL2uscMMpWqwSeWicQrjxijmogsXCSAgcEn5AzP2eeGL2lEk5TLOYegqsGzMSqVeCVUFi
PswENaGzuHalGuVX+jXjqDppboZIACsuswEXmWWDgDDpGzzdyrCR6oQkH5tbHklAmUKSgawzoj0J
+gUqaKVMga1zYJ8kkw4RDJIRAq6ZWrNPTOPyllAwsVyAcZyc9xP47KcfGnthYNVTPPEHWhJfXGkK
8HIs2a6pSWklAbgywwr5Y9X6YjNXIfyPyA37hPofE3lyXJB9c/+N8ZXbYeTk80R/kNhkY7XAThxc
xstj0J/NGnQ/AqLk/ofhoGKN7yPZ2NRt8V05bJzUa1jYtTTnG5VwCqPx7MW25Ehu8l7szmvm9qzm
FH4RA16yKJdYbv63WFxRxOI488S6SwOdWe4exW/9DwqhWG1UxaueMo1UjhxJWOMmDZvIIzMVWs2b
OwWhkEOIV02lUVKJqhFfWUuzUCkyY2eU1fEEWh8h8rDiO3TZFgMmW5EFhBzUVBLgFGVZxa8vrqNe
Eu3RWvph6F2ECSEPeFfGsWetD5iyqelPHMSrCW6wciY5ylpK1xoNx45OdTVquo4V3q5J27AgwRcA
+LwXlxf7sM/ZSrbeXVqIwJvEaQsdBopSeivdSdecBnhP8h6rYtD1Fg3UCf0fJez/yMjng2ZpjpF2
j2URHY5Ll4VLO34DDOMxs09MtoJq6/+ANz23irwdkk9gnd07gp4v+wSvO7gn6zTOYpVdI1yWvVF9
DlxP8dUeWKLHOYhDZbrg96t67ZLW46PeZ/fDo3u27aYM09/5me2qAE4P6bfNYEbFu34zUVrYLSJh
dHdo5qQ+c1YRsLRzkLreBdiuEliPIh/9nPdr8meH56oWznBrxmaiPvv9fWpI7Ha5PRBDyuLXMIbt
w35WijBKagqhYt7kzoXQUsyTqe3N44RMLnqLc1jcrR5c0ulfAY6h04EL3MHZalHx2N10mj+lxVNS
pGP8Ds1bdv5izEbOEkvBOPYRCrn4ybj1jHrNUlZVC+h3LSnm1lsZtkT6NxieMcRg4sDnA4aEO2ln
yTHHn6tW8hBy9mcDcFptXxZIBeMspjjCqf4l/+sWSfQ5atPoraHThDODiXp88t7jFm1jg1XHiHTY
uOLNEJsfqgaVaQD6fcw4QJA2TAVlT/H/4w7pZvzSksciGpwNWUCuAOpxUVAWMW4+vFq15+Mltls9
eAsxkl/UgQZiIldh3VixT3TLrX8iLrWTJ6eUywncmVYbkOihHecf72uZUxcuUxsPE2umjfPQfH8p
FlN5gueF1q5d353lKObd6MzUYCiAJGFN5PYwF8xgbGKf1JETcQRN/NoYLw5f3rzUJYocaKu+MjPk
meZ2Zw91mDAku6V+bwqMe9OTkoLWvR6nSqutVPzKwhoYg+2OdL/5fXyaoGWQjFDIaDM1zpFEcQpi
+BpZmncNcKhsAd8lRf4zEP99UMUkPCYekqBpnRNKSyxV0Y+G6tiBJuK+onK5bD/0ENGQFjVkBYvT
PP5DwrnkkFvNUdHjB5pH8rnrghLHD9FtdOdLU6prsUNt90cu1ymMV2QnzOTPgcPdpacMs4AYn0aT
TANylfDnCixqoDxdOqCpc3vlwre/1Ud91Mip9KUWjzuRa8KkdpkB3wAdkSAx0FloEWIR6oWxHAkO
fNxrU8hyso0MNd6Q2JkQyg9oPRIhhLL0z60e47As4O2EwzkOai7KuGOq0kdXlvqsVPXnkpXwje/0
gN0R+95JHCnRLy0W8IH+TI4YNhSk9lxslAkUaK609zc/BwgGKYtprln+UfbxpAkzmzOongCIBMvk
IRH/soYa1L7WxTFoPhLG2JcuZBJ1XZ0JAbUXMyaYZhLWWpjIREV29/peIG9G2Jq0fY4hjPZdelEs
+NMEETkVf2yitBaKVvEL6wf80XSjUOXeLaQv7kQFRlPr17EzLR2l4gkTvgVWqgclvmFteK2/kgTJ
tan5+/TIv601sw6yKrN17BvzloGodaw02wGjWPb7t4/D5nwdtyY9M0davYLclLOEqMLFMlCMG6Rb
mSZ5qdLqN2904ehWB+Cpi/+J3THlngeh6IglZUV7ckZvRCpNcu0H6P1AaY2zdACwGt1w+3sItqNT
F1tu6gh4rnw4g2YkmkIz/SUVbTj/b6FnkR8vaxIOG9bgNYdw/wbiOzsPl52Vb45igXjJsvVIDncl
mTOoGeT6Cok8MIk5utzXjVd/f1lbSL1PK8eSa6qYyfeVkeh0/A29Z/677gVrCfQyiz/E+RPB5Qbn
HNS4Rp4DPPm/+8RDtQsi8oxgrsQ3Lnih+gbignsC/i/BwDFVxEflT366cM+JUm/8GeV3wnM1xkzb
L199wy6XWR8P/r6QdiSXhNQx9DaZG6lxJZ0w6zVHh3SHKe2vdPmmvVwbFiI/YfmmLq7HJOs8cj81
OVPpe4eRqo2TTva3k+D307CxGI2ErAiRAgNKbYdbucM48D2YidXo2qh+2AD8SYKHCWztc2vnC6y/
VA8Ww8r6F3/TAm6ik+N6XtXVSSwzT9AsSopVG4vJXxjqS8FWGjAzsE8roS9TiHHJmY1Iv/mrn9tZ
u9gIiHcQnhFXad6+jRS6Gd77HyWkEi5u0pFJlzXANLYA0ldyY5JFsvGqeErUzizo+mxJ36A7wviy
l+KVnfoEnZlz/9ci+/+0fncnbCnEJaLYrHNqQwK1t10GllCnhMBttdav0AbCzp/e6QkFr6o85XqJ
YW0oaze+DkXurndVdHj/U51Jlyu20Hk0tH/Qltrlh/Jpi8ZPtH1GH6qb50CN8n5LV/eaHvFclu0m
oLqGCQ5tJCcnGyCZMYojbPRJXlUQXac9ZopqwJQ3UNXzYEGrYyx9ggIFr2bs/eXrMNk/RfQ8iXPT
1IHr0GRw+UHr15VugW+TS4wRFejH3fwLAdB0McsPnAVj6h2+z5Se8g/UgXf7MnIkxz15Jlnn2nQM
3heMb46Kn5f9+Do5P8vevzcKGilkyYANbjW8CIxEoH79/JshdTi1fGmQubcLBxkOYvAAzzk7gBxW
JpIbaDS2Jz6aZlk6AVHcd2sYphvPEitMKj8VS16uhoz/ndYyx5noJWIhvg9y+NFExPy62Z+sY+sQ
b1JA2GYh+2+UV3VX+87HA50I3uhoeMHDkLZAE7v0wMIIh6JpnIhJQKbMzU4MT/JTV6jTx6kT8foi
eZw5E+hKO68Q/8EwCt9GvKA9nEJT3COpM27HVcHk2tiIXeWVgCl8s1zC3oDuUM2t6ZS7+173nSXm
BhxbagAhX/muAEzwpKnfV9UDmy4MDhVruVHOOlOImHffYnlZ5jOpwNMsNiLnJX1+Dch8u9KAAU0y
dejpVuS5QJwNQhh1SyGNFNLNPa2Q37YC2MH4dpAqOlDksSghyRjgsiswmzm8QAlt/n7+CdjM8Ds1
4TXjfI0YPWQ1Yhk1oRZ+CYHw99ttZmIyBjaLJEaBEcs7zLRQYdKYd7MweORZiazL5EcJzgtR/Jkn
OVADo0heCTsBtGikPmu+R76aOq7dIpZ3BHW/RTla9BfN9q8XvlGTS4EPJv4nR34WkEX+N19jOOtV
TOs/2hyz5dAWcjEelNeK3NnLd7cvPGr/RYqw2nTCmPs6Zsgivy+Jo7CXSkPRrP0181Nu/61nkXZi
+JRjIMW9ogBYaEgKHN9Gk9TuB40IZiEd+lFqytDhPSUDStVX8IuKTzLab7Aky14IEXOJYkJo0lSX
HL6u8xZyh6CE/JPikdvXlQZu6IJLSqI9dT4Xh73d+JebLGeJrjIhiXvwd3lEym4njqIkCul6d6li
k948vCTI1l5PHGWPboiK5nTwUm1Q9ideEoUvi8w8QxeyH9NeuWa3vZksiiNuRwQ63nU2T8b8bpqR
km6WZrUwZQMB5jb7GQER6FZBpnPuj419K5HpdpT6YoIdcvsm+PlUmQ9pOzD6aqiTzQEbifFsBo0y
uMhnrTkK612fcIlgMrB6oiMGZdWnpxp77Ii939N4ODAjDvzjW7rU/4kHUCVH3HMUMD/LxgmKiva3
WqzNrlLzi+I3BgfoSvEPm27EAsrXGYaj0s8Jf+S5woyoAZdKOr5H2lprV87hm7/Cy/03QlvvFuqw
SZxgVF3NpPKb9zVGwk0V54Y8bbjyGhS0/ZckQCFhbTGwFqkparcdPPxDYJmqgxRroLo76DvB16GS
9HR73451ZGkt3Wry7vlvPpGk+N4WiGmxrv4ScipY3a8fs1AliowI9sfT4/Uq1PskTodzQk8eo+Rm
gUGSGLNoLzc9A8j5BE8vLokvBmvU2wWxB9IM8zbfOwEPialg2ZAGz8M+FoW1W7fZRa39PdF2GvCh
eC8GEWkcW/B/CXWzj9prJuxDZyHpG9uZxZFsXcHwMznrcDd87niKnf9E9Oei5J63Anj7zkAWyxGs
13oMbgoqAUypZ0tTOcgbEWYio/CwJ2yhnYzr0WZR1mZPuJbwSQMN+1/BAZ2LXMXKEW+vLFMhWdw4
lZ1FKun6Ld3vxuOmSOCJPuKAJK455gI5ZI4iHOe7NQV3g6g6d1quqYvIFYp0H3G+L7Ak/5dYTFi1
Hr7OYnNC5y/PZiG3/vgBziAcVvh5ctDa/kFwZ+vL4QIeq0RABxppu4VpJ62tzdJxsbMh28Q5viqE
E+5073K0Oa1diDDW1cTDjs7fDkA9av2dg2At8djcFZSB+MR0WLTo8uErjvASiGcnlypWBNeQoobr
WaorrmXdEyl3vMFBd85dVldbtxbY5LsmH5ZHfhPremAzyZX+Rbo+v+aj4iD/ld3UYZRRfDbSwIkd
ILUN5o1szYa+YKX+U1QWwMC4LJvE3Q3gH7bmmJLCHJ/TwmShLwqczkvL2BDhHQUer05C/4R1CstY
gGqajI6FOLrkWnjDpAq2mTnm7cbv1Sn8Tbvf5v1+KSblDniUpxzysT9hfwFlhDxc8sALzuueVHTP
bqATcTihZ3xHl6QEOHgv5m9ov6YMLQFflxfGMPfHmqCgs/N9kczL+oX0Fq2mcwMLKLkSONYikRBj
pUJC6cCNOawhXBhZH0FdlG+YYFP76IDVA+tXrABSseLZrQNrMFjtp72/kYpMevEMmPz1ep9cG41a
7W9PYID48aoyBqykM6HcoZMmBPPemnLJWuoEfHruQQ7SWQpI7o4wMEbcM0sSEp5Pu7muy3LI1Xz/
+8Xp3Poh8LpvBS92LHJg8AT1bYkPCLG/KDSevkZ+WD/KO0/iTlSkPK7VVyY5GRDeyCwLXSjkel/A
2si0D1/KF/SGE4RwKMnXyOBdtfsKpblbOOyvBGNc2aHm1iwY/cns1fRlLvYugy23TgjUvCMA5GDH
YF0dV6KkZtY1fA/PxjkKbgpLluQ6EuslBb5GxyK3Fze0qStkQr0m1SqmPgXhfhwN9MPg8gTcSAO3
3wQfKq5qJDDHrvDBWoMjkGAIlG4NOetuTBWjNxj/nF36W+/72jAFfXBj+M06/rbbs1pV6/Xcpafd
uT5FOiQosngwujzKObClILE1C2kMuKKYFIBC73BH0twyBDu03u8kYRs9MQD+hCbFsAMStHyQFunT
caEUHtRim+5baLZIaU+iPBpBmsXXF2KSi6+eWdUNT9zTN0fr5Qk8tPo636kj/mlsUS6ibP55rq01
xho05Kq3YGvWm2Qjroo0WA4gA8+w2evxEU67mQt9krnA6oZ4ywUxfaBE5xLUTofS72EXjdwqsXtk
2pia2zsBK2DcYcIdfrcCUnO6ED7QdPnJCzhgFxoP/oV5LWmTix6vc+N82OEMwIAiZCviWXvuO0SB
whIrg83d/EE+bzrbMgNuBOX7877rgpO7LG/Uv8SRXPj0GXwof2quCFIRtFAXlDolqGabh07HutL8
Wrk9CCpx06Ivcw3QmlJCUM/mDjwvQC77nup+3SmkRZLXoV6MP7FmO7uprI4C6iGF6lweisHli/US
swdo2nEnzC1ZC43EN+SosLoKj1gQZlm3F7e3uEo0CZqEc19aqGluFU/oInNVn6Szi8fzOA+9am4+
d7R6D5nZZ3NUCUgCSYAFjVtyTBs+8e4lchGplxBH7uyHTPJHmaBuRNy4lbn9WWhb/3o9pbPKkLge
At4mTNj7OZvGfLjNjBqwMq4DywpgRYrW7oXWsH31kcONDvsmVWFGbTNLhuEm07EetT1GUIxJLwIe
/Y/Bt/xco8BbHG7ui/THhIR30a7XthNqwhDkf61Pju9sZqg9eraaMqYxyp6kiIFpeTnKfYqOLM4e
eBB0tytQiZb2upv8Ha7DVjcS8XUkRUCyc/IZYa02c6udiUebXbcVA7MuTOkGqb6zEohMNpHjGRym
FVXCcsiRo74Vgzqy9CdZMMGcHq/UOwI9czfFU0xR42fKpLIQ8K6/SwjlPQTAkBdUopy6d6t/c4Xm
Ly5wiNOYhRgq2RP716BXzypRQfaKDYLe5FYI8LuRpuJHz6Kc2XRXLYPMzyLIeDpr7AoKOSTN4Fcd
KKKtVasGmOvL8S8oUr3lp2Eh43adnXTMw5RVF48Nk+WzRiBNxRuWecFEPmwJAyJ7o1PVju3nXD4j
o0lhXAqCdn3ePYikHrPf/jznJA4jsVlu28hv2sq/WhR2ITgljh849G2gfH8LhQtjqMV3B98N+Sbk
KvpS/tbQ5NYNhaLTTj15WtaEYRul1slRCYBF+Qe5SRQ47xed6j7PL33K/bnzqXaQYg2ksLpUZ6yB
ktLq+kh40ZDHhCpEFtC7zWWKr6TmWdRODx8TMSZxDiByoxDS3FtweTTBB++LYLIdopwJqfthF7wX
2Dpm6GhUC9Xg5qruvvFH/Y1JT02R0ADpNWmFUW1WHbHjONpnqDYtR4lhXtq35fEqqEBu9avAC18q
Fwxs+BiBHhZnoIupunWm9STCOmtvEuFIP5XPWbdwTh2vMBhdueVtOxC3eITAaTTbOIYO7b/TrAwo
7DvAPU6aWacnQB0Hpbz7BhsJW87deai6ApyDGSk3Q0PXKXRdaCl+cnRMVMcQ8wJT+0/+E687Igna
INtuUNlM8AM8YF6sM/ejJDDQjw9RO+ISyFEj+z3ilw7Q8sAeq1JKF20NqqJq/PSM7N3WTKgVVZ5h
wfvf5cJaf4DVnqqOIyot25Lm6yf0MfjMdvLuVbAqr9JfmXkkZaB4tFyaCQUq2Qq6YUMYmiRmwH3n
3fsdjWS+kkwHR9ZWcvptuefUN8iepaCHuB2hfAyNwYZlQ1BOtu7zXMcgXxD8DX2LEeTlMx98jpfc
HoxXaRHumIzHRf6fRoEYREWwJqW99VAE9Cy07E2Pb2A4UUCpWjinnZ+MhIvlEufL/WyvBBRUP/6j
YIdw/qLJ6X3OEoWBXSSWsdvnDA8erZ4uEy1Ma3yj40t16gjv15wDJSH+L73/SzQHEvU98evLJD0g
70VHkNuswvdDMAUnU9XH+zPqem8hZIpCYdhDuEq51kxk6NsupFWRM7mhLR03JNO8TC1C02dnikx5
igXoE7a9Pt6GvTXOKigD8VOsa19kdHhmMVSnq0zeu8H+8pKRRguc2tVocy60DJEWKey/DwyDSZ2g
PxNgJIAIcXs3RmwqjNWaHqKbkB384Y7eWEYO5jEH0CbpfGIS3P00Um7oG7xOr3V1WaoVRSIAgceC
h7POTkY+IlKVzLhx4j6RAfTdnHuHr8dwyJvEQaFpBfDpttKodTcB2KJUAWToZ/IYY3d5serHK7Kr
zVocgcv4fBL1TLDlnEu0FQyktVGqId9WYi6aOm6tVd3qo7Yap/+k/FidNL52xC3NBafw78QDHHwK
/VsyyeTjwAVXJZ8sN9BtQdnB8y7NzkmhPksQTeeH1cIkDTmpfjJ5vN23zLUGr9eqjmNWL7qXTsVx
byXCrAiSlqyD7Q2vYAtnt8wTmYpzCfON3CK5XeIM0i955PahYmhvbqmRZeiznunQyNdMANlDhKb8
OtxRoESdD1MRysUjJPrEjCK/Yexmon0LMPh2hVjwg65Ug8u3PjzoHlQaNpatnpcvXKe+7IFG+XaM
GamUwq1G5i12vsZKKl1N8KNAIwb4tKewyr1e4F/3B5VwIWS9V6O+F4JyYy0OFPjzCfLEt+lINX0F
K6dy5jCo+l+rGrZCUr/YspVPA69CVt+AJ5SGWL29yAIIJ8J6TbN4XqcDLLfcxagt6g3IwxSSGuwf
bXf42knTF6CbCk3H/r5YMl71T0p0D5BThuaoR5eizZwz6UNqu+j/p3HojPJZJI3pJBg07uKbB1rj
wYRwXF6UjRBKMFdEZ/f8KilqKG/VWfz/AD8aLwt8MOL3vYNj3mWs9DiVmrcRgC/6kcS69Nt4rQz6
o7JN/SH/yGYTrXDaILwIfjmPlLgdp4FkItBnNWBo54kxA3vw9UnVD41uQaBqSaL2jzTrAykDaSKS
nn6xriwSMLO4Qtje9qnkGdjiias+AfUEXBjlkNUdFrsolu/MNS4Zs7uUeur4U+x89gf9Xb/SCExN
v0pZ7BXQ9+tepJ1F/8gXqItZChkEuO7Hmn9B2CJVzYyU6qrLNYN4f0rOxl37eCkyqskLBqj0ChAT
1rNy7PS5OVTM0N7NV2FYsiAb2/FyrtR5Yp/7dSdPVxQBmFQmUUxh6J2Vw9KYGI2xSU9yQbvLINRJ
vrPVlzYywBDrZxGCcJaOZprL1tQ+C78xN350t4fnzVmgMxOCP4RVGiPPSo6g4VbE2GAOtoOqAZmW
XlPUGiZBRZH/0C7Mi7bgTnwIW+dJXB9pMsL63GlCF9+NcCxMRW0GqxwrjQ3/S5ojQXCaIqzXARE3
TXOm3TBojcQ2M32cOE6gDAVAsPWBcGuf8GlbsH6PLfNseeQ24VqfV7hIqkzOraUBpeb0UPayuS7c
ZZEWeA9Xv9rxmMGMmdrxoo+XGcXW85+gzEHFKGYQ+bsNr2K9WkCU+bbx01MaHKC1f7NdirHJTwIr
LD6UyJPfpCcs3H1GheumknxujxMgB/n5FOunuZykaQqpKds6N5lcEHVuANW9SWfgFk8LJ5hhl734
FbkehwYNVqPSjy4zx0Qcgz/5kgEM2CzhbP8PcV8HGibdZ7EWtet7nIjaEqkXBsSNeN7bPrNE0p1v
0CmDP1HCwLfSbhNBATdx1kKxkKfFbkIbuL74VwWuzX/2nRgNA2gnlJlpHx+KRD6ALv0QtdG1mBOM
rATja9CPWmPv1ABWD6OeK+qtkBLmgyu0w4MOn6LveIoOGWWZ2zj0toFpall1WYxshRK/rFN4FooA
NP9XLDLQzLqBMDpQgQliy9TyH/H71dX88q5jKm0sBTHi7paPEqcaet/Ufl6Fq3C8EwioWOKC5GLK
u4iVlWC8Evexr/aubgUHCH8Eh2UzCSJvwFuuiOYpyK0NF70I8OL0/Q4yMxZghhbnkD+9jcuh6Fj5
LM4jddWzSOv5Rat/Kai8pUqy0nDDfzJWiC7vavEWNj4wsyEmAwKepJd1KBxnHGG8j2X45E/vHgJP
mrcjCJpY7RNvEyBa28g1GQLotEnGRxwU4O98Xvzc65Z1Z77RvUoRqsyUctvJqEEjccoNAs4u0rDs
V1x1FXT7dVM1M47m8a6M8O/FGt0dMLlq3Yx3hUAcJp+KzZXrygnT63Aq+ImvWca6Y3Cq1VbkOycR
RAVoIVjLqqKu6ql6VTdVsPFscg8hFUWqOtz4H0bxkCwK47Z6SjGouQaJ4rK0cZyv0piJPs/ybjya
SQSkH3/KirAUwgXbKmsl7FVX41ronNLkxzEyfWK6SGGLX1xlHiP39S6zJR52LqZodDrnMijL1lZp
vXte+kTzAclAwjGlL2tXvZys2BUAVBYXq1iQpY+teQe9+JuposFUr/rSFJ/U6ZvBcvJ2Mg1ZzAIj
HXgmGUPeKHqkodXJJDavgVBpXvNxf4J2uXCHL3nXnEn9PDJMfWWcQDUJD0nz92C4STklrqSTFVjB
vllVVfd73zNPjddWU6lxkubKjOfeQW6z3K3lBrPsgWyjF4aYLZBqwLaFHCntl0DdunuYm/NgBp3L
FO8h6bcktwE0tAxRfPpwrlubyUgwxPeJAqxAcsPBiOizvPgwLddhtGQspGxdtQgLJ8EyYm2ODH2t
n3L4RqfSMbY+/9zYjxNYv3HzmucRGawnJVHpTFm4ADKHRXTK0UjIuSFbw45tShu0i1Zc4OfnOz11
VkZLy5o29n5KjSKfxVWDNVK9DlXwUqRSsmBww/kDGkgCeOrm2nErWs8KwJxgVw6eciDtO65R1APG
z1YgAGXDb+oNiv/039b/J06NQd3G6gePJpRcDIwqDn+4YiJL1kThavSBZhiuHuijG1s4uWkbwuLw
mYSkOtZhfy9oNh3GNKrj27MQz7ctmcvQ5ibdLUg28K+mMQf2U9rTwhyjKlT9LefzNz6OKJMbk+ek
hxdoevNiK7Icv8aBy09Whm+6xA5t0BKpcmu2/L71JouB3V/ID+iyDAkoikfSOBRtAn38fVkzGVwj
vDIt11+2cK1mYgvvcvTtUlMVyKxO9oXDKcdK5yfDVxQhRa58USDZ8dpz1lL++9QXNqvG+y3iLzVA
pJbSKo+wYXbCs4HMPEv7o8xVc3xX7VK9eUMg3WEoCVjGQboMMtiXiTUWEquU+TuwbsCsitfzLFG3
L5QyLnN8Y82tBmywZkQ+iqPVeaGTf70nUY3LVl+6nZAaSUkIAluMUA7ZihbVw6QR2x/xgSPi54Tk
Nw7/MdVYzVpamZR5ENsdkRmvOfMwdJxEWKdkbcunmefeNPUyDmQRHLAu+3gksjKDWZndzmprhPtR
h2bRpk/xTEvIPKbUsoi9xhl8OCwZkheVZVlMlsabQON2/Q70aOOdHCl4xzrUnMw0CZHsO1C0R/rF
Ylj91dOI9YwnAflwdwOdJDEL7iGq48wKLyJSl7r6Frhjpe7TZQQhWgLiREZ+oZ3pGFz6gLmsOcu0
9Njm4RBXEsgnsdpJ1iF2R2+U0E9G/BglbDoxC4T29eqvk5y05sHi+EbwVzIJLx9CmzNA2NH5AgxX
x/YJCEaXyXQAOB9OrC77AkTMDvAR6c6IUxjo8DPmoVNViUqYe29Mlhcqc9mqnwrUPGqqUyhKNPn2
41WynoT3x+3J+9PtR0XvbURMazuzpQdQFi2h8L9pGfPX3rlJHIFNZHGkRswBEqC37XYIN+lWObRf
blyjpc/++Y8igbxVt8BxmZJ+GgIHLKhbPz1LKj4pNnzbpA4ApJ2dPb/lujOcwjg+Xp1PN9V1ZC/6
EpBZSbT0Q4F7R7Q/ieeeuKU4yfvOtsgyOGaHmS0cBW2sNKJwRcolWEzamX86qBeDyobqVjBwfvva
qmDWuZf6iRnrRvtYw5IL2mfOBVFVcjMp7a+TF5OwPXTBk4hhqFntlLcIJohdsKmmw2qLieB53h5V
GKfhlwZkL0tEhNddB3MbfWkvwttoWKZ55Ireb2Yu3aWn8MgYv4iNgGjVVMLnCX9mGz3yv0DXShI0
ICKh1bG3Pyu/wHMVd2Rj9zgkDuQxgd6c0h/+HLSborw5/eFZkRVpaEbJrmhXAicKednXvkU4KQkf
hp1aW3XlGwisTnDqxuyOm4d/hJ9CHBCg294Tfds8JuMXjpciIx8OzeUIhkZa1Nk3JbA3EzdsaeMe
9TNK9FL4uu0dc3hAFEfdamu6/M3V6eE9hJCEZni5UZsGfmMEydUD2QVKVm86sckcb47XCeMHhdKO
WmMxG/j/EQYQ993Ut2wjtK0DwlK5k7kYEKXuJ1YddJ22+9AKDC15/R6NhQrr5ynNg5azPs/oayF1
N2282zUpeXeDJVrHNYvcUmlpGN0dszZqK+e8hBjAvbAHDa1xnIefgDaGrF1e+DXVCCHcrFvR7tEv
qfK00fP1iUYM2aOfdxodZdaQRDQk/wnm2QJ1ufVkZ7EuF78qKNY2h0cmv3RDh8AMx2KsElKMseDA
/amCBFFg/UKbfvU874iIxNumVayB4lo87w+hydT+tu5sjCXS/NiPq6F2hIKxTkmDc5gJ/J/ljGvM
++pU0k+kIiO4zz1iTwC51FnMlXTYE3maVcEDFmO6x4WmFQtF/HLK7lVmCYQUClR0boU71tXZMIxd
5bwjIZiSrJV7cZ1bJGsYSiBm0/eUUOAsQGwz2L1RKEce0hipkLYY7xEadtqVSuvcB+GwYDpt3yh9
dzYEp/G+qUmx8D9sDB9iHwsT0j1MzYWLhdGGYRzssbsNwQxmUXWNhUD9F6EHXcTHf9gxWczCCMeQ
BlfDshIj0TSCxQPhvo1Pbs7wjX/hWi78sz0Upt9PgL2/SHdjQPTdWbXMggcus5ZIMb2gBDA1MI+k
ZxU6ffZvSCUcI4hx9D4QlRN5w/RbI6M2OneFSwCsDTD2+pQrByY0XkdDt/b0Q/5FqMepUVtGD7CY
WsQPHOlnumIzcygwsSWEjk5LSyVMEyMz4pZCpw5AFodvguuN4vpPszphmKIk7zxX9Q9p1T90h0xS
ViWbgIs+2jJM2kIPBq4Gk4xGenZlHu+Mafymon+Tmy+Zc4xQWJ2m88sBIymJjqImegAi0fMI7UVe
jeudH3fATflMYAGqstK4fU9/a8ZvN+iQUnML4RpyzUXYNX5BMMkS1+2p17TNj48LttBbEhpui3lp
+yV1ctD0t6xploNjnX38B7uUx32B6Nh4H8lYJUiBpD0xEKRoqQegxtC8LJpszQxH2I/PN8Y36Dba
s5WT/7dGQjey4lX07oXHxxPfczKt6fE3zFogpskBymh9/yXYpkrRrpP0/UUJ98+F7LjZXe85+PFR
aTL6x6P2EBlLt15XPTLFFTt1tcGkYgl/QV+62Z6BNqGlRjsUB3jgT9ZtiWrR6q91u17SneW8DnYK
llMdqWNbLarOEDGWt3tQ/1DhNZpzAL7h66MsLkk/+wL/3ornkwPjy+P4vh9maVuX+buj7MRqc9VJ
JbFtxc38/DnVDnGZeujNPTfK1Zj0PlfU/BnIcle+VYxUx0SVYwHQ8tfxbahpm8irgdPhISw2R+QX
hyv7q/FJ2MaFhA43TN9mUnBOzfbcREZgIbfzDLIC3DWDSr7joRMZglkhfjoF5WmNfwxG/BszNufv
UQ4Wdswsam7mMkaC3z3lLOWZnGoDQTHKRvfk5LWWimhRji8VltIxJQ9/piMdl6M1grNztJP2oj4D
KclNnqpibKE1YvceUjkBdso6xtF4bJKyDArdWWZZnrQOYaMsz2p3OsG9OlxgC8t8N0aDuFZ6XBaB
nL8TBcqI0V5JbGEZTqLs7YyWFbGqNTOa+rFbimhDxethg9AKfsFLVdz4dgsxWXMlZFu5RJREVyyr
Ge6U+MDKGj9tdCA48Ox628R7ndXt2MBJRyapiliZ9w3yucKp8uvyX3V9EKuOu2rsmR5eCf6H7ny2
+Wm40W/is91EhBs8vZJHPP0fbzgRugS2VA+R0F1r94Fc/bpfxSqoMP0he4Y6N7AWf31nmClGNs+S
g8BXbfElmrMTU1bG4sYrQdjaEzkeBXRhvtEGKFTmgXk+6mfc363ZCI7p0nVZnEpQYpj2YE38cWZM
+9pB+JCayipOj5f/eUZpPF+7E42a2vaykc8Y8lGQw/TGZJOxYyrEV9MdXtuToD1dN1LVHohyHlAi
eRXfuuV5pVbK7siAPDL0/xVfa9FNaTeEycndshp23ROqLTbB06EElRoNxwl7T6bBucuiLTXHR7oe
a7Kl2nUAx4fm6OfdKAJkZnqNTt06W61/1hQF1W+i4xUPnd7xZ0rbNGXfprqw6FzoEk8vXQlKySgp
u903pami0R9PFGNdqHacmIU7XFYNLo3Xex+rs4BMczwvnrWX0GBoDkGVHm/oED3HlAEFdXohAMD9
OyyVz+akhoczgaqsNc1dYV0bd89Umc3K6fWqZaTwOKyFkfrSVbvQCRntimkitLgpSee1Iu8RuIlg
4NVXgML3+ZU9bA4iwRN7K3qXUHqoiDmIotankr076EPzxUgeWyEhf/40CDc5pPpuLyV9XBGr8vTb
V5f93j5Gj5U23kj1cBoNXgD7o6wTGSmLG///DlEQDPZH2GOByZXS4EbHZFg/Ms7zaF9+n962cNjk
rnBTRMr0Gv6jyGYPeG59z2bJ0CVgBURi7hFrFu9LPhq4wG0cZzqDw4a/ahAUqnU2wo3o+F6wicUE
y4J4kZiY40G0egSQhXtYqc5Vb4xyuJu8BgHqVVCQAejnryjyjEknWYHogHFEkXas5Pp9IlDVieTT
wOi7Hcs7dlX+TPTuZgTJStURCxfh7Ob/lanqMDPxdxKWKNmbVTW5AE5r1Suem8Vc8kEnoreFVYhf
DxpaQg823Ib4EuYga+CfNHlWYTyPi8J974nbQBDiXvpd81LVkp6i5CltHK91bgVRBKab4jn0Fsfo
GwsYsZi99T853JQVHnZ567mpqM/8tMa1LGb0yQgjQzvGAgApHwTPzLiYafJAhetHbpxi/fUo/I17
KzjfZsb8798FoHEFWJ4jMfn+vcw02ilgnE5cf6m+fwcliYbvPEahUxOpCyLq0dDt8GlU5PsN1ywr
QthvgbD4Ef3KOLINc1dnWZRf8pa3Bc3OXurqlOad5CdzWQg9yoh1YjgWexmHsfRhe5e+an3HtnQK
MwkMStRhImZ6R0clDgAx4ciA+134Cpsy2ZYF6eX4hnzUCdGVYa5URd6NsWizcCz60WvSdbBZX6+v
TLgQWebVahvO2j8Ng9kFA7qH9nvYZl7zwNTUV2ww2HUxH7QAC/N9Q+g2Lle341/EsOY3d1X67mJb
mA1sJDSpVAdYM9dIHGw58sL9uA7p3zV32D4nPswh8Dl9bFWv3Z02O2EsuOhwuqjRTqaD05snXchr
Mwlit6FuW7PqZcHgHCzu050SGHYLxuZ8qBlSxwzX6IkEZx8Sw2FdxT99R2ktEE/6bbikh9sIPqYT
pnKmvewOWJ6/v8hh2vgKJ/9IXljJDeZJGQt7u0hUUDgezBVaSXukwX2Fy2yQJZ3z3I74gD1O71gn
Rm1gmAPLlHiNl5PGSiwRcHlBc7gIxzr58ey2ms0ylR/l7QD5yxhwavO0qHwuKcZGox5u8bpUzyBy
2ZDH+HxctTMMeM9YRC5ClKO/a/VMuLgiu06fOaeXDSh8LV4hWcjFDMmjnziBTTUhj2cJvgLcqTQE
WbBASt+AclrH2Pc9IVOTJrILdrRDcfADKG7S9NS94Gx1V2HMXWJ3HX7d/Bh8MEB6rsJ+IZI511rc
i46bKRgPa6b6DFUcVbCH7aNFJjTxnDk/94wyHbeHAXcN8e+9CMsm40l6/j0x1hr31oG3/XnpWG7A
elAjEETLK27LjZ6QRSp2VsmVs5dth7QGstbFvCV3G7hRf73fKJMyeTxoLB+ZS4qyIhe1vfe23g/c
o8I6dKyASUBhuYy1lDqLMXxHrBj7WLlPfmeCt5nmoOhNQvvEaF/mDx7LVxZEbxr91W7PpvHUtpIT
7hbPJZahCmz2fckas3z5qO6hYDwpvLLL3f2VGFrFESbC3dY0btEapnVbTZm7U+8t1GKPXkzYJDpr
UfB0Ymm2BQ5h7eblKEr2ds9TcRT5dbWYIeoDwY437dNp2lwOqh1MOumgoQmvaSLJ4Xbe1Fohxtaq
Ik/95w8X1Qst+svxGE+nIYx6FfhMe9Smntw4wjujUwgDhagzAEA9e31rV0BOm5wze/CXqqCemgJe
B1P7jqXajvC/+0OJD3vyVt1DCHnemMB4wM6F4dbipoX8XF+tVBeyTY7yesgtvuMLyyAvIHlkyz4s
iGXxz+7QZwsWngE2oQa1l/tN/xFE/UFxtv/7xmGPv1k2X3FoK2dL98Kv/Lz6HrNYMDAzgTMAzYvp
9EqCdWlvcuaSKdgO7msGxWySqvyhBKeQyAQgOiZE+/xB5iT1p5bEVrY3y/hqvo7g+lAJ6noVnpSp
6dHAlxVrVlTlZKmuWLYwfNUdMgC0SxZMrYEr8MVmsEHW9BoD+5yXi8wXFgzgqQkVD7cDfpSEh+yI
lW0IKseL3bzf9ccLRG+1ErEQJ1xxNcvvKHyR8ftlpJBq2Dsi+8QDTxcv8OHMxl38wY3qAovrL2gx
T3lh6gPrYVx/RGt7CzIybiTRX5DWYSiOdlTGbAK2nRswI/BkV1JluRVeXVQW4aNweNXQkPEktwpm
0swpEVHDX9gz9nSNcvq+TP4TrH6p+Zp/ztkgGN+Wv5g2eoi9HAJL+kio8et9cgg819wSeMkSxBeN
pDEl0aWphnrcOsuiZBV+xxG21jwfbQ2zIS8ciPk5LJU3PAoTyhUbLu4/l8sGO7Fa9+7WRgIt7Cco
iv1JmkHGUnC3m31/zy7B9vbONblSrnhuG0XXI0VP/0UML6BPjyR05K0HHsw2eArJbPEPmJM6F27O
aXedBN6BuODVkDXFONA9TtWkf1J1bsHdpjbFAcXQgAI3BlW+lnuWikNfl9eTlxnW01oa8HhV2ifo
eZ8OHh6EkqCfIz2j6zj37C0EHflDNBqpAZ7M5EWqD2gH0k9CCZriYkJDROZzN646iwvxh2rNk+62
R6vr0GqgoJsGuBF1mzqoq+ndGO6+ebAeo5ReD1jAR9QwbUjq5PjBW9ebbEl7mT/Au74DqAljeap3
z4raXiZ6utols/Ei9JrklAt3ubIGISn2R5zFAzPs2Y+itM/YCj87Ag2NiPwtBMKK2jIQyy8KmzaR
ZsZcnRLmB6py/KMzKr9NM6thH2WyfPhTwAxfi6TSpI0gONRrRExY6DkOXUMctC+MiCFs1HbpKHQZ
mm1+ZUYQQ2F46XzNr03EVPRoirca4D5FzHvKlBtT1WvYCycJkZSVqXG61prv5FZY4BpI2471k6Pr
Byn+oxKYkUoQQ+6pkhdBGdgqANwk+DlXHtNwgmTg5K5OfQsaQvhnum5N5/ZadQGXZa1+tz3HXrFW
HxSV2IcHJTx+FbUH5c6IZZQlUkcfKcjhpe4WvXBcaOZGfmtOMIXmaUfMMsH7SZHIq7nDNfX7CAKj
YEWzj91DRR6x7nMQgIWsumBRyxS97cIyDTwYMJYxL5xN0oUhDTGp8tt6dIqEtrm58BcR46r4TOUi
PHcgmSkSSx3M+S7b4fYoV/HT0j3wC3BO8kN5x0H/TH36dr7VAlaVOUkZBjl82z+KffBCAJbWFD87
Po1EF8WOqUsnAVPY46h7vjQxuBEO2xj84IdKpmqJt0DbyXC9x1Edn7Qdt3qnfxHCUKEwMBGN6Te7
sVDV4FCB/kF0JBMY23sFOSkoOkbtQMEh+FQdyP74a0G2WGGqaTTO42YY6YC5B5X+ds0DOvjHnYB5
fCiPh8sq+8HLfd7y4zIfiLc9NoYeF0T4SuXGSoL5L1r9lwYULhhVBMLRmwFqc6oGvLyuo7/k64bE
xYr09pKSVo+08h5frRKi/pwNi7lEnEHGfTIdUw3nucJDoUnSqymRIXGjwdx3NeayYr96NjSBR0xs
Q6OTC1RKbhVAnRevOFZIMHSfZ4NrgwSKol4UjL+GyiyWP5X7bhsiI06dOL5dAXdb/gvfDSOx7bhc
j1DG5CplatW3Epf03mgatgG3NaD8y6GBQWc7W8QTlmofuTtORLVj0R9AMSQiWq+au0peIDaWB95W
YlR0YYWITiTHvgHEvopKftXKxK0hLmy3mxDw16hD4t/3wn3tMD1NSezYrHyNUJN4fTZQFEx5gouh
NovM3Ubo4bA/fOolLmHuWVkJCdr2SfSsBIKNHVfAOFvgCV+Sr4Q2a/Q0XGBTswqpo7Fb0hvGUDwq
6SKTHFR28LkNqcauE79R05T+SpUmLjZh/NbJZQwTd5YchQ1pA3a3LJsk1+annByRj2M16hrneuN0
yvs4TL8j7KWBzFRQjPGWyVlY8e+NmDXdLaDhhSdXLm0qaJbPMIP2JwFGh+sE9kMVyW4OBK+KhNEJ
7hWp3vxohvFN4lrzmNVyaoeRAYDfWTVe6OVbVwrXEIXx2xmh3TtdY7bckufdqJk+SBKoxr3sXc3L
4xGtpj2pTdf+gKYvAw4JOdBEDXP9XFxvO2ECGKdHSmA+UMFLqGWimeHBjx2mDJfHmcW/GqXt29d7
hXd3Oxug+AAqf4E7uhZAd/roKafvmh68Dja86ZSA4YeLq8YULKBmAPGLMubtZnlT9MDtrWBGR+c4
DXe4OvH8liUydaQnGPdbvU7AIOS+Wn08Lx1iHavuluy3e9w0Ng3sUu2Slfa+eedgIlrRg2kMoav4
IEt+y8YZc1uCU6XV/Dhj13P+ORJXcl5j62+9/mOD3WbM9IOs3tnvpPu/vYm/Ipok0WtjhxukN9VQ
gmsAq9ucEhHZ5dzBrf7QkdVTD5J8yRldBDYwGr5mrVY73rkWJRnV4hIYLf1zWerSLpFjkeUY3u3p
J5yhftbDOidiBATjyciU0n7MgBROQ40UOe8LNGVDexMcof17G1FbjXJBOqFBarv8X7Q89a9gV4BR
kmMvzr6HOXavcKThNR9KjvrP7lhZO+QcJQvsrFlZmyipDAjpsryGvjCmDs6QuZXOUFylps4s2+QM
sr46ltAa0T4EyonYMjz8L5Qc46qldBvtDCKqelqA//JLjo96KrSmHJgPSJSfVXPcFOiPzJSSKCnO
GWOGadVv0imGUgDiG+xelT9dr1B3c3Z2ZxxxYXWJx6kw5mvGrn5hSeOOhhhpKZaeV1Cp8fAFCnWM
bK611zCJVv68odh/aKjYBFtkzT8GZSK+uyqM/KuoojpoXbt9GVyFxwR0fC/e605WunKn9A6MxviH
wclT2GJdbWHnR8fVbXsN+BQ5fmipsfvZSIRK7wFhl5Jt7OWGo0674nieYON2uhgaW/jZqHkcS9wF
lvKiZ8hqtDaYWa56OCrYh+COqjCshAtWPXFD95kGFfPmBUZWXcsHqvaes32ueMvD5lT5ccdes16P
EHuUG58MLj/azqH2cR/P9B60vrG/lNEE23vZuJgf4KgN33KsxX/VoUmfgtoMtz3G/Me4k5OXvK73
pESKrN1pQJrqktSmnTJ45RrSAym1VoG5AAptgcahgy42VUlqZkcjtuwYdWJXLkTYfbX/UItFdfa7
6ZnsQgSPQCtLLGpJ5ZAR8ivgsRHxkQ6kq6mbvU7f8TQ+TmauKj+R2pYDqOPK1M1MzklHtRJvn964
SjosOMw9V8csuq4dC2UIIaUNpDYQkTehHCkfOczD587zpJ4eRqvoh1ME+uj+6RO9byh5wUZg59c0
eLz2ca+siDlwHurx94BmkaFGSFHEjfapvjd2RVnShiYvSAJO4Tfn3NiCGrmX3CoHxbdgRMTfM4Kz
NDzxAYdzpNGJ1OegZw9ZmKfVEn/hlQxat7kCs09GbMdNLUEH3Q4ZVjsQc8xhhNrObyT6Eu/N2eIz
L71szfhGTVbA5aXYh526vpR8GIioIvXM7vi7V6OFYcm76K4/+E+I+4wtt3WDUAARdr7PxfWtYAak
KNwzcOzex/f2w+3sLk2KkcmaR8WiCscZCvw9oTaLfRbvnwEKb31BkTdLgwuwc+oEkl24syLh6ls2
wIDdu2PPTSKuL04BfMuNR5NypWpolFP7Jn5eIJEWIVmoanHnrGZ+Zokx0OG5ZdjKxPhRygGgszMl
NGLs0dFQskPiczJKLlVTI2NHk6f9i60l7/NsQNEhNSmkmKB5cu+erqn3qcajw0KL0k1EFpxOtM/n
5qrelZfUzEbYeNzcvfPhiDO0NgiI3nDhxFfgmcrsEf87gYudyY9JOUtc7c6mnj4UHxWt7w+z5pPe
uxOLMpsAk4+KiBtqkJEqT6u7NZD2wIQeYH1PaCQqblI7nOQoIIIMFhxRq+AnLLg0yLbe2aY6QYMi
Z0LTDl+j3a2pB6RYhRoO3limK8TO9IvuStHfmQ3K74Qm8dgMQKseRCU56MtfKOC2WNIuEygvmp5T
Bpc4vN+dHQPk9xuP5fWfpjhyWtZwFbZa0LZbdvdYecIwcWi5UG4rOXmG82nbWnUFK9CB1P1RMTd3
CF2cMwjmiGLJJ0NCm73U9mXJ+jIAfIVyoGXCaAtrha9/jeM1vCvOfXPaWNlRFk6dDnmzrVaUuW2k
2LN2F2VFIh7jeHmmdaWAdh5dOwvrt2FkZUs55z6dZp4LfkCnoxNBI0TK5ceJPB/S/84w75yUtsae
4wZhojgefGa0mDguOzH+CnBJaoimAQSZVRm12wIhzoeoihYDsRalI/FsI0rNd/v1X5N6smn/+mfh
MFUZHA1tgRahnW5zFRNMy5evrZOtzE2wqlCb2YoeS6/xT3bYyhblrtegJHGzmlSPm2KVzcUJnmJQ
Yun8TW7/e1q4biHoPU2jEH3llCaGlqHO2nSs9puOlY8w2Fqpfm4E/iHHcSRGG30ssf0CZTM9ouf2
ZqfwYnZksSIXd1p4a/pGGnr3LFKfa8l0gu+9x3fVf803V820xnfrT9GRioaaycI4O7x7L/V/s+iE
mGrmaRsN3ZfGESt1PjSEvdaMUK5M208z2z8eOYDcDBLjWFvuAfOvEW8uG+ZENtSOT7s3K+tAalqf
RGIHNjhXGG03rGHonHdm86hnRKL1KgGsP2iHEv8BH0T2SU7IVCn+DpVruzqcbid19rnvrcBOOC33
y7OPqGnargJ82xpHqNWdUC0x+fHWf7lN8q2kccn/AtY1wwXVSBZmgO7OUvOgvM7Ykw5xg9YwT4bu
iOv05w1fV9KB1VMLlxHZiBC54kKxMGaLUYoadM+pg2oDakSoQjZLVRbTYbt7gxBqT9BEE5PWgWoD
pOHYpvvq7l7w9TgYTm1jPxz7RZSvxfgaGeka556Rsm7kunsFaMqE92B0APsGRRb4BN2rqB8kTuGP
4JPR6UJ0XP1xzyOefE58a0eyJQq75n6U+dxS8S7htHeYQsAwf9r0Zoyf2gb4vi2uKmNn5O6czefF
MLMgnQglqbn5Fqi8xb1q3auhbyFwAhHi3J7Pm1AC9gB/QVWDFtplO+YQ8rFJteoplgJpWnofcuTI
v4/MwLkOwufMJtLwtBgeLMYbaImx4Q/MJ8rrJnw07i/UNPX5N+NmIoAFztRTylpYg/VMmMm5jYYo
sx0oJ1gWiH3pa5/GAI0Iu8QQfkFCwAWvzfCuV1Xg+Dwitn4joSMUUcrh3B6vl11QasMcXCV/lfE6
rEyVa0DSRLGhOydo4evpLT9/msyd08KgvbyoUvD2Jci/I4Xi3Af5YiT+o3IyP4Er82FsF9Q4GtRm
aZnoDRz0C/STpXU2jvEID7x7bDjMwSSzteIKMyMwz3eSTghfkbB37JCZYQrqTc1gIre39phfP7ij
aRmNug3TQJ9EVcHWAdoDQMCxNepmjgPJmKGzS/GL1lwi4xeH5xar7djsWYc1nm0dyr/9eKRs/ry5
R4YTXSUpehp0br1cuPjS2O6sm7h/q3PYa5KMRUkOnFPwdIKO1Uub+Jv0UKaDBSM8hezVSa+lwhDC
GLgsQwreNRK5CeWjzYhqnO5UR7ue+u4B2iIDHfx5kyV6obwkqKduRsx/Y4vYdF1Q2QFGslKXd4/x
I74lmc+f/aEz3FlK42e7f/w1KvscCEbU56r2XlQz/KCn7I//u1C2pFLKoLumHFLadRcytzwspMMP
HoFJYtexPeO4YaLvx/sTdtUBgsWefLbMVbEtJKHNFST1nhqXC1kw0GcYV502nWJ/q64LjN/bYEfi
jNsxvxM5tJlOt+LtEz8BJUZGQbLDPvpySIkWoz5Qu25GNRkksMOV0k8wF3WrEcy88JrDblddDsz7
geFVv4DcvPdjEjRRozdrCNuvfsxn4RElnzcQzqcKMS3Y1WMmxD1q0jKdN6OgYiwGUbBxln1/59FH
+SQQrKWdoKWHazZY8PR6xZDo4xqXkoFc5dAN39EddD93bfcA14s9aWCKDRnIAnlHkVNaHcJWCZig
cAsM4BvGjD2gVl04wa3MSs4FudPA5aw7kyWeSfLjoSZVG6XkTxyDZmXO5iq2dxvtD0NgejZGQvu0
7t6+52Ad26KhMNEDW35VlpnXJbsTl4BxXv5Cep3vktapypnCF5788E+5vYqkzCpDgbWqRW59yfn9
Ll2f4Qdfr7xyrLA+BeBC9ETwfsW8einPWjUTevf0IxC5w1wbdVWuB23tgerz2bAt/fjaghHEWZEL
7/vASKEn3lPUvum64CLmc9fQpsWxfc+we7bGLRHE65dkBtnKt70imNrDgmI561DZWO0x2lTr8tJa
n59TB/WWwBuD+oQNt4JFGpSRg5B4i1RYDk1hIsSd0YosPl5NC0nKnFV0+chbibbBy5tbL1EBswrg
4J12PCvbSNRibqKHjf3ReJWoFEwm8xS0RyhBPY0E91thII2iFVOaDxTh8Avyl4ZQSE110y4QJmQu
quVu5QS9//v0WGPbnfp5KmqE44xCknNilYttnhZArk5uIqf2XZot/6MZVGsBtRvsDuzOi4fk9CFR
0uWWi1iCfNEC3+KdJ9pUEje4Uc6sh95REOynDymVGdtnmSlyP3ti43pdMEzlRE/BxahU/M7N80ri
w+fNq3AiSJgBMPz3+kVY+giCkE0BGNyYTlWwGvs1fJw64oH8UQZ73v55Q2Hg7wuCXrQAmuPLLiW1
FkrDyTHtpmTBO8m/5gRSjNFDiOD9GwxkRzVOo23yR8vQDfEFxQMtjgrXjRHC6+T00DFQ1Ktd/NVg
UUQcZeCmnBTOz5UUUkuV9RrRd2g4sf3SUqcMmSO7auBj8i/geFublpsq4TEkjluy2K7MTuVo812p
zLYabReRzfXs6wJ8o3JBeFZU8268irGcx/wMpeiHwcV8NV1+VgbGLMHxVLr5ajjQRAn6YZBi0ttb
N2zCg8cK/f6uwTg8MI3DVn9chAHcxeexwEsycOROem6WthDlTum53g5ude81r3QekwxirCVwa77w
5ao9nk4f7aJD4ygvdk0L1x4rASYxGo3UdwLbnjfvCfDpJULxpsrSyYkMO5uPUIFDpMjMtgI7UPiK
2Dz6apAZRpsDkjLCUMoj8v8WSJYRSsakRD0EzhviaOMd6tG3vlqOq4IlpjY9Je/1B2VQpvGeB9DD
V+XC5BcaS6cPicIaqBoBQIMVx9RKcfr9b5IaLK1UutffThTNICaCVD83qT5Zg00vOgup6ep+rZ/e
nG+ML3HvHe4/kCq4Rk47dRbxhBFZXDU/fNYiKUOkzDwfsBWZoBDf/5z0cX80bart1Uze3RvmRF1K
3u3uvm3hvOAlJbKzmFcK3pNNbBFk1qSL11hbwIe3EevLq3ArxXGiXhldD/kLAFkEx0cQWVKZC4Rs
ClytCjdHRzc5OjmG6UTBxkNNwhGVWyRZkxzF1cxsmB4w37IJ4oCTpAq8AIs3p3OCrFVOwyhpXHkU
1M+WhrS51yoN2BUoI9DfrLQYnkI3wJ21oBiGZlIhTvdgN7aH7oyV7fWySyPkx72Fv+eKvUfwc6nt
+xnVlHaYAq52YWs73lQ1IElxadoFZ97khX0hp14j2SBhygrBhH1cx94WQEchV0NnMFOq9ijUFilb
yxuUsnW8ksAUUAgzQhMVy7RryWSPuj8OHdOb+jvGDEamNn1HQRfmZ0m116mYSLtlBCH/fr/Tvs4n
s6CiIwEXHnkakPxr5Rp2ODB15jIY8MXKFM5Jq6Rq1M91bD9Qw0KVTRvNRD2BiVh6Cjnwj5ES0w56
HH9kio7+q007ygdnmeuaMx62mLkeTEKGDCliZbW1+q7V1eOWBCgFMdCiAMeEbJs8k6ZLCGK/Iomv
09iWME7hcNkwjnCkDMJdcWcGaBbIH/lpzrvrnTWzB8DxCEffJsdus7sMUwIUe+8D2eZlgCEjS6Lm
pqS3NNZJdhKnDOkW23mblk9yLavoJivt5Lii2JZpfpFWBzTpmkLWj3AXK9ZYPLXr7EtYDszfxqcA
RQ5V2K0CzIGrav0lRkp03PD1haJ5748hGkunhzt0RXLC1HjyzKf1KjGwaDWJKwOMYoCUhdB58ZlJ
4EvPN31lzxP+SeFOgLLlC8Y6cAq5a34XxSb95HhVi330zrxdj3Emwjmj2QDYNZWbGvB7OfcwsO5S
682lwOMycI78wrTambJRGkKhj+0gcFu6elqVN37PZIspRHL4ybqbRS7J0g06yIgUspnNT+HqCTle
i+du8MgkkBWCTxJVLfYq/WZPX6MdOiIsONcJB3m9rFmLV5C2O51IVrVGcl7txMU0HNAiYROx0EBZ
Q0HU5EzhSRntNFkGgacmS3+FGBiD6IUYtr+QuyWoh38mfgfCovaicRB3mYJjvDJMuXa2CQvjHtlp
djdVCQSUDBmEg5kwMuaXwuklDaC7v1H4OVA0anE42LrMl8VbhzRTJnvZqYiWMVwq9Xh9xWYy/kRJ
k3ogwJjwBBqhR5TT0fAeleG8kTTea5EOUbdw2PjGW6wlOhKFbm8IfnDYY50YTas8pMialuvFRJd9
TVwVNrGgcvjynBVDKkZFb+idLcFxk9tA6zRAtkBgiEulUtQW+JSRouUUkq1rcVO8G+RJdD13NrWk
g6ohx40+j8hXuBsp263Fpc8Bh82T6E/hqInfteG//8IbQ+A/si3IWUjMe1UVTVQ+3CW5Ov5eAWXT
75fSap3Phoz+rI/Vxt7apzZaib+mV6/bSFXPxp+kfI/DOf4O29e2R+ZrKMpgiMGe2QkZMjiUy4hV
pPRmjFuonRfRNTBC0Le3vQ/PrD/dE6PN33RXcwmUf7PkIUiP2kIfer7KpUMArShyEoOr0qS7jTT5
33TiI54OypIVs4fQqKSaJLmedLMrdwkqBbhw4Jrhlshx3BYBh4REGiGilcn54yWDD87PHmuo0kje
UR8PkIiIwAKg9fBgJ3ICal/YYthB4FuVfYHfRnVQb0GfrUqKB1ViNPg1vi6H40197J2IcAVKQonI
NUoBK9mYgKj5A9gyL+pqf1iZ7iYRNRGfWcFtjvRljAbfqIx6MFZslW3mPCKaPpLvxkZYXIwSLbTq
B/x28AP6rzeS0K2CA0+ndQgS/Gs2lkSVKJrfSLB2rsPijyESrMLim36quGy08vf+gDEQpZvf9ze9
IUjZqAPgAtuLJL6u9a9U7qNdQveXjhxEpidEq8yXknv2rzKZWC+JxptO50fSAPPeDVDkLILL/lOz
fuLKKPTkaoB3boNuglU14OdjkjReUgbOw9R8cwxgNd3EQT8CHvVcmBNryxK3X6QI70FtS+QhlaKm
MroRhSv3chQWdfzoAzS/zWezSt+WzpNdB9IKvWARi2aJhTSBOyuNsKnRPRt88OjZK0IBXlrBkgLQ
1JrCDpa/6egeekaqbA33sNbJabN27O16bHVwiNCafTIhY4wK0yQ/mKD59kgilOgJK/OAaeTJHo3H
YYOKEzy1lAGHpVdJwM27C8g1Uy183/N6Ur90WvfQdv3jlk3zrvva1OrfaAGGxEyZxx9mw2+3Pg8G
EBMsllNIn9dzvpnYH6YPU4gkmMIntZ0EZ7TUgaOf7jTL2JYH/6ehNzYxdRV09gRBuE6uiySsOdpK
79bO5xdOeGJxxYuawim32Pudh9KhdIPrYJ2W5dVNBxqbo4mT00tY1Vk4RopnsOfZJuHG7kVAOHWx
ah/B9dJXsvBfk6Y8hbhozt6kkWDn0JaoBwFW1u7IgCgrI+zfxLVAxE38IsgQTfSLr2S6uNYjitXl
pgwBxQAYenYRhM5oQnZkOJuqrjByUpwnZ/oewWpcwDde6PYblkpcenKCYZqizxns9NYGvd/GcjlX
mncH/gTLn9mfEXIch0+biW/EZDk3tVDP5WoQgQLrTfUcAMEJp1tu1mBhfU0Pg9kj+LfLbeg4Wghk
I7m6sur9DopvMalGp5OIMnwdRLZjZtl0I+pVDhBSzLAAdGlVqENMpRWfbhgyJtM9gj6fxFoPaDzh
jnqztewprABscIXa8ktf27M7cRPn8fol/8qNd11RsABcLahqAgY8uEJT/EBIdG0lhONctEVCwQoC
Fg0cGN44w9Du0LlKUyx8LMrOxLTDkJfVep11CGGAsdyEZToHFHtjIy3bMHVb/7BVral3yKxctE/J
HOhqSSJKA0Xn+8H9LQ9aGJ84gEaE3ZQCJy+6ergo5bxqAzWJYg1YfYxsG/aJuvmxyk8AcVXJOVFd
3e547AhgkUiNkGSXsg/IgXKEvZRxjkh10DB42Kua1Dpt132t+Yn/MzAtOoDW5vl69LZ4tErfwdZi
z3+DMDmgJKsDy9NVZDNdm6zCeQvx+kPJ+yw2j6FfEVOYs7lsjtcJ5wHk1fLSIlwMm8tjbEaqIgeS
J8vMWk0JoT5B/dv8/qH+ghJjpxPZ+1wVJLSgXIYoEdeKUt0okHROBdeSAk3EvRTG8r4lx9EkFfPI
Dor/1iZFrthFynvvduROUURPiMMsg5ml7Zn91LA7ZghC9wHErJ/pl9ZhZndzItk5O/46idA57akZ
G8NOcBxnUjHvRe49vLjGZPv55yJC+kt5hKJ1sNetKSxYrpCs+oZSUfuGZY95wmVgvSyybDfx8NsC
2ec7tXh1dmrIz99KOKUsik8G7ayhiWbkQ4/QDpYDFjwX47NoNQyVx98cvdkp2g+WkPL9AndEehhA
lbfKFgwlac6USz6wcA7GDz26uzWnxQDtWRoXfIwZaQE2tq/vGWcTRMbeMVt7xD6XHxrsNlHLBPa/
tSojpvN66mkeRrhvznvT2wQDu0IqJGgehUGTZyNIWp50dCy5q5anprNmmicakBs7L7yK6FryfX52
rP37g5XyoBHCA/WctH+fwRd5C8HJ0UfCDwsN7WOrQD9CUH5em+TaxO3F59ltPpOQom+O7MIfFq93
lfpUOchUnOEr79egkQcvxOeEaWW96jwlo96MTpu6NloHxWoAHWw+ljQHvF7meQKCCvXzXTAamKw4
8T4uzWXepkxdHKJkysdR3Gz9TGBtzf1LJiu0sUtHV+qEEcVqEx6yW7rRrgD3d9rh/vEBWy83dJB1
Xt9CMQnB66JexgBipaY4jZPBTLMGTR6HgAM9S6+wTq/i1Wk+NObHtMP155r9Gvxhe/iIs04n0PiG
9oCVdJJGX2REwilSeTUCRyx7Uhs7HXo9yNKNyiEpNS3H7rRM1mFJViIiMjh+Fkdg9VzSLGTZAOn7
j7M+CV+UgD4vC95/GiptYH+58XkEBJXNnZ1V1B/vcU2HTM0vV4AmqO0iMzL6pDTVDfzvAnN8l/wt
g1qdEAgnH1eNfc8AY+HC2AZvkI856/TnGgVi4V1YH4tMq9d1HA41RGfdtrC3WfeyrNrSumx3zPUw
Vb7nkQBXRVlgQg5vYGXRI04dFB2O2xJGzYmfOBoe7VMVfVwu5IqW8UplZBVHk1gf8u/CR201ME5P
I1XxnfqPc1gMO71EIGfWofHKL3DOrI5LmE8aKby0x//WU501oeVuusWPIm8qprBW2tPy4tYpXmDJ
Ss2HUSh+95KHGYcNm+BIYBE18D2ehWqmiI23TgABKCvy+MUEPmOGZhMT0S6GWwNbK8njy6PRfa8j
JMHyc5F5E11Id1iKL+cIhkOgxXyi4UPIlU5U9KWgc7t9COfulqAMKiMNSDdjXW0V8gYso9djQcDB
aCSrd1pf2n2zH7BiDi4+RCCklCVwLqVA5+kSLlC1j7BQlnZCxvD8JcuhXR26Ys9u4/QaoNWFGIq9
BYbTs50KBefgxN8o0AZZT9BJU2EyvPcE9HHlwp92LEQMSe7WCdg3V4DSeabNqYO8+vT2xovCDN+A
QRuqZc0d2l2LTqQE5BABsxm2c/Dfen+gmsWKUQ92mnoqrynJWCFy29fBL4UKoPaGKxS1ZPDnY0F7
EoAjuAWUNRX6v3sUfD+1J0d83rc7h+YONT0uYV1RZVLxbnFUI04fQRJOF6jOpqwhG0zgJKkkVIv8
wsJwTUHUpg4AIZHTCinO42QfZRaBHGlGPeVgSHNWB9gTRL3pigNwgb78JQzcC2BLG5MulVW9Wzjx
ioSmtdprzmZV+K4IPsYekkJ0aSfuar0WzwZrMOzvC+/7FuuGwb9oc+SLl14EkKPYDsgLJug8XVC/
gvzH8WuHJpHSgAloO55uj3l7prucqtFzYb/5aP+2uQZz1dgaNLSoi2Bj8H9XotqbEpu7cma3X/la
B5tPm06+LWQ1ICJ8lqgAMD7P8S7T/ro6SLoHEsl+jjb7kjzD0KRP7GG+KB3DTwMI2Au1uikMUlH3
f3ciIpNlOMTg1i5drYauNsNJHOCE4TG4Jjzymp3Uou9Hk+VbXK5XXoWQ63W4+z40WKz+O+u9nIYf
F1yJOX2toWttJQ9jgu5tupA/0GT6ZYVGVPQueQkW+p3smOXJHS3B8yWh3MJNTbJRmXHaO2+ONbPu
A3xIamr136gYfF6NS6/8IfNRp4Dw6oUsQZxcJGPb1ylfBey6T0ide+2yw1+EQbazvPivUsDBg4W7
QfI2HZ0Y+BtkKLoTKY+8Pu005Makuz//RtH2cVP5O5yjZHB7XDcesR8TSQo9DWi4PaE7gjl520Go
6uupL0BgrNNNheU7/H2mx3W9JLWWblkjsxEmsJI1QPxzTMKRD76a3DPriVOkUgiIgmGUJhYo94Ji
n0VfMkdM2Y8A99GBohs+GJuTtJVxsdgHFR7eHfQF2kGKYilysNbu+L2i7ZY4XkHxM5AZUkcqGgN6
+JwlI4Bf73VMrnMlXqGU5EeEUNcJr/9yC6Rl8/5oymzVwfhHG8/5g4JZ75syGkmasDdTcWEDBsCA
tAn5+JmTJBzZMVIDO3DzWijdIMmIEyRyyJ26ZUsSX1fwTB13cQQsSSHaALXyi1phdvxciqmxXj34
utVgCgHeyKKRWlAP1gD2UuLUnsiSymVvJF9RDS/QH7enlQ0EN8U6gwxNJbG1YGHJSO6dzZI6iwOM
ZjcUfb53ikTFv+UlC+Ji/ffud2XMWkhB7YM6SbJYsZopQKRskF4srB4MqFyARPd1btlWnaHiq2P9
7aqgSJr8TPgcCnZQZM+V7lJb/ZhHZCdN9/kwcX2E3F9m8ePMElbYQm870NnUZDb5Q2jC7wK52hVd
gobomh2kp2z5aToVQojKyu9BhW4HpGKvahQ/9qPntYNxJwnmXmrPzkaDr0f7R6p7rrSiccNZWdZe
lcRXAj4R76TlCYzbTLAdgxC61t1SSHlzB5vejwvVOsPDyKeASCCYL3LnqGj3x784G6i1BAGbK68n
xH/bZZOpa7iS/lqjzMmuud1yNvOB3danMB38enL0hM1JH27o7mZffauxyG5BebaqK7NTJfzuLbjD
Nxb8kUFHzz6QtVtsHBAnCp2nPy+ZTxWp2KW61WxBqf+SphTS82/pt9xeGnPVzNR9E55EpAQ/d/5o
mxC9xhCeG0eA/+u05iEhBzLUAmSjWQtZLtfVw1bFRd/rjMN6VpolohW3NReAE7dKt2NdQ8rbgWUu
YIZUsk1l8/mAXazqrfjCKOSewrvN87+0dPwOYyNd1iBFcByNujMKP5Wjg3uNJrE7kcbTSlmKgjwp
oy7JxH8OUWdIlrlbbpqNuGmAw6y46AH/vUa+xyZnZH9TJUMn5eIDV3SBsemsltHK02h53Vz4OUjK
0mH8tX9nv8KBEzGMvVupRoRfjImgN7wEIknmId9xIBqNUuDJmtdreV2y0yWYPydO8+AXz7emHT05
Kb/AiPy3vMgyhKlsD3E3z3oWiWLELuu5qfjNepzsazfbbqtP6b3lXZ94IXd+niDQsLAhNR0kjy6A
ynJeWNpBhmT4GXSLU3uF1/A/+/YSHLzEpmxj12JchwHu296cFmg6q/5doF3Gh9AOhp+oM9Afe6/E
7ZcSSFxUUNiizKJ8MKD/YVpFJU3mdB/+OC9oG0TJbMDq8mSoZ8dJpyPjQ7T5Wt5r2k1UybHtAzem
6o3P0JKhKYWeokiLmDOlGqfTz1hP2/AbJXj4AmlouCBcMMF0TxbBp7LFnp+JZ6UyyRMtwBDEN9V5
tgx+aUlAqQyGHUExfYOnbVSlzxBbii1is65BKkhPWm7EblVYprh5kpPDoz2ljBnEGcpde9mBCxWs
wHeeyRLVBFgIJpKRrM/3If1dK9ZTKN+wuaQ+fIp4Xht9COC0FcGer8nHHlNG4QSQZPcM2o5yeMHN
Lo2uu/5j+iYMgxFVVofHYppMd3rnZrG+cvLH7nhUZxN/YhzkhZir1ZAEprFL4RWR1qX8B4DNFVQg
VNtGfN3De2CETxWAxoxjVr+v08NyYIAH+eSqcd3CIJ5u+tHTGIs16DfQfyLbFNfk8Id16UonTxns
t8EEMyYMHHN0XgHkDqyJPwKm3A7+hnhdlOSs2cbYGhhqWzFu67zU+us8Dzx5YptnTTJ0uuvzNbaO
sBjhhakpsULoqpJURlsEF+RJcFntpFrXo+FbM6uqVNzqv/nm2kHORhjHc8x5tKWeKC8qF657NBcc
XqrrxQA5jq+EszbILK+FCTBf3w+ZQgFs1fjoAgD2MorNWnwSkP2e6gNbUGshC32ohYM8a837x+ss
atgZFnOsXl0QvAPU0zwvNWQKWgJMqSsJhzroQSeSDfw0Eq7uw4AcdIxm93+C0lGVjFl6xOMAdSdS
LNWtffEX0Fvr74hmpTF+rR3/C/rHMqMwzbFbTrw3nib6Vtx44gIXSCFso1i1kKesTNxDcWnGztuw
hlpqZdUPRIloCBVKUhz2UDC2u2BvnrMbDForMqY0HkozSXJNrR6ZqEQfiSIuFs8IpV/CYFq66Vlf
9UTfNeUsvQqzJJ/+D6BiA61Z1v8L25mEjzQRnF+eV5X4VfOY7KSxuKorspeX1cilInqL5GzYL4vj
YEj38tO3Il8SPcVHaLjhDvoLyy6scqvmG3kutUCZQGUqJqevyFQcHmMVzOc5aO71loHo+9QV0o2i
yFrUBYonSvnyamCEnkjlGYXTX8WEJLrIc7a9gVOFuSo/nFiq1NS9txZy7Auo7DRGtXtQdcvJwHd8
EgPAZIWKuRxsEeCzfjrnyRaVfnEXPZevEcZtrEpGNN+GcxuWUXrDHtmFmsIPXDxP5fEQlFtpSHmP
vUUCyC0jaIr/UgYZ9UftHkAjXBlDzzhItYLbLkjlP+amvOJ/JbX4pdqYzDfz1zjZW+jNiKARM0AI
BpVDozmTtzSiWJf3P4ep/t5rsl/scaAXaCsAEc+goLjQ330T+uWI6eR4pAFBLQaZLne58QlkNmwN
LsdrIYYMvmuVJdSMOhoev6nsLFY+Z+h/K5F63N5j4aRQ1czRsdkUqyo+dC+ZGIdNWpHxxPN854UD
qRqJb5tKvyqgk5o0csXky+2FY9dyZchea7mAEeADyW9SMhgYxciAAQn7mb3N/43pPQDcCSkt9nds
ZulDvvhv1omOCgOasA44XljLzvZyoPS6vq8zCWmIIpq6lFKVwGu+dMTFi02Bwe/Ys9hVITYazNj0
o5tEiUqEPmrcwq/eFBaZmOojiFOSndSnHIEA+PqZJimVyQtKajjrcQmdx+JXs2NtayFRLpZf3ROm
++xlAih2EQksLIzsltKWUEqpDglFjkyy3YWb3L5OmNI0QDF1JO6DSLGL1lfbYEjfIWNDbLALrURm
GAIVmezCxu43PUT1uMLDmVHoYx9CvmLZLpGrkqcby8KaquB5aivZ6ODb/J5b839FfCxwyOVoROow
69YNckxmtZvbQvgVbmT+mzgXz5M6o70B6kvEh998jktaCWgTL0J4RiUo0BWDWsYnNaMHlf5vnbfL
r+FtuotKb9jOFEektyPRoLlDI8uyBmXD3u7TaDnkolaWdhAlpImw+1RpwFSc3zhdtiQ+iMNaXymm
XyxZv23WToRhben1gvrJ3tJLVI8asLuOuNeQ9O6P+Yhavnn5AijFGiAC+sVZL8MENxLxCGXQ6+Q/
v3LqtDmV4h39qrDy3QnqOGlUpOlACkiYsO60MQTCwmmR0TSD5Ur9/4XrQGjnacHzSvRgz+AkRF4X
QK0e2q3GE2MhK2E7xl+hkVTDAFth7SsYqESmxtZ5skWRUNTAXV/5zO4MCLwL6k3IHUCN2voIUEZl
+ypjiCLHZNkoIks+HUSdNfraixZ9Guoiz9zn17wph2Peq4SaxjiTd7a4YIFcx+AVMiEmZN3IsI+r
lHZO1OnUNI+EIuA1EE0tsXgrhdD3Og77bWWbp4BiFEAMsjwRfSsiEkAaRB2uBycu7HdN8aVn0ciD
lqxQhLaXixZkEE3c556gmAJruwJiUDBGlgNnYBk45h+DRhXUsuOPFq9Je/RxNFRDKPZgbDzxuv1M
WpD6FzMI1QvgoVye5LK9svB6NoZ3YHydC1955iQOe63uoi2PaT+NDbRMZdDkEuDPLrPG1DBpn+QE
+uQaTGnc0lBKZFxbWuhavm33MYDzdwWTVtpMuy22tqNuJL9EyjuFzS9KR5rcISwjzUe7aqBmjB/w
UcAFxtoUz/olnB+M+mQCPv9FfykcqY0bIT4lO7AASjET7mCHw06UwtW/qIIkTM72JXDBi+Hvo4qP
vnwR77PCRuQebOxiBqBykU26VcUsNpIgOz6H0dA16VYryp2mn1tTp9ElRIrEmvLRrzflcuIanNaw
sH2sBIi3BI4BLgn8EhAOZtcGmippZW1PYfA6yyvwbuIK927/2V76ig0dBS8nSot9BXM+xBrkGjnZ
yvO5neKO3N1UMhgYFAubeBJImyjE+NFhWX2XX6bWWcw+qqDQVoajxtnToB6nLUujNpfMVIcDGIMU
AfRakIpaAS4oW7DGzjklyGj+px8zZ4VZRVWa29jVmpxUSezB6oc5XU3q+FzMsVcLmWdJJYayhsHT
uaoRP9GMg1jbKlyuhlnbUXEBnXOiNm+MYuFA+MiIaAcBtMB7BWRC3iQ/xoeKBWmZL0kCmHuP+RjB
spC1arXOKtv6RS45268Lrjxw/3qMuh4Glij5Hp5mmXPsJ59D9wme/W/q4HoSjCmKuHTronpFzN9V
lPiah0ZedcTAEUp8EvPa+N8VG/cAd0RSMt0RxZgeV9YSlqfr00kttjsKxou+WuOfqwwrj9PgOl2t
XiH32BJZ3itbAELSvnyg0jD3LugneSXsm4hodHblBOmxgCyDTBrQf3QcQWmyroR+MGnJJnvis6yP
0N1AGdghobSftaoXfg5gV4WoBUUF4rbuimiADg9rHturzGoh6Z4Cs3XxWa1tNF4sj6P3vHKIqG74
bG8UniMCiIvDmAm6MSZbaZCMwNGPEoTsxP35pCbYd+zXfhvR15lk1lYHokwrC1UVA+9qco8/pxOL
1l1ELM/73ix1QtTliUbxA0/HCGcpiIGtO8CpxGpIfuv/3uUwhSuDr1IQJK+C6ndLHwFKCUo9IRWW
m8WAb65PmqUIRRxPMNx2UkWWxqWDGq+i/OI6bOnDX2dkhrXlLDpZUrfN6rqz5TWtEdXP0pg5tWeq
DbSdcGdSACLT9HCWt/I51O+8gxZ0INeF4rVY4+q4bqLJFG3UaeZnCsqi8PAAXxbwlbAlSIjeA5Kk
DyVgpJrQeWFdtQxbwfZcaOyqEYVUZew+ZWCKSnnH6j3FHYWkBfnBu74EMmXBXX9Smw1fiALHwuQy
lqri9HFapRJyzwgbCni/cYJhoxfAHfyz9DMjMFM1YbxzzxqNWy3occcgnQkSSv0sl/4yX0vPchmK
z+ekorVOorWr1T5G3fEQ/uqSC0+UfJxc9WrAmK5BGi9MoCYT09xv+9A5wae9mHiYsoPfM4IKx3WU
40Uqrk02Qofb13ylvll5epS/0uOj4jr6WFm6DVi3Uxj42SrAzMkScemdaSaTGlPGMfK8RPCE/88m
rtAq0IhFLyshxb1s+Hygbi4lUUiNHfyntB/W/j3N0nJpSKyt+soUHXV+5y3/EWHYwSAmmBgoYeIA
FcKpnIgssm/6jc3Xf6K6NvcErxbsAm0c5DKkPLy/s1th1PM9HZtZ0QsnuqVB+sTZMNcsmbnrHysi
4ElzsBPePwtKPNHYP94pgCBYcw6MHOx5K5O5CuYLuIX8obQ+pqreg268StGszMQ0KXG4j0cT4zOd
ZpjR0rOlLxTahE6sTgULp0bBe5P1TEsjVFBg4WaElOiDJ5yGNCirZVFdg6sFiNfWKp8Hs613EUER
buA78GXuYOY3Ebx3wb1xX6fiMKAj3M5MnV2D85/wqUxWiQe8m/Hx4iYaSnS2KX3m8ZaLEiI/Ltns
eWFuwMBNK/zZOPLuH3RLBIgn6z3hQPIL7zeb6SghMIu6tCpEMVyMTa6JG0KxUcMQqj+ugLuVPqMv
wdNg/wYOy3e/ac3BYkI0NCoNj0yZj0F7bKijKke/dBmJF9k/8ro1U0jeHVYrVIdmkJ0DgTSxogT6
p0NISbOd9KeIBKW339eFj5p36IasSmQc6lg7Jf3kfKGtP+AaXXQ+f9iD9TsTkLtgbcVHrw+4A1MG
BYLWHz9j8/QtR0Y/+159JUsVr+DhlUdG/INxpfGatsLccwSleR+SDsXVrFfxRBdcb0OjfmMBOmbK
pVY2oRtQ9LPTK6Vn59eXvrKMhRQVrYSCoYQEqmW1p8pUZlIm2AU5Z408nYekWmCsa51ngHUzuU+p
u+o1BebjyPAix2tZ83HOW1cqQksbcJbKWCNrPwn3wd/3jbY4p3CtkZ31e7uH+mtrO8wVHaqZgod0
EGkchun+Zd7uzpE5SyfTvo4Y+XHXXqmMTgfd0opK1LWxkw3W/fh9/Yyy78G4pecCKGijlpPD6mIc
c4tLUcmG/rZioRUOdiBBO7ImDG6S9+hEWlbwy2w9P5PLNIaRSqLXx/RA3vbvTYfgEeMfFoNAisiN
1jJtBtgS41lVJ+QhIqIO+b8C6RSRG9a0xIKqgSjcDzLdL22APMZxPNhMp4og7HbJTI5bGoJzXs5m
dopbCHtQOdiwwsd4saAiBICOstjlmOEBiE7ZK4HYLz6M+RLJGFhGkEvn1RqdkPDOsHpm1USxBVGv
BzL+/UBEX3KKyjNAwmOEHvr6NHCTR/nz4B6r1cU25PFBCa7zuT0ZiBp9qqmFpy+Hgz6M0hg8sRKX
5NEGO08+BYYNl9e0xag2aYjsBI8F0BM3CpHyhE7muqZdPX8JThKFd7l8hP5M4XQ3GvHvoUqAc3rx
CwKS3VVXCVkXB4OKjQXM1A94urjEB65QbfsbQZZh3ScDsOjzCTlenUFIygww1z9T0SdKk9S89E7a
e5fC3QbQyLLyMPUz5mUWd/BN7BYMuXFdVZBEIbzDWUm2Yrhn/XNKe9jBjSZcDgIINQpyQJUfFSOt
KoVldM81Z82c8f70MOjFd+auMLZVQFpxwtWiHKbYXz8fZGo3+IcJj6hRV2GAQhhLiUUCEscSw1Rz
XhgwaQmgyXB4N+GIgOTsYZ9Z4TtkS10BczkEc/lga/jtae1jwVNuMFNMkb024VMAqmT7P8m2bPzu
q7o1kDwEomBX6A3VQP+wBbSoLkHCtrO4lqpqcopljsl9NWT4S7D7TgaiVVpZYEOnLngShpyzEd/m
KMgP/HjHLozhO/r76K2eWrNp4NU4oQ1yrIdMXruA6jEdPIblpVONRhuPaGY3OyE37QgscR8mw5yc
ob3+UfahIVXdZysfz4M6o3sz+pGjaAPSvFUCtTfZBo+aAI1d+4G2tn6MGa9BYhcfpTrkk6gu8ex5
VJToDU3o96latk+Xmlp73+ToOp9ADsB20KoDQH+RghV6zY2FchbtP8n9gun2y/12v2lJzNOc326h
1dHjk3Twt0OCxugd2zF5wYXutW0KJ87VdHFmkY+mW42WaoXjKl7PNE8WlIZ9xy7rtk447nMe4eV4
6jDo6fo5FWRYaVl9thhXCONq7p/w2vAjojagOuRL4SS0Joga3RXyQ+HuV+EKmKoXNbo/BhbTst4h
haNn46P+RTr6QEK79XTYuKfRGcO4Cu5zQeWUzjvPZhj9CdIcd9dRH4EDExgJH99G8wqV0QkoHTVR
JnHoUTWz9/zU9o2RTDX0mncmfYOlsFrnmYYr9H7PygkwtWw5yncePLctwP98Np17O+SmkpuDRh+H
ErenHxPMV1xvdPVMPFHaIa4M8X8JrJsD2tYai+rbqCFUTVVDXIk+Uwyn1ykWeTMlPACruHP6F26/
VwRaQvptLKAZRyEavgU8mlujl4F1owBrdQ8LQ8la06BY/Z2i30ZPkFBgzMSgJBfPqQEiw/96f6ao
evuA9UMawW8MQHIkT7KWlrhCcz8aKd5OUfrXHaeTWuTlX8FPG+MCQu6Cv6oRPuhPoMsS+IXR8AKn
7nocbNTWpXgOboD2HsImGYwspeBYHlU4BBNJRgaVupvAYqfBNztGC6uKhwTiYg9EyocsaEEVvSPt
481JkpNKFxS2wxKxVsZ/vdYXxkI9vEneB7b47Ocf15KxY/nlk0a9iZKDu7S3t/QsOz0++zdvwBjs
ASvwJVfHsp3zbT8If+K5zUGDVIWBvTNQIzHMUZ66bu7OAOwtkF6MSBRhXS5xLmHuaJBJ+JCBfTIh
RaldYUNfWVCfbplTVSC8gcbZ/7HFjvFxRI8dbEUnUTMGT6J7eEsAK67Yjq6XB6xCKrfGkDRUbNFp
JN5L2riDOuwo9Bq5FD9GfCwxWHYlvavmkhaBGLHsHvpByQeRIzoTUP+aai5AFl+loZQRBRFOmgN0
kX9jETi5b/TO2fm+OEKLRxfM+JmYp8dNu9D30N68xGtTUT2QxNR34tvoSWt1cfT1YFA8thYI2uVr
QNSf2iEsDbV82wt+zwLrlUL9Q6VPOhh7IwNNwMexn0othXLoK286QtDOp1lelEmII/b33EuqtNFj
wlt7WxH5UD627O1rvNeRkQKty7QthGVM1Cpw1WTwLvwt2yUTSbcslPmigg7Tmr0f+g9TFtL7GJYf
WukVsS4KPsfCyUQ5i0MCeD+Z3dZDhLgb+TOabpeax1Xh6yyOzSGJNXZth38XQs5IKquL3TsdEzit
raf2TvAIE151S58WOtuORjdVpoRzlOycVCR8Yl/EfPeoBjxnJqhiSAv8KakGiXfYRLJ4jHKAuxcS
pMVb24P8L8HOmuf3U20BxgSIw0HlRWrw1wv8y9gvqrTwdYYm99aES844jxUjy/4zE5mfx8H0JTpG
7b1PfB1YrS06iRfidbAUzNKvno/LGkSrFmkjdm4vWMPemTqU1DOre0iOqARcc6ksihImQAxT9dbp
c8hDtmwb9z0c17Nhg1xZ2wXINzTGlF8IJkVBwDW6e12DMgag89wL8Q5CiAk1fpL1uCzTYAI9Cnf6
NX0mvPXyK3+JnX0Kj9EKk0RZQAeDQlAnMjjujY+XobUw/fTNs/gVraXhIVS0cPcU9P7brPpcmbvQ
rzLQF+qzbNMUOCTNVUU8Vl7TSaZvAyYd5bsmGF6tQjwrRDmtut5xvJgesB1lmQyhT70OJStpEZwO
9so2s/WKZ201Kp7ghDPcN2R+PKFUubMlon1v6cISLqzSe+mc1dhGIOp9khk0IfSxNvGQN78TS+kP
Drp7Go8ahbLcGtMm0Z3qTDLetL/XENsniL2X1DVmNpXlwHYsl3IaqjOGrzyzBi7hxCIyROWvwdsO
ue92OLf+ChH70X03CCYk6tcGGHMzsMXLaJAnuqsScVxaqOZc5f1A4/909UzWAXreiu/R6n9t3Z+B
a2GLagYCNfZ5xvhzJBz/QXJu13u0tgvlZXO4GiXHPfmm6DQDd2u3TKivEEWaKYlK4XYqubO2+MvO
ekaoc7xPwblgZl6PHU8hPwwGmJvXhkIjkP4nBnSFzm9fM+tXh42gYaw8TneYBtqgJWqi4d9SpXQF
HVyaa8uet2bI7vOmJXDYf8h0bdAGK29mLO2NF3ZWKnyx/va0K0CTR8NZn7aqdG84OdJ8SV7afM65
oEhJYxUyiruka/nbJro/eNsSSVX/9LgWmH/szGhWXCmARBQAMeXZJL0BTpy5bBV8m1ChqlzDGBVQ
Bm40xD7xzJ2nbFuqG2tSbyad526x2KTSEi3Z9/xqaCcof2R7Ic04xYdSlIXGoUBPgs+dgaaJ1URG
BLnvIKVGEjgi0YcTBMQk7zy0rcoVMc52VRFVs4lvsoRi0aRpnce4DinSDJ97vNvYUMzDXzbzHLTS
YdNM/akTh86Y8ZUIDezSDDXnJrUUG4+92ZT6S34AT2iSb620QaQgG3r72M4kjuAoCjqeaBmA6axM
dlgBpTUfGEOpDo6Bw9eda1bBU+UZO+LZk3vs/Vea3aGCj4kHK2YUyi5sGCwkbGKGPGwf3FcLApj1
sI5OJr5BmOtJzxIzYA8hEEg32MHdbODFeGC5V0h4UTn/O/s36bAUoOvpS/2vwHdlYH+OZn12diJg
zafYfGmOs9WzDzPmkFdGrzhd/UesoE/yEVs95FoeGj3OVauPOSLoUHxprM1IfqdfWUJ/lsRZpx2o
qSxFkq1E8i+czjTMyjvjKoeR8GBi9FcFhU6OwtsG7yeXXQA/+CrKAEoKWq+gLkxJJmU7yPXgo37k
5ypzC4cQ7WqNNqafebG+ZC83vJaAsvdckP6Rq4WAW9wDnNj4eXvJolvYneY1xjll844QNs1fUdGM
8UsFsHikzaznumOHxn5LkU2J29keFOOat6n0sR5CHK5Ns/sI+3IZiWO/I363Y1+uXBxzsPDUwccO
zqvrx76a8Ok51r5ZDu9kalYwkJaSjy5L94cb2vIs+1+e5wPpIyARqZqPY5O1IPPE9wHpcDA8SI2F
PC0ShJLc47yOQrwU6pKFsiEQ8sMsXl+gnf2fDsjHv+Zl711DE8l/BjpyT9AaZO5/LopkER0Yk6YH
+MvskkViqH+jhe4Px7RapJKC6xx78WQ/H/gSuyJeiyD3tQY1kYxTde5AsQCxcoMCawdTtqO1XCQ4
X6hN2T6TvlmFjenfr+7wJG4OOc+IsvlWHsfCcnS+lNfaxNUK+s0x6dPMQ5+p00K9yEfaJeRg+WR3
qA4mbcD3yfhX4YHFNi6NhBXaWxOfui7mVTo6WoqhnMbVU3NvH+QICXKRnZxf4FfgHN+RVLBK3AGm
e74BOaJQFk+kdoOygSH73D2FTzsVvYTmhNwdwZMEVjIkqdXTvsbQ/IWdb8AZkPEl7y+EL+Ck8FcS
zniwtLTFBXWLRipJl1r1jvM8UekJae0M1GMSM+Vapzb0vVJ3txdlgTrWcAgRNaM4pNhCYe1A7Pc9
XrZ8tx4RmkUIp47nQKIhieLgqBO0u7cRynEz0/1SLmQuW77CayHiV9ZL/5O40fYVR/d3dlQ7/7ox
gVt9U0vpiV3CE3Oz0ThGHtwuPz+G/Y2pNw+D6ewA5qxuwSsgfY3kZNq0b4ex1DLP8gqIknw+YaAA
DGnyztZ4YDrEHYBmO6t/3i9ur2HIEn+++Uvtt74Dv8x2YHSs5pZyEKFU9mNrH/fpokA5lHoWeCxK
H0mtQTmhhl7QZIKpw/tWG/t6WfrYz1PzrtoDGJ9sQGYtagHPvgGactECI2TjSjVxwZhmIDRuaqPh
DlnK4HhxR1K6pFzJuNCKpe1fvB9Mg4jBgjobqY7rppBHrvvxZqNpqxMRPWRV5l1TMlJd5MB6QL3F
xAQxfgcIwxUcfyjATZaQKri0nGKanuyAwTRQvBYxpY8VhQ1hi7oXfQi2tJ4yEQ7mC8IsVsXtvZMI
gdcRHyAkyzkYBwnoewKDbLGAxtzYNPFftEkJ/528fZhaTYjtzmyYpWt3RIkyfkO/H2WAAAPQIwPc
0jS031TAD8KDpw4wpZZjzczsZFEsS+uehBtDDBRBpg+xjSztOmHao8UDFhk+ESvdgC04QPtxGIvX
airwakM2KAJBS4axVNsYHi7maiYV2+QCuYX0UEdRlwv+GY49JVBuQw7uzwvDEoPLiGU4BOEpq4mY
xesJ+83XMBHRS0ZdBjprUdM3Rj89SQG9iGxlGB1D0iT3qFSGfslLW+32bXZgxZ9heiiq6wdWw/Mj
4u9vTatwVB89hyGiAwWqx27vdHHyEd/+lP0N14S0587oGMuk2sLolTYaj70/D1VYyQvG9P3Pg6Ct
MDZ/OTIuZIJzWvU8EV/N1xu4Gjy9IFYRHshqzn99hkIDx827oD8kLIAfJoPR+NBKXQ6X/KaE6LiP
gTRGqspTebBixxH0ZPy9ZmNUCs9dvInIB0Qk13JLUXPcOABK5srOhbf7wyIKIN9/AnLGvZsAeLTH
Z+L6TEkYyOZNFYhWjUzx4dstoyq2hPCEQsUCP+BeoP4mBi+HRG9zMbRo6ZEAA7lNcOIPPp6H9dKY
yhJgoAzq9p4zhtOxBlgPVXPbacufwCAe/I2cQwkt4xgzXFyXJv4U2DBM7o2znbfgrpWtiZ2JFzgx
oYm4fnlCNMa7QAR5aWHkByDgmSxg08nBKmpLkhGKFG7TFJGu9yY86ci7OLS7Yjf3m/wAHygTB+ko
98JuYSGdnwyrmFjLsEZRznsiCtWE1IAXmHSt4YpqGTkZ0N6JAA4ctbu/k/gTNJdrO13b8YuxLWY7
TzxXocw1rF5/NJn1Xlhvf4Cq0I0U4RpEsHiKFO2+87uiyLUFIHVPxqUYM/DwTpWdHmJdnIHmiwy4
VIv9/PfonsUmEsDk33NBgaFc6bNghhpCmpWM9JnvNyBkx8R00fs7Ob0x4s50ZZz8gsafLqDVDzV5
RPpn6Kh8DGza9svlDtMHTENNnxNxqzS4CqIDH8bMZcE6r5ROuXar6NzTVfAWcwr1sgztDC8lzGKz
WeYkd27ocvsUCizT82e7g0pgYl8lriax4PeHL1Aw/RASGuZU3lGOQx6U7+r4t6g0ttm7mcrqEWcH
ulaJ4F8lQ8wC0y+5It8rI3a00SUoRoJMGuAT2uiWhC+YVxDfM/t7ETWXUz9J161rk2T92n1FOFUV
dLNC891aRxup53oooIREgE6zOzfO+jc13SeRDJoDUqSxftq/6C+gaz6MNj9i2SxEM8ujD1wN+ApL
y3viKMVq3QZe/Q3xbbYHJU/ibC7gHmpSPGBCCsylSaYHv24m2rxxtrsARzNPdssPV2B9h2Wg0CW7
lCnRQptpd3kViAeAY4TsQFW22CVEjqWmUi62wTkEYGaQhDWJb54KxBFMn8OUsHMDuiOcxzmDnRTf
lZyh4v7QTI5AxltKetMmgoqaH7aTE+8ocBvdPiNdA2AlbamomQasaqIx3foxHXileDZjJ64Vq+6r
+q51iiEAoeRJzQGLT81jcAtDiBSaT65H16sW85cB01tK3ms+my9xnNeAHBS3lBAWJ1EYi+e0ToxD
J8titmSHSVwrWbxOY0hzo3TwLdE66Pazah28qRfC11omp64RDEx04UVR0BKHgGpBZ6w500RcvJOf
/dNt1nymW8DRqI5c9KVTPjxdVqHIdpnJ7K97G8EqThy3fw4cg8/A4HeQ/tGMTxOtBoM4I4jOwEZ3
4z0tlbcSQXmftSIUm2V9ENkOwwrTPw2fiHLqr0kM1xTnpcHmfoAbmzEJxFr/zuE6Uc6zrDEALkGY
hCKbPZTNYFg4dq6v+26MiQZRabwWFrR4zcnAJfEcfVmPyOPQpJofIacLAUGzd8luV9X/czoXR9Yn
Ddz3dccuyeNFJREFnzHGQGozb6dv0fLaYW36DZqfHob6/piVT+nfLnb8v7tFfBvxMWv8tgGeuv26
x7JMhSTLkZWcGsgX96HZIKohnIz/tXH5MrS8ZkZCGNYmuqnBiUnWfmEYyYSiVTbhi/0OrSD4Zwi4
VUB7WYE5SdCxYzJn8ftQ9D6gwRM7BJdpMN8bSQ7a51KiaV/epHR+KbCKaVrHNLygXX+Df/+fEi8J
HPcgo4ciPJ9mHeSrWBSPuJzvxwyV5psucDClNO6qgfge5mv5SuALlt3pQY8HRPUZ7NBygpJtZGMK
0yOHKIs66SLO4n+BW+SekbU9lUScg5vDtU8BP5GFG9KPrcCCZRaf/fW8w4342FirnuBu+GE1Oevm
3rXw+XbJkYpwaPdHpnNbgnA0y7lay1JZDFV09rikgZXqFIroPHXqg/Q23Scq5GQmzIsyaR7dVyCm
hyCEe78PYVZ+6n9EacLHncumv8alXkiqA2CqoreLKIHAzSg2q5fQrhPpqjFZmGocoCHoiaPQamgF
k5iSWBCKWJJOaUiSpPg+jdnPt+ohOap/pjxjNxcEMDgd1YkjzktLuXwPg8R4gqGI8CxZbz2NuSoO
aBq6zzV/ggpHdCwa9CQZ8zlV4xFSWtY+MfZxSrFaWmXbN/CSTE8fkiEpUo0ehnkqFSJXu4Wp3hQF
QV/R4McPQz5xmlPHj04RoJPbg8zhkk6qN92/TG+9T9i/BPHcbK0gz479G2J8XiAsysU7Yo9hc6La
px4cMiT9oUrNaIcNqXDLJbi1Oa3VciVCSpsnmEyJG9CoZPpc8fnKvWMvWuYrZ8x860FqrhcMw5wB
cYtFQvJjIodsk/XztGj/1xB71ytqDhoLqff5z/V9ebhJKvkhaLVj3SBhQvffmilvWawR9UnSnS36
LZqNGzU8QTzSZjpq8t8GJjIrQZWWZUHr0y+N/1VkR8h/RyajaSJw9TrGzeY9c744iHLO84HrCags
gJpICnsYtkptlOwMUJHJdTBNV13lv0ikQJmsjjSqyHrpEfiXrMDjmJl/etNNeo2CtxFkGgWQJxhc
9ILgSYVhi1u5PiHbMzWHOWyko8iE42wW6rSAeKJkttGcWP01m5nGovrOXxJhrAE4PoT+iWeyqqd5
csLfXmH8ep9emCwCRipDoKhbSpa5AKKVyBq1SpdtFbmQFp1QwDHcBntyH+iZrURlXcMDRFATnPzp
aAINNXk2lpf60U7QWzSFfe4KUA0T42YaKFvhA+KsNUtmJVAury1HAOzKSzcT0WZ8sFY1p+p+9BEO
pwV9Kru4jn6DUnA8ENZu98Zu/EODB3kDaO4/DXMJ0gGbpcIOoiG68nc7pu4bWl8Nq8+vPD0I9oyb
cUD5m4COvAa60TgcWZ2jnnMeL1CLpsJxSke64H+S7T1vO6RzyBoiERl7UMBfOXH+NUDkMD9KbRIq
jnEhCnj12Q10z2IKXugxAoYWwIEK6hcaFk7qtGAiV0Ecxd6faxblUHs66Cxx+Jgt3fwrxR50sTZI
v4LVUoFVhuKvW38nTaE3sB6xCIGP12g/3Eutd+77vaMZ/4bEwVlGoxMh11WEtf+mPCLmfuiivhzf
KAXmNh3PrCLteMGXBU8chT/zsuv5J3f6lEXkhAKU7Xz0DpY820f9SyuRjI4uPbSGs969A0x0EWvT
Ws96wjf1yq7E4cuoU3DpyGYhiHe50M7ts7s5ePbvHuhCyH3cv75k+DvkojvZmKXnwMs+C/jat14U
lVSYDYbgUlitdRYw29qgOSLT0omyvcsLmSPHgariDB4FYe2FWnI5dqXmFX+g0dbE5PZVxrCFSjtv
iEfyEQcj++xWMo8TGPHWOsR++COlqlShf1qQWKg5wCsGyaZJcygFG0MI8nZzqTjQq01T/VJVUas8
G37a5m973WPudt8DMGfV312+eatr4OmfO0Po5h8g7lo6i1jIFilQhzIscxXJUPrsAlmuxcNuy7Aw
meO4kubQxN9PDcRvzQwOlZiQsML3V8rjRg3MXpZBoK55kSBgW7aORkN6zDCAf9lGTIdOB4Md3q2S
13x+bFKW5RAZVVxAOydC5sSsO5+ElSjB88vjl/ZP6np5aN6mAU1VDnUvyZzPXLmMD2ALU+Vsd3IL
R9vHHpL00Oy2gJq2pv2IENFkqKXnSCgo+otmyGPY6dULZsDi4x2rBBfsyU4pQaPgdw/Q4lie3b0d
5k04XDc0j6B7DFZ+aX81FngDTxjfxi9Mj/fRSKPlD5v6yEudRyMb2WLfotkxOHgTlR22N/uURNCV
z/ofn0uZHXvmlJAbiYPj7VGt/4/oh/uR++1vtWhOrL800mHPuDiGirhB323AgEPcPCUgJfikPL/Y
e59+djBGLaDUxpxq8htjFdhUaF9ED7KPPRa40DMBROSPrtKHecGS7Y5nKOhrcqRNCsX79Lf6ppn6
IvB8OrVFBRlPnlFg41qPMvMmfs3DQxyn25laDnvs5HA2EcPK7DvtSztGGEn5s+bMJv59qSZSa0PR
FPMIDOqEFemw+vRPjhThYjYIUMtfhtyo0TMBUWz7Ir3rTLJ/V/kvUmuy8oG39Zdnp7nBKKQtTQmf
TGGsRbHkRlmblHxqQd+P+gcn3sS8LFc20O+ToRM1BGhrgl5yhKw4uahn9sWvuDdxdS1cKylaEZJh
UJwb0rpf1TdWJbjkkhMeT2IU3C+pBwOzyG61J9Qc2fLvytN0pNZwZdnJBA8rSG+9YlnQaG9uvTz3
e3gGuNcgNyMySLnlh4K7wc9Hda98xeArRBtI1kWBcWlHa2nFmikaderhp+ivBOEfAxKdhubqjFRx
LasT1mz+rjkQLQezucupsazhylnRWp9DeNYZYeA3wUSNEQl5OF8o8tCCvHUjRQOGQPX8Ko2BsSCW
dZMbj7/OIRRwSNVA7VesU2q6YbWdcLmv9ci4JKGyr51pSEFLyw+Uuqq12bHtA8QNQYZudQtKN75t
JfjnrRiCS1133nGXY4RAs616K8ybp4/IZiPTXQM6eGOFU9aBIZKhFZqk7TYCOuLZ90S0mZQU81Ro
ejxhFSybHp/+uszk2RmI8B4VyW7u5h+SpyJyS0+DxoBjBLLpAsDs/4vixLY4Dz/vVBcBXJa6wSkW
f4jmDo+WAYIaOW8eyGon0O+S+rrrLAe7Fu30Gd2Rbh5dK6Np6ATJnuHhSYrspCxI3Xug5CzyM4Cv
hjY71riQScHncZY8AVz4znyhIoYjbIZJd7LrzeiZ7YnSaQkFJ06JruRfLp/qtCuCgpqshZED4bfE
78VcgWDynPpBgHeppVoRIbIyCYbVIPtGS0Rl7uKsQkzUv1YXXTxFHBcvrJ/k6A2wHlSiuJBhr375
3ABoTbfkhbYzlTvTCGEZ4bsnquu4Lhp5t2LfMKIEOVXas+j1jXRi2eqXYJiSqBf48cnea+3ZNVs9
xVSOXrfoqLcrWnRGtdmGJyHGunZoTbG6DKf/hjPRtdJc4fK9BOJLRSK1zwKPfKCzWCfW9V+oNS7I
k5rlBYZu7oCWgYx2RWHyuwxGLu0nvxKq/aomuAv/HR7bHIZjcDHOzmDKq1RDPJS7pjEAJFOcxRbY
suHFxYD2NMvAbZtrp+Hmntx7+6kwcE4Htffv+2loeHfidE8RmEb18iHwTQh4jYon2CMjwauzquV3
TxNDrsKhdEBOTbWl2OWsbCXH9KpiB0tXBp4Mn/dbfmXM0p2lLkg0XP1+uwhu9UsN9cLuigkZ8qrJ
S+P21XzsRDuPR/QM2SFti+Uvn7yEqsp0PlaTfKpSqBxu5FDgBmfaf7g+lz3IUDHLPXKY9ZLbnDZY
r5HnZCXLo+MUf1do6nl9zGM9YLYN6YDV4agKM4pclg3egG8qnFMIh0otR4IVFWLJMPvIMKWmltSC
0PxyvFjqFoea4M12t5fRGxmQhkI5dpjdOtu2EeOt1IRNFBoQtUNV4jihnwnOaK0jAB0S3OVDEICx
E0p/sqS29ZJ3BZ+vkEJImGUhQFZrHFrB/KdXzv8OI9ZCb4e4KkDkKUI4CQyBAgLErFQKmyhVx2WP
1CS0EQSrPXj9ZbAarqEuSJHM7/h6CDez00JpcFceUT/k3fsh6CpKsqjjUFE4qMlfdeheG6DhPseb
vrWMb8ar6L9ESDQm66rOSEHJYNR5+DVdBtSvcFbam0bb356s9LnEXC+8+aNIJ2Yx4xiwR4HMDlrZ
ECr9PsmDJNRVG99oWkir7A9CvUZUNyV6uDkplUmh4yrx3bgNL8dTdVs4kro3tg1VvkYoXUeUF4ee
eJbYeO5vzXKjgRM4VVqM4vJk6/qYxqnmr3vCyak2vJqE3ejTmqCTv0lmZo2/oJveHT4y9WljsFNz
e0L7MXbNXAn9Kd3Bp6KuNqtdNd7Hrho5pFUfjzSG++HQkyyoGFrG+MmOJNFMjorX7ho8J9v6zGOw
cVnTDzGAiJFdsDg9J1RLqaJb/jh9CmQFaC++3bKh16ouSTe65XQp4Ssr1Wew8ni5HSDAlNRBEHJ0
jFL+EPTtg+WZXpFbxlovLY81KUhGD5cAJ1tuCtdS7qx8APqfSGPMOGkjbDlA9GNlg2L0EIE+Liw+
/QyH6Pm2f4+Phc7goVujpSy0LeYm3evubKSFRqPZqS+U8zV0UEPIGAt35BCPQR2L4OM8HXNHauW4
xRGe86kJlyPOScr5WKfBSRwmOYazGZS2YfIXtkSqZZPwrfX0QxLgIY05ZdD5tVASXwYqkg7Wia+Z
HNT1mQnScyS4VBfcSoUEkuFQf1ooA5srwX2wbnAw3L8DYpEkIgMgy+qCynKRFjDJIpEUsZKStXBC
Sf6pIs0/Nz+VcL7udAZewsCFahyaFPQC9hFsJgXbHU9itob63dmsz8aOtJeGFw3ovQTvCeAitK9x
lL4YiNGP9WBjNtUBF4XFs8jH0mPV63rKNpAeE8Y1/I6JJsp1ZDTuX2n8ZZ9X9pi6sZ9fYKGoEiX7
DLXHGuZynauqJ6qrMzdmXVYKA8xIgjAUAdt5tBy7WROYSlU8UyyIQ5HjslCEKpAlL3KYaE8H8el5
7JfURiD8Ej6Hj69yo2OzCSO2gN5sbYxcZ7iAOHoTzpLrhnl+nRwzxyx/uf/1q80LXBDW+6mdeDxE
eYoPiIrYjbKRJiSvHekDUSAQJQej1joOyAOKtTSHHNrgXNf93oIl0twVrR7MwYauN2sSdHq+uZAR
8+l7lec6ErhGjZheZXtmpeV6+Y9doGzg3Bqkb/swis4sIOCXvJThSCd9UP6OePFlTzwKurVlAhqf
kCQOfWuYWVURQkeJGPf2DDq33oyKTW6bafhzqtW78hgFAma74RgnbdXNHsEGC3q5yvyTE7zDoVU1
ylwk3zxjxajP8CGXFcSQzYdj0QOsg09e6G7aG9DZ+bTmdBnk7L5t427Hb8/Hn0XxJcDiknObQWn1
bkgSA6/DUz67VSyPp47vrOgqGPc4UmgbNSlMlkC2YnTzqD681zUudy6QzLvu0wGNIkjjbDRUMik9
AdqH+HDmVC1rKIN02gySqZNWWXrwt7nyN9ltOnvrq7oZFS24yYVDg6Iq750nuVqWui4XFge/04PJ
cCjV5JG7HQewb7hWjLTW/jkFxknHjcHHyt4YoZqz4MUSFGNDOQDWfcf/j0+drkdF7U57o6+aWxyL
uTnOYmGE/wCv/1F1zAYJNwZa2PENcjY63dtTCjB5pAHjzkfcr3FO3yMBlTM04OsyDXQDq8BAEkQj
ViJagfISZsdlYUrNn51TNbdpCnn2uazQYmn/x/1zUpxy+xM9peQmlwZpB9xOEEEPqvYryeehj/TD
LmNtZIgBdGaw2IPindpADvCvj6LVefl5AxYWEM4gf1nYRorVpjsVNrKRQbLYop213FRsl0rfZU/Y
b+mfsq2ybo6vX74PsWezdOvj0D1WtOpN2/TIivR+flS2DJoPCc9pGEJo7ICOIuFLnPZ87XG44HiM
p4DvDLl6jnY76SroseDGBfLnhZ9wy7tFHPYUhxAnFepo62jAAiJzpNN0cQIJb6MzPAAp+owP/MSo
bRrdAkF5FnmRk0WqsNH3t0kgK7xhVzSX0Sw+GvoL6i6+uaU3oJOL9M/K/69tsG87lzuwGeuBVlWd
oDayu9I+HPDtO14eNiqDgJ4qGv519pSOD/hl7nhzZz0TtB1XfD0FIxYyp9nx5HWqA9gnN3qau+cE
A044AMMDjfB7gR/mXVLwy7tWi8iUcJo6O/shLKn1HnPDPaWtUBQX0mwOJknjiM+msJbT8FQK4gni
HBus6UBB+MBPP31Eiq/hkIDbX4dqpkkdh7AuOgAWQkfyBkmZoy5sCzAR2HMJ8uG3Nt97sO1xV9mU
ioGZ44eIar8f4b2EXeB97yGqX5fuMHUxRwaHAxx03KW8ZeVTuQZxSShXO82YkHa4Fa6CLA9F7v9P
Ljz/YwPJd8N8TSR0mogol2UqTVzdTruuaQBUdaEo169v4+DsAStbNwBfDgeQXTp/5e5UhOZtf4F8
5F38YT0wYyVPsTcT2IT5Yu65XS5BQc1NCjQ77U1gWmatfPE8nABiXpWRfTxg5L07PsXnL1KpL75s
fxlqZnBFV7FWThtgKw0OPtGVcldsVv37z94g/6EHbLV3id5i+qtbvueUhjCFwDfoYUEw7Y5Vs4p7
B8F4YhXlgK9b+fM0Ca8aSV94MKIx0vFC+T3bRJzO1PkiQ5UcwV2tsdUtBOt/eIxY6xd6AYu6ED1w
udfam3LtACd8zbNJ2W3aDbZhbem+1SdLzkQ1E/MD+J1Mm1cBqcI4zn05u5sgLo8L70f3MjBLqRM9
Yv5BjzIfj8mhmxiwxYIvZ2n892TF/1BfWxm55xCrBQkEQsMdpAZviztHfxyBqcSTKKz7zjCEbRLy
E07Qx689KRxsvUzza4kQ09tSmkvRt2uAFoLLgLpBlUEwdVdtSv4nKbZWIKinEpkdDs7PfrGAnlGz
E0DOjMk7wD6HhQCwBgv/Getph34YBMDYV22RKJP+97bZLE+Rde29Ib6Fo9Niy49YJdBqsGd3ju/V
JRGcJwzCLgejwtM1ayX4bCZTBxkuo+4z3TgG5lgKJ4kz4WaYe6qVwL1O6yEtninsRsqIIUHPs9LO
vtzwGiQBwDaH4xbZY4iCtEnQEtp+5xL2rilyeTCz1eYRq4Ei6X31KdOdQiARSfFjNRQnJOhtswiC
bREizkvOTa1uQsHr7ZxTNlC9yCq1mSTJYxt9rM2N71I9UgNx6K/m/w4uZQypugBEXueQfvxhsaCU
CHEQdJ35LAN8Sh6l9YFFCLmMePi8ePJQ546o9OGsI6NdZchgkZ23M/cW0sTnCLm0o3zL+IpEz6Qx
bphQCqufXgRjmjw8iUv5jknvtGFxFR3lWhPlUQaSYjLDD65AazCYAivPAoBdW4RWAomS/3URGW+s
gAVr0Vc0b4xLuRNVdCug4g0puTgSERRHw2u0x1uYcnDrYBOcKjUXzU88iOanRi2uPDlzao9qf8qq
J6MBXuojVs9ZCv/B7n9NZTHo8Buv7gMMvgJhsSqT8l8xXuJEmG7NxepKK9e1nDaGbrsJeQKmAnBw
mVc8Q+a2JZ68AKu8ol9hKP8cvBxI7nf+pPfKj0hWjNaKKeE4zlwbXr0i59Y/tRd93YEu8gOvSvcU
SMPjJFPSDNoH0vJleQxMnMRAt+jNxzXZPL26f2YVW+S4lGZZbfFg0pBKAscI0Uh2NFWYHIaPCdnn
5y4LRN5lLuSXO/xmsVRhUyYJkzr4SJk/+6S0kgUYzHCEANth9Qu2EY7Sm6CJZ79XEbbFsEdnBq0P
gvAmR6kGmSw898SMAQh8P13lXJBo4Y/ikU00+oghY4TKbv5V8vhTHfs9OUNyLGrgQ20404HvAOz6
05vEvU5QX6SYtyHyUt1bpEF2GqwK7BC89QrfS6vewSSeXad1IrnzLHp15/vaphCaBdOjv5zMOVZb
z8dSrVTHah5yz8SnnSgFFh/7GgbyCD1mhY5oY04I4bxY+IsDR7L8+YsjEs+T6KzIYKd8xGdMCZ0V
etlOUxaNJ8umDFUdoi0Eg/BnBrAX7Gr9GQjQUGP62Fe0NWqMoHp6e2ng6qupDUAnR++Edqo4pmEk
IVEiztuRCoUSSWfsrfThpkuVZjm0xwd+SJSLuczmvjHD6gFaaSnv2bi/+hhzoInIIzv4+470pvZy
XVQ6ad5x2Qs+Tn7CQBu6b/nwOrADVDMmwu5UqTuk/J9aushW822vtTTS6CbHrRAd5C7jCizVSiFO
SBWA0I8TE6TPomZCiUPIRXziZ2Uw7EpfD2kvuGduXrImqFLmtvLBxRQczepRsX2wEl7wX2lTuj4o
d2BkfMKavrL0DjGCCvhTSZeUh6qL8px1hw0ChrrcMrPLR4Tj0LNndMBk2OysX3A77JOGcHslLpLC
URgqela5tjEeJd3ar21dXh+7xKxx7w5ILYbiEU//DFBctnD6esJwt2mi3ukLoA+bYBNiGtyzvNIu
9KXUSNmYWow867R0nn76BqzmFe5NUw0THjXlo1w4Y92qgEvxVAdXKBlndR1zkB+4Q9wagGkUCIrB
zOGANR7JNTtbGiKoeWUtgecwEtzx+3UgVNw385VT2weT1onm7pSPDCDqSx9KVh0FT7KlgsSdpw/F
LzwIpHM3UNFxqBLhW1SLiyHhML5K3y1Q3UwpaT9KUBZf1ItN6MhXYKHZHExZv6JrcDc44oLlEB5V
92D9viHvRdcnwI9d35Wff5jRynt0eeW7c7bU67vDAQj6awbUkKhqvLjURzE4hAZ+U3DwAEkfl61y
isASXWce6J3ZAsL0vWFVcN4gQCJh+dZdDvI5r5Gpurgk44CTCSGhtrqvhkjR6UeMHHwxS9HPEde+
CQWjhFDEM/gr/BuPYJdE3T2GClIwKttCUG/uHuzaqJv/BD8h1APelW1Ac0bFB6u4D5i7WvvCSnfh
ZD4KS2Y04V+oLFr/Bqs/OU1qK0/ppKKi8Lk5YBbxAlzmWq3uO3zKGADvP6+Rw82uXMXipd8eAJ21
0sdHNixDisGOuFTIw3G9RAxfgOGNQuNMYHcIsTE3+f1/NRFBVoMJJXSWgM9A9nRCJn53CqAh2m+q
b1ONZ8iP3ly7roc2ceoO4sv3evE/XZ+sRX63v1wFfJfzb+FualU5u6qPJ2qJDBtaq/gwVPqOb3bI
2c31VRZHvA44/teRF8LLOSkqnCZRj/pDcDas3fISyy9BpMWUtzA1VIlyHN5EIidcMwHKInItSzRh
7egAwTj2j2x1bLWhFXdGXF1rXReOBRQ++JS3zgEZsH4vm92Ts0gltM9qddUGUV9alelx1Iv90Yfh
d5L7jUf0k0vtMQqRn/infrrWshc9eom0py31UOoDnwvqf1UTzq9yFGc5GDe3HKw/re/4Bsp/883A
TCYlrbQgPCCHXH9vT7es3XP2ArhiPS5JrWyR8DVqcICWXSLjhNy/ejnB0i1NbdTBUg8v3kavGYQp
t4vktKC7X/0zFMJot3NxOX1wOnzJD2LSNr8NIMOy/uwVsZ08Xes2/5j8l0w6+PrlMckYtmL9SpeK
fAmX+1knERN5sRlFJGIUPhnZ+fPcca+nw0/WtT+aNNRKuqKlFMofFLcOiB00ssIRzC8291118AyJ
kmekukcbEqRvIDxnYcSkZ531yfiq2i0qjpsdD3QPutEfT+y+zzDfKUPjQVYwBDrcKylzP8JGqp8Y
zr4pc88HZ7tYVQJS/ScvPbwCG9Nr1mZPZRm64o6Sq4Sszgd9S1+QUsOZ9pESkbBfbI3+oUJxnXGq
nKeBbFjlpdt0KLDMP1eouGgkdnuEKszDHaciGBsg5i85iMW0UdekycUSRffbRju+qBm4Qx9LQSpV
LLRqwhyA9HrNo1xAgfjenYTgOZfociJB48apwfq//ljrnm2SzUn575GuLHr8KWTOhhgoHIfBwqoj
FJaOybZ6GfRfSKMJxqze1fOismDoWum3mlHrK6EAwEWH0tz4Nm9SF6Xof2HADtV4YDPlUmobLvto
N5WP4EJlk76zpI1FwK1rBABSVwRTQIcVt83lRwZ2bi0UMa8LHSHzlE5MTuZN2My6e6a0OTa7/7Q8
eoSJtAMy7G1tlJSKwGc01DlbskVOAEtuJGiJD+afUe0+J/zBqTyH5eANMTBidq0+aYyyRVWfBLqe
gv+fNIFoBatXDRM9cI34rZBIGdxDV1gtcgNRFMY2NJNr/wqZDFM7pWpylAVY32SiuGSu5w91Lddb
xVQ8qMumoZqNg+YoTEGHtHb9nJR67i42ZTXjGnMBlvJ20FLDo52Ty4Qdjlo05vC0OykDw8i9ex6A
0S4d0BXucdKTKciu824lEZgWE87avg9UXCzSyMBfkipveeWKqe2/cKCKkfKKMg0z
`pragma protect end_protected
