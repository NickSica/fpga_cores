`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
V82h/mp8FbHcv3//3zVZ5VW10Mue/LSt5dvjsUkiSGtG5WaH8H9Fv7j37k+xy+3/pQvfXcpqBF/k
iaz4/vETUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n4WSOWV3uUjyMD/l4IGcKD1bHONRRplCKgax9lu4YRYlORLHEpckVBvOD9geZHtnlLIjTLNUcuHS
rc4oO2K5x66eEf5+m+hNzaPYWCrVKWQI7/tyX0imMAsD4JQXzU2CP3ATsQoldRyYOQZmggmbIMiB
stLQ3uoRuVc4t0kXI7U=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zgo3FUzRcS1G0FRTCr4C/JBs44dp3dv5CUvkYU2vM2fDyGtu9ekJcjDXnFGi3Qx2X0BV1gEyWxsJ
xqQkFlu/f/1mutspkUjOMtKZNCgPGDHkGfwBEPN/xT22fOBwQJUR+Oj5KSeDWe2U4t5UJ4XXcGMb
ZV9syPFreDWYOTWkkl85cAKcf/WXC6oz+tOUowqV4nSLA1PaSrK4ohf8oaOGNVX+4Ji/w6ViTIJJ
OqmPJQ151npm7Kbt4RW80tp1OmABkNI+o6h4rwtTS1IHzM6bJ1Krrp0V+2aEmmqoZkuKINjX5Pw3
P4Vi6iUmJI0uMpdsCPr3MEC8HH4v95WCnjh0Qg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A45QQ9IEoKpoNXpmniz3AuFZmGAAZIhtA2hP4/pi+Iwurx8nPI4ZkKpYXPnn4DfH42bSsec35aiS
Ve+A8f1Q00bmFgtclspinRe4YgFesk40ftn1mzy6g6sLCNXhUm/IIjCSNk+ie6jVQS7STfOdio+z
cvSm8QQePoJjzlJz/jkNhsD110PhDAevJWb+C5fforY6kT0k7ZmJmE7btahod6wU3o7t2HM6+XGU
DDNZ5E+RLS+IiJYVCOwsdqQFDuRaWwS0k8Mk4UuDiVWtU0+QLFZ/8UGJhy2ZDSYlL/8TrrsWcD/1
Vku2N+fkWCj38RSMWEEe5TmUHSSzP7uBI6QwVQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b+wEsHDGMmVXUM545W/2toIjDItLsHFsIOyFDid8Fv6KhzBePVZlc9t2c1LfdAa6UEpdqcx5kgIr
+oVEglJG3R/fb6dRp2mvlu6+x0AYh7FK0My5t84q7uKZ6EPBxHnDds9FLGQdMDUFv8E10WtGrG31
lkto5q+L5WLAzYgiD3//MgdbP+aqLc/75XWIRhw/PfRn4OqyBU7xSBeoK9TDxBwOscUv0cQ+dauJ
dUQ0W2ZCXwF6cP5c47k76Ikfu69J0/IO+FTLKMkjAB7Wzsyqbpl6RMVdJ/iYscNROh1xxo2k+52w
4l9VnVKN7wTWZdW75B3V/MsNTrKb2I6dBdveDg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyn/owx08GdB/M0CwlYM5XwpK1DLRGgNdNGvCa53fvz5ftb1LM2R7yhWTTXlm8iqXlg1S70wvPmw
WVO2ZNZ0csmDdQcX4HNMiokrI2gpR08Dk8n3nzdOhqyFyh79/eVJzQItyKMQmJZNCvFfww0mtX5K
FbNe2x6ria5jEBEBp3U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J8WwILioFJtk4e6vNsFHYZhWTjvAMbsqHcnvhYKYzsY6fpaoYuWnjTNNNxS6JYZj7bKOFgPjdnBA
rKaGPLghV6UU9fx6UcBVLjNOj95AU3CZPEjWGC/GqjGRPxOkhGtDka91PZuOBRTBqJT8F+5qIgQR
vO7WJHaKezpaUm2zbeC7+ShM5p4Wm9L4dzJ1OuUGZNm39p9FbORAZNzAWa35wpfJ6PPOgATFMi7Z
sN0Hg00oxMFCKSg1bxvN3p4iC3rVT+wV6yuzOecq97B7Fu+tfvP+shqnUhodTpF0WYfGWHeK9ocM
Mg7nt62XJybi4Tm5rgYGMIIM0i67934etK5Aig==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AF8EDKLpUnsf5U27caIfzjHsL1dKCT4FvrlOxjBwD3ZJ9vsXwbWO+EJTOJOFymKnoSSFnuslr7C8
ZCAbkJJLJrLXJwfvC9hiPRksxuYzuxWrtwsjJd+5KWtue3gL5kHClD8Tbo/V+Dnr3gvKzMRNdFRz
i+4p8dC6/32xR0/NITJMYT1uOYu0oBFDHGLR02Wn4PqghcTR3gQMVeL0RsDhJibeNnf4Q0NsKqCF
7OscDpis6r9ZAFao+mdpLGI93rreTlZvJBUPh2RcpqOjL/8IUv0iM922KOCZ6j1LtvD0igXehvHa
5hOx0DDcMjOoejqJiwIqLij0FB13lDBsu+fjWw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 142256)
`pragma protect data_block
BMP9G5RAk03qFRu5UmzfhPRa2E8EtqJjN3D5ol0ioUhd1Y/pnI+Z9bsxRy89+HCs+ZLbtnwytuQj
294k7ud4UXrXma329SxCtsgGHomzjQoQlIpv1W7xtWBQ5Uo0WbV46cFfgvZLtnEWdDebGekeHw+7
H2wGCqx3W8wzs07Hq/X+h+ynA6ATyU+BBSX02UnnB4i+1grO3DtziDbJtZu0gMMhS4hI06gDMDai
S09+ZvA3xCIc+BSB5Skb9MluyQrMaBFZJbGTcVspRpy0R2RUoj4qb7ikGhnA2oXT5kEVvEUsY98a
vlu+ap+u75IzRLtK2lI4vJP8XW/nxF7GUOfUrtWr0D02urAdQ0AKBqz35T7+g+vMg0mkg7ClmzeE
v288fAuhUFBNrjd1x/BZ1xYyzbKcM1LRmwBeR5ZZEMY7BzTDye6BwgjZvwEYy8ZoSn6LwKBDJqVI
70x0iRiSoagOxf1idakDXglsT4zX9jFR9ggjkTQld8xr1SMyk9EPWoiNcnf0/udk9buwnNxETSqE
cUDMBseTRqB6uqqlp9TtZgqBbppagnr9v5ShK2oCf89ThZdTKQbjMUTw3zyCP4DVZvs4xQBh4ygy
k5FgaJYKPME3yMsA/82srjUGvI7Cxh3D36HuGzCMGwg1lwTSjoGudkjkx9FjB+Zn8jb9E5QjyNzO
QdflUgIvtIh/LrxsnH1g1xzngCrEBfEs76JafuSYRe935Z0LM0XAm895ing0fRWuxDKFllED1g5X
GoEuAFjhV9EDHElfSWQ8QaVz+OjJ9icP1kGMVLfV/8gcYDT38S+HiIH8+g9gAw3ort5tccrKKfbO
QxKol7RDOyErerl0wXdfJ0vao+7hzE8D2IpkKmc7Qr7lOAwXBgoBGJdwMsfrVCm1f83gXwPNpfgL
0bql4i4gh2AmkMeSPU7+IIL1SLatuJE/hiajDtwxAW2k6oT+YZR4bpu9K4M0athPa/SwLzzmNa0k
68B0UyueTnpFUaYD2h1zkXURrmTG6I3+yzTa5N+yApGOsBrv4Ikemtu5vZWqywFaJTpDRdjUlyHR
Al5DcCOVkvh+GvYy7NCnjWftE2JiHWnVVf5HuAOLFdSTNAr9+veKt/0fd20Hzm2tSfXDoi8Om6My
OW5fn0fHpSfiGdBXa4efAC4gaXYZHlkYPzXnRSgEmUtZ9sqdr8YLfkmJYtuhsSl8wKRNoqrAwoEZ
IulqGFI1An13jUvK/1eogaJuNnC7X8knjqOiEdLEDHa82cEKF3tn4NWcr4oFm1QGfcHqzlmdYX4l
AloAGH3oYDEDYCbhK0lYHNRG5duY3dCSJweOW2AX9klO3G3k4P7TQbrDBlc87pkJh/SLZjNQSgXH
yGdvXkE69dU7MlXRjkHc9fxkUu/6ANOWMtyr2RLDeFlma3M+/pr2Dx9pjBhg48s6E8wKb49nl/Pl
4bITES4kdb48QecnMl0s9r0fEX3zfIRpAvmspiV00XZiPeNSjV9DmFX2LdtjcIIP3XUDfqestEp8
okaxLj4Kdilbt0DKjzryPLKhYuG9QTq4JNotKTMsE45loB0r38dF1earVuqZ4WLQoVPqUL5KBviI
YOrm7alYvmsrOEVBr+hIrg1a0CS9KsKrlfuL0Uc07JaGcHqwJESScBzolQrdjde1AG8kwOxqtz0Q
0994XHAVr0bweT75PkLYUZIjmP43/O8P+AYNuZN6XWmKcoDW65OrNKmhV0EfCjy+ihBRAK0afOXr
g/PmqrQTRisaO9NLgsPRatwBYBrzkMMlzMcqeQb2QdiIDQdiDvNdL7g0MLh2IZRQOZoAFyJ3VGan
T7bYqQ6nnzeJYkDqOC/HT1z6wCT+ADoX1QUCzYU1lX5twoyQ6u9Qqo9x0fuJUttY9u9rvHCKs4z+
tLtLwkqsEJoKIb4pcANxzRSO8j5kR1cEgS+on93OI8omjvvpJjtpgTQjiC6uISZ79b3GsmyvTO4D
H/WuycE19Sypbx5Kn6qQ7bel0BmGj9aQN+TY+R7Y2PWYbLglwhV/pZ3gklrxLwhKlXPSjtV0yTmo
TccZsVxwadfzQtbzV5gLAUpZcKR3qqAnJV4AVrm1PwzF+vEHDrAnhgVsSq0qHyZfhDgFpKW/tkYM
Y1923VWb/DKzx3gW2djYAK2UzXdbyMKekyoUdDufhRh1BU0wIOR4zS4XCO1VXmkLKBVgLavvZboI
lheTt/Vu0PF0MjFmj4EpS9HTT6PUpsUjmtsVuBdSlN91LAZSLqwUpmP6J47QYNb+qRHSa39TA6MI
2he9cQwd2lKO5Y1UG8mClh5QsATogGX5zfq3XzKltsHw1rkqjVickdGBT5UD/JqXAi0LZ15piUlK
ueU+xeKHeoCjNdcUAPH6dfYQV12wzWTrKjUlWDDBeitQGJ8X9tByXmVgS7YuMlztLSdw18PX0Trh
Dk+VluqkQZ/Mpoa2vuql394R31OJIQxyeeNPW6457Yb3D57iu7ZE84o4aWtAwjW7HJjdCWBXkosv
3S05u9w6pVD0+AbEaI/aSNl748YCtF7sgS+TEQCfj52Uud7VrrIC6Sb+LLwhETAC4eoTRVo3HCMs
3mRAVnvLymkfprGgQqqyX/ksiPQ+d1dBwRfiEyHKe8ELcSrvoQiBpN3TmSAIzp/Xxrjo4Sto0tj5
sOF+DzgvzrLzyx6qXrxg606a6x0nWX/1G+BH4glvfBUAuHmkV+bndQOeCPY8lC57fb21H1MqulQ3
eJ2nuU8PLh+WPG5s+ExzanvFDsM7/T3Q7tPn6AJjaZJbjqp+TUtzdafg5lvD35Wmm8HZSOfMS/9G
A5LQZmGJSe4Yc/P8oW8dOog00AfM+9t1zK6fBaZQzN1D0CEImk2P/DZJXBFthzm3X4/iQsKc8tcT
AwcsuxLaS0tys2vqiXs+3oYIC7UL5J0yXPH/j0OhutOBt9EhBlYmIk8lVhi23mxsIOGlTvtoXZTR
j5Z8u/JE2T88D/OiS/1/OD2eWVtGpHKHXttFx9OuIfUIFG3pAU4aGRLzSzASq2/CeszDGog/alWm
nsP/sRajzbIrM+DYkBH38KK8OrrbDWehUfumJuWfuyMm9c/ESsNIxIBruNF8S7VStEZzKPURXA1u
iiSUFwCqPTIvzq0y0naf5qW93ydOf40EsiFJbRMhMxKOy2/Mwc8SK0Gz5FDpImb3Q+vok9tu1DxO
asAxsCQOYarDJZy9AvRpQ4iVUTtfH504z0qhWcEJY8DK6Kn5kFaXOpGvAOgHp8Q+Up/CkYLyrdlp
LKZpMHTjnJ1VxamAYymqtbo9ERiZWATyaqQYq97RTudk93iOyFYH3HLYJc86NMq8m5ObZrmFVjY9
kNFg6LrKtXhYYk+3Q0dotQgclxCiWeADb0A2M5F0R/JG+QbD5TZK2Ks+vrDSKhyejzMvHMiIcrtI
FiABIhRoy9S+rVfswNG0ZTPurBeg6ZBdiyDWLD4JL5eDf2u/QLSYeY36ayxyaqFZjlRqCAWcvRzv
/H1PZK+UUq+6B0tD043R1E+ZDDIFVimlf3N/b6crpGmwB5cC+6PyaSu0NUYNI0In/cndh2ezWpX/
Kzy/NEUYOP/wyCBse/fVhI+/51AmhiQ93PJ8ffROS+P1sKYJVfCG6wNWtubBf9ZW8OK4dp7ecB+/
riLO9zwoI1ZNxlc0i42XWtYB9Effo+BxZ/DqPweMknrb9L8lA6kAs71i3GUNIvagb0GupqiGQME0
X/74E2jXxTv1ZXBGyGUY62xWZY6kUQHc0AkUPi7Qo9Qa2Uhh/XaOs78V7hZsAFcuh4SYHy8MgRSh
Ev5wX/XLIk1LkxuMTTnadi3mP9ic54yCzqL1gQEV2I5CkAOET0nz8JyQVqAgU0tBEIuc9DkjQ/jp
5hd5iON81eSynWQqhF1P0G/0ZuDY9qdMZOcjXcNiuc7bfLypgt/5U/INYYN9p2uMr/aMZqLJKDQw
AtMr7PcHb3+2G5zTsCe2/znT3f7aG9i+iLEDNgZMtNTzvJt9Z2gs97afWyUlEp30GwXFuks/1Ylj
OCxs1wHFpqDlAt1cUlqIu24Z+PNfy6F9uP36Zz0B+YESnNEcKz0iF03Q5OxemlPxQBFm0RiFPelq
TyXYXHpAFTThJGcxTs19iAJz4c0mtu5SqbxRjWjvywuW3YpOh7lwQmx/jIXQ/MAVk+Oe7Iaqwub5
jWB4XcsUoI5BO1niM8DYwfpD6fEnwKYedFNnDBwH5mCnQ7nRrfcljOdDY0lr0rPg845MPaskkpco
ZYJ1UeNLAaqIYeiNst6eTS6TDVufRUk7nqA94xTe/kHcHQ2vLWS+L4MbnJoXvr9wdQ8cIpWjIomH
mmNTCPwvVYUq7WAgoKART7aREt64NollHwmpriX516eilcPZ/6eDDI0SvC48FU0uHTuPUc5nD7Xc
OctM9kHpF6bJS0yrW8GHTXWmy7ewRvFscLlMSaSVDhBvs/W7F8YY+sLPr/gSUmHr6OOpdWMejG/v
s7WQn9DY1AvOVDKT0WutX3yZdW7aoP6r2SfcrzyEkp40JWc/Y88kXnGzNQFW+UXLcmKHfVKgDOIB
Thjv3cgixFXl4/xs8L6fQZq4caPtX2eTQ2lG74yDWlZFTpcdyFcCH5Vu01FBikBme84sBr4Yz5ke
9XjejdAwqTn3HQQNs/YXPwT+hfr3M2HOKNx5JslDl9+INh8Rn5AwgEmkztW8NSnrUuFVNojtZ/6s
IdPh09cO7vCy8nvx8PRcXUjGfz+IE+AEWpoYZIboNJbtm5OVALU327J5zfPS5s14cIa789jmPkH5
B9KKypgekF618dSdmrlCg3LRNE0/FJ0DfDMJmAyLwnjBB/t5hPRjrY/RA1SBJCSNrYrIunUeou8/
SFN5B3lN0CpHzhuFzzm9eOrQ3804uo95/J+0ATbGsc6pTdpzbht5fh0y+LLMic8elFcZoy9cw0lg
QRUqkrpst6NdqRoJGDxFCX3W0o646ZgzRw7bsRatkc0xVQQ/fT7gW2+zpMJUcAQ0gqBwqBxM4tbi
ff6xexRwBECiJ5SqGkieCzvqoWIbOkFNHaVhMLeiG2EAfF4uZ9lqJD/JLM0bnWmw1XXLKUZCnbLZ
081QBlatBNvNlLev5yaBjP9H5ydK/XPC2HxGCsrb4byjzoxkqQlFEmybaegzwx4hFme6ve0l+aJD
47sczpjGUOexi3op/zjBzEvy5JB1RNEjcrC4R0VFTTErkvrGpRRRpd4wAflZlgQIA1tFmknsgvhW
5zt0zBg9ukri8b3zULkEx5pjd1Eks0yFcp+Of3L4CLbEEjumvV0cAdOcDPe4sxtC6caRRp7bCbg3
cAUMKslFpmNW1D79yoVtPEl/++Yr+KP8qZbYboW68HuqI72tlt2AkbuOHyUS4xZgBCe4Yq55VwP4
LnsNqU0pcFP9FLHkiPFnl47AF0BB+GBhovGFE1a6M5f37NmC4+NKPahIBthsLNb2GSzUAxWc8Fyu
zJ79Y8ekar8RBOF6IHSBrrHrUio1QoubNWEenFoglWFScTZpgyb4V+1DAVd6FHV7lNIW+eiSFdn3
4lmCxObQ2w+sf8hQQZkhOfofXI0w6u/y2J8Ekh4Z0bhjDozvFZte+5XybB3adhusLo0weTs7Vqx5
qPzdtcJqRlERBo6KqPFtUrvuXYJHliQLr40IbqOLMLHl5EYSF2bk/g5EMcyupHOwkTAS/M9lmtPg
fKP+tMJCKKabU7rULB2srutHVWVB1MoEW6qUeZA9eVaGLnUzUle1wdVk4zdQAK3b5yLqcZK5rZgv
JZk2gUluCcGgo7/xD/geUioMzTV2ZZi9YJVgvaU3sVmqErMQyseWxbmcuIZYoFIjpFjDh3349+fD
eT2ELW/IilwT3SSjjA8df2GF324sXWx587I8Bqk5fs/4yZoGsZIj6qhiGLbc8S7ptRy/tHmtsqrB
mmSFxlQOI6D7thESw3kkJjWVFcAd2u9pH2T8xFLC6MZ0tUWKY0Y8TJ178hT+VN22DeLqMdAAqo5P
up579/8MJ3qUX8RO7B/iVCbSTF8zG1Fhrom5kPRJ+hK9uT95vG2GoHLq7kuU2tXVtf0ktYaTYrwb
EcdlgWImwRIbiy8QJOQYTh2VrcYEDlHe5G+OC64uyqdyiMUjQCBia7JqcRyyjFtZRY/VTdDhZwB4
J0DtfQNJuUMp89eHoMdrIOsTgRPDXyGOpKnsZuA/D2ajIuRuVeiCQcawi+j0XSsoWFmTwcs0po5T
TneRnaPmwWu+gD+hNTqgvz/zaH4vvzcT0iGSjV5tLjPbuPFgAI6jRwLWcSnHxVqUpFX+xsWo+yTz
Dz5tD3qOX8LLns1tLuxLDsOjAZu/fLUV6g54UosfOs+x+kBX35kZgh6VB53E1j4wEnKaOkduzTAB
sfpyKa5yyiza5/hCREGOG03VMXMwLH5lkvxvGXa3ljofXOj9PlFz1MLm/vm+N67OYhi057mlcpfV
ABwX1OxQdxV0dgZ4Drpr2ORpZV6s7Rf71WOeUX5mh0MusF8appFb7eSvYYHUJDlpRLgKTrnhVP99
z+RDLGNdEvfCSTTlKFbRW/MX66WLEeNAW3zp55c+mFVUOtoQ4q0VRRaKC2dOWk4lCEBFhq0qiHjC
d2mz9J/lGfTCjRPyBdE8/SjA1OEdvbfho5Ev3iEayabierta8tv8OLzZOov+5VLjmJh3tH75b+De
rfAlSPn10SQAiFyrKfM9jhfd2ShjxGer6te72gu0AnyNWtB9uRWQxDp6P8rcjeD2xzMdW+4BouJL
balqVkP5+4Y+Xt/7oAGTCsm9EmCGvn6QRvQrgEpnxNKMzGlc1MPWXkipZHiktmzwC0XLu+U6PmMv
4bzV9VCH/90nThjTch0R1UshSmcHcsY8uhN5+WAQv9Y0LfYP+hPQG+jk1//Maue3RMck4kVCzUPp
EBptdWKQ9mtGC74/paIHblggPh7G6xWXIBUsvEnXG583Z22Ya/bqXWHQoTK5coECtKGWcllyzY3p
NcDgV0B4QkhwlnxUxeyJ52MH+h3jbiTOCdbsMeB2sSIh/bFhEwLAXzzJjKjv+icBU6dawVmE7siH
0/Vh1u71pfXvqO6a8b6Mi1is1MY7kjHKoj27t+N64ZMNzzMjC6T/r+DSHJ48XHlIJHARxurvriZP
KbrMAHRf/t0oXGp+SwM61NfUGQxM6xxNK5RjTDdOp86/mLoAo9ccRukG3FH5SEJJhzj9RGbRopkx
sbAz0SX52LECMkQjVfVyonvT+tKr18bY4eS4ZLc777EFrloD3zzF8SZz+DYU125LB8rQj3YULAY0
gsgIKAbXMYhPSPRlx+Ld6WjVXEkFdWPtZGr3lT8c5ZchrMPAnE4ewRa4QBir3rO39EHiY/FJbdkv
IyAupUGq1mIl3BQ9eOTokeWEtppXzFLm2UYSnnPzEcWUUy4iAjPFQpELXUNT1KftzjCx8iQfw3aj
oD0jqmXIlLYS6z9RktNYVMFIi65PWUy115/YJNJcQctpEZkP2GISqcs6ttsvPI+g9uGuueNzp2ca
QE8v7ULKvaaVDVX/BsIyhKD9fB4eM/Y5wTxSQDMNFnKyXhWCyWCdx02eJ9h5wucGQhYdTkqnj6Sf
XDkwdneh7c5XHjzJ7HJlcEj/ZppWzRO76nGKDPpHVvkuARbwcGR6vkhaaBfj/yM+6IXxIC+nB4RQ
0BFxoYNKP/o6+ezFvJeHr2ch7bTg/JjEdCx9XdbZo/NwkSM56PCPJWL5UnFE4rKxvioO1Zl/XyKt
V6ECOnhUSMRRXACgYSpaEIonSWmVUu7Jt/ApqlfDatBHD3icOHbZyaWyIUSgmHn/P+lafKKeqPWH
rm9hf/tt0llVZcOK88yrT5Tq9Fj1fv48XykJsI77KzA3X4IXhDq1dksF351wkvMt4aiP1Idh0uGg
vnFSLTXZc/RNxcQ9MH303Uj/WUATNpi4B/VNi2MdRZ3F7Xi/FptqHZOLeb/S3B+bcYX1zFee011O
zGG7vwIuVJXpFmH0YwlRCkgWHKzlPIGYy4gAuRcBf2OWOd9dm262Ks/4pfgUDe7clKksUkIB26Hb
6UWGyJaVkNg49HWh9yrLPXk1okBplHV4tK7Rl/gLVNz+VJjv0EIVeOL/cnlRKoOBEJ+aw41R3yDQ
LmsmWtp2uKjOnC0nCGRIzJXuxhfzqYyG7LqRlmtfC+NjfUshoEg4NwnUgkHj6Az/nUDUbx2tf7/X
ECiXgobJypvKgEssiQ50k1O0RIAClp+izXqdmBjJ5D68cnAxn3jVxPe/2jmEkWmvnytdHVRM0nXQ
NVPiywtmUCvKx2kbRmRJL6wR4gHlceaWnMgklNdPIHfOdaJpbyp9CyLZHdHkRqdsL6RF+iSv7HER
J2lAa37vWQlhfodsjrLQhMKsHkBswb7fao+Lji36R9Jh+fmzDbFZHbmVC3iIBGgxuxTZNnycJStF
1dyoDyn39a/hFJs+fJczrsA64OECaDieqsVUP8y0tWRT5Ui9OGsF7wdwrRNLXDJadbR5LXD8mxEj
f/PDXS1ScSUtj30QvYbUSg1EBskYOT2tBpPr42dfF7IFiG0lbJkOeK3WehjdSV8Bj1JvE8evQ+l/
VezNf2uea0kvBy6JaMPZpS5V3RmXIJZdk2SD+LKijY5n6T8KQhi8+Ms1vjqcMUGnSjxmhoje3beU
Wgq4kc2h8LybVPdp+fU3unFyiZkdQPUFaEx/JnzSA6O+i/h+ANFMaWUO/gboX3w8NCaPwZ5mPQ0D
UAuWLgjc2z7UOPUIDQUIyBPL3KpTs0vUwe2lEhFqA6X3W07mV2B94TFJ3KcAYuo555l3tcpflOiQ
lqB1v6ExSugbNNHxqWuZwP8+posfxetSxcb/YDZYTyUlfRwv9Tzwy/FqxL0udtCskD7JEaYRqF1k
qmuZBKy9//iwif/Uv+osG6micsDuXhnz5YHFFJ1wfE9x3DpXzlWrLDUDS+5q3ZgRMVqj226WaV1s
boMsjn9uh4NXFa1UytjN1eagKKrDs/nT+6l11wly0WwJyXj+03oyk9/SfpDAHsDgc1V1XH2UPWFg
Mg42ZDRfPTMSUaEzzWjTIP+AMbMnL4x0zxExvCOFS6N3SnvxWrKqniSwEPZUDzvxZx5K/L+FCTcG
kTf7nPffQyvILuofDrJzfpOtebZshVk3op9vGIN9u/AJf9U35MSDXtvozGhzl+jYxwd7YGyU/GfD
MMbW7qqsYtfU8Mc+Qm25uy5WUEhij8i0ky7E0sx2lQur7cGGkFANJydn1pxRYBHU8NlS/MLeBKzV
DAs9G2hK/ZAsTeAW9JH1Ar4Em5pgzbTSBZLHydaxjM6xOjESeS0uxt4wP/SY7GdCNZPqsILKjaC9
FzHkYkY+TEHSAnPYhyVnHFOXvsunTDTVp6VIRAvZ2iuAGzr9532wuNQqUYAOG7XL1IK533B4erd8
c2FLpG8+2fSMDY/ryvRTJGU27yn1uFlVJmSKjoUOAh609cCA84y7qn12Nl7CnmGGO80JqEsPdeZ0
yJVpDKEN61HoBf9APadj5D2llAKrprFutJ/oGcReOs39aVtKQxZmq0ORwSqIOS6ubHH/sFbPF8oD
lGoNd6vC+0Y335I50G3RbdahlsqwgeQ/8YIsMUJXMi6srlI5b7UmWewp+QNdRm/SafB5qkBv4lDd
49PHThxZSIz6O75wDJ3qXUDopNwgMdf7l1kqe4G5csNBWEyIMSkpgSu6OGGNO5VEPQcBsxbyfRDY
Bqoo6dP/k77zjTCb+wp9bhm2Ay1IuzfT6ylsvdD0cZNf8KI7c9WISxk+Szsy0G0LELi3IRE3Cdwc
xMsuXjzsfS9+hTUovcOfdbsGhCYa1RSlmiwIn0LsFCXTffEmaPWVI04yfJ0fvSLoQ31IdiF/fOKB
xBc8Rb47mG494abyFgEqVueP6hGUIYpFybHcUSio+ZznPisLhw4SCAo7oCXavQRvon5pJEfZoeDr
YVOmdFQbBX3xqenoRd6vL5rtfZgIVck9+Skn4a0rYMbEvNlcUY2bvIKAQ0G+tAt9lX2N/3l7ekD+
eHuXqLqcJM2W/xVU0JJTF5I4dcUmIN3Q2gi5WTeetZCGT4MFOettwQCI8XOA8agK8fT9cX1Z7bFB
9um9PkDfFjYkxcxFywrUUI4EEUbkB7h9GQ+R0UmdDjSiXG8DU1AubQuZQe9fir+ZuRmtIVRwRktB
eixDr4li2gl8+g6eK/0kBPx1zA4GXNJ8qFNabxzoW2U88JA79/9VZUNUjDbDVoj9mAdVccDmjptb
r6vXqt5s0QWFKgiuw2aq0Rfl6sbM2AK0tU+KmZCeASSbhjb2XGWlKmtj5wnAMbhA8rQ9XIO8rD32
1U5frXycuII7slKNKzcQk9aa1yyP0pA4qif+xuv+y0KLeOVkGYKJkdyTex1jp/5ZWCbjbb8qpR7V
/FCXHURRXd8sobzN4WoIfdWu0nr2el9uI3DeexSikEoQCNePRxcHvq7ImiYWlOz9BvLZQYb/pd54
CJ7EUqVhiOzHk31BXr54QVy4dt7T2anXWXadCxp/Q+i+C+smnFPpnfrfNUU2a8qC2QYW1r/UnQJv
kvt3keHQ95+ry/QNQ3UG2rqEU2gwpgnAtEW5k0le0aMV8Kkl0dxU7HUUYfoUuV14qgW8KC8uD3VP
K3GdlsVlRrfudHPa+XVwQITInSUQVcB1tSjQ4q+k0q2b/HrLQGlyFxQvCv+rS5GsINU9ShErbYup
vOBCOOX+1Y7UFM5wjlqXsB7oY7SYwI1f48bdTjtDPC5qBsFsypHWcpsLZGVxqeNsH1NsqznFdY1W
kb8QCfM43qxHou3QBlv6xUUX8GEXc3HCjK2LPneYcMMNADnNT4uqh67MD5AwO0ZDZGCwwssWiHw7
LM5HRciZZvFM2WkwecvkzVSShnuC67zhlQ/IzXLkoBGHHXmpa9eTTzufVuXoYyxBVoYrCaGP4oLP
pXZeWianKeg+3nA8cphfwr64PjMNWg58th+BWJbUGvSgZOlf26R2KUKEeAk5GZEKN6aKgDsvAgVT
JbqM1rJ5Yn6lGcvFByz2qv8nHyN+NRvXzIR/TAOvxym0mFEtXQsHsk6gAaQBavDtLJtopbfyLlH4
8g82zoZxc9KnMV9tLM3o6qASd8un7piVqFzkEkq23grj/ftVxAipNzuTgwUO2Yfidj037ohQ/0Xo
NNMIN2BSEj1IfZ9m7Io5W01+cC6Th7fjtY8OKgBik0kKKHzp0UvNpSN2NxwxfDhmjZ3svy0r7qNK
K7ZClYtKmpgT7NbgN5iyu2Dij5QZHH85ZZEBz1owf4lJHmDoEkWupw7VMreT+0raRYlhOxMf8r5V
q9v9R6iNfxknjK9M6GEMnETnLFDzawezSVF4fjm1NrGRNAaCtCwk1CT5u0i6bThwYhVjXYsVvuWa
ac2CXza6WfYCLphAoDzSJVu12xNit00lVE0IG7yNChUG5jKI0gEnKP+U9ol08zoMwmjiWsPEFF+B
y8LldxAxw9Q7Q/SaT/hyCkBOqTrWMmTcV/HI+KwpnRBbXNeOkfbT4/MoHeKV9pGLlSAc25AM5Y7r
FJOK99Opgx+4x6pUtGegp3CRnC1BMsURmS1SHr/LgWqKL8okUjBigXGA2OrxzdJ9TB7Vd3Rg0ETq
kiieNJhOiU0PTPPaK9d4EHYMs4xkGu3K0rNdkSgAQlS1zIsIOmCHPZf7OYa1X2elxWrh10XSPc97
yyOZMPaCy3uSboGPbt0W0MN7NMiFuXXhTV/gTJK2xTYYF17KWBVEIV4SoPprpo/naska66CAKzS7
ZT/s10+0+oK5OpcoXDbR0PGd+cSeobya8GviR/40zzozxg5amfB1O5AwsIMNAhnTgE+GQhaUB9QP
07qMo3BjcwH5C3Ujdmxxprtqm9X6iUKBsUMEt/MagEohWWPr0N37wuymLcPmRWh5wV/2XlC4Y4Io
A5pJ7jHzNHWXRtUIdi72rV+T88BlW5q8e0+WWjoVmytdeMvRraY7mxrDXlRFLl1qssw9OUM6aHVw
tTo1T2P7Nx5dHozJ1L/oRm9cFl0ocqCVQ/K6OiWY6LSOgo8cDsDMDPWzKIilTXamKu1b2V3PGZhE
WFBaltBs9+qkCv9ktSV3p0UTYa15eaIRRiwSCnysPe/x8xHqWDpiBgAkIz4otj4UxaHkdyI+lfIb
/Azc64mYwoUr3VGe9IkgryA6yYOEwi3wOYnUwQ060dA7VdU+2b435CYIlivvrhpcBUBfBr66tGgW
wXgwY6U/ufzh/Nej8iYiAuZjebdAwDQoV9ShMeFoF3A8RBRE6vsc+NSF9n++/zWvdQIqE2k7z8nK
N/3M4QxdsBewDokoQEP97O6tJrthmaxByPKj7ZV4f3owbyUp654jmwg0Zw09Tv2byMZg9cMq3tEm
WTb360HSqXPuSWbc1qXDKlfVMBjPHocDrmnCABr8ZXJk0SSrhpK6RxqahJGoY4cnODhiX35AOtXl
v1b8tVKdkxRK40ESMbcwRza7v1o8637pJw3u0eHeemuuZf/1NhUCPSSZyYmZX6uiCyNgj1kpPo9L
Eo1BW2wZbrtpTqbtmgPq1w2q9IAY8zR6dDTxLod0LzoMcqvAMWJ/oZ0xT534wKNjY5c1mFGUr7x7
9GPjRYYy+H1xpwMs2c5n//jMGvBrx1TQezM+KuhBEltUhGp6c3/59GLfv8j+lcyeg1F8794DxNK8
a2ACl53llCBJdrSXGCMPJvP8azE3iBzI6Rea+vF8EOBUuuFQYlCZ+OBVs5deD78e2qsqe+7J+WgD
GXoh2anqlwBHZ6/MvqBfQux/uwN9Ywp/zVg+bDm43GclCLrHiO7Qaunrp/TXNsKI9a8FeLyE4mPY
NsDfOx9CqasWe1k5uq52hXsO3Xli+98SgjRluR/lYt498z4mGnkLHIwM+nWf8fZyhqT7CnwzK6of
jxINy47GkGg9QI8P8sqgAPLb+puh6iv+4fwn90xAVNBaVvJszCo1+Jv+xvP7u2kXuGw/IBfydttE
wUc3qbAWF19Fq66y0frd1whooTS/4BxSEKrreccrMq2mkEVjGkrSkMQwCm7zqwX6xhNoCaAQSW+E
U2vOkf4t/15FCLtnAJSdohfEneLgQqw6FQQ+0Tid+j+e2KP5ZhyofaZt5Wv1PSSJI2bBKYP/jrJk
XYsOUpVybptuKWImC8dsPsjIZ0OKunQzheVrEv+cTJ3SxcLpLhPkXRiJH8Pl2hUDcDUTLUoofH0d
sdD37hMRQqfYQqOMRNZJ+diy2iOkogLtKIjmXsRsar/mkmSTCI9GpLRUKibB6bYrm3GHhvFCNWHm
/WvXlvucOhGjznXYLnme1/i4zon2G7/pqjQgVqZrZho0eaxgPx+BBGxHgyWfls09yFOtJdlEioV7
LIZnJvxDJlIyCktgDXau0uZR77lqGpFSt0o9Emc4sKPNEClvQJ1K4nQdRsVRrDdlOTJYves8dsKe
nioFCINCp+A1hpNzK2RD+vKaYPB0i2vwXNSqLbLf1c1My1c7cJ9xblJFeEdoh9uSfAUeLAwepSsv
UMu2xR6zJc8aqv1Hta/6MYj9oK2G6rczgPO9B6xD1DZOKay1bcSEjcFVOqtadg1XmgZD2lP3XJfQ
k/kqzRlxfbEMlkKwqvtMyKUDVw4gxL2+9XFUs3Axje/LEK7pPzGEB+IHZXTiSHIwphLSLKb4Hv3m
E7/33GzcMxts48PpV8b8co07TlJFzTbnPuBombsICFHxdr0DASD/AmVhs3XaGTfNNe1d59d2M/7V
xE1No2nxN4icSyvS52YtzlDZCV1ql9pvbEN1oEQuu0WQn9O9imqb/qRGMyjIhm8d6DrCcaRzvl0T
Lq1MgXKbdw8Z/zG83wbi5RTXSp7zBUn6G/s6lWFDR3y+X6ntfIFELibcn3+4lzNcRyDTeISeibm0
Ih7+0ZHSP9SemnL/gyXO3fln+Jpw4BdsrczRY5/pT5z/8LsKWBIHgUHpOY9T517GH2tmz9MIo7/a
oW7oEzWCF5FA12hrRvldhR4Pyq0cw6rBei5peJIhRFP6vUAG/vjb2/rQzuSVK7vGMoLPyIBshSLb
/ij9j3zdB3Tf4qRUh6xkQckswjHRqeFi7CbT9kapKC7YQOWLOK0KKRkCAxzcsDTOVPbygHyh6XZS
1L+qLfAzlL9eg5ulHb3ZvJ5XhRbu1tGH+waYoHlbkwllJ4//CtKEYP+hnE5UdMZdsY9Dw5+j5HUp
nJLd5Fp3bO2OskXHGPrRHW5a5oupXHbS7Pk0hXiehnT7Hmi4czdRYg06g4WyQKP9diR4irojLGyj
GfCMP+R3ocy3FPzJ+2BWUHSJqIVgCviXPmrNP4+Fpi2+VdhEk/uAdbjKYs7Q9o0af298wi8sIhHC
0FUKEYhDB0cA1J/NCbfTXzbWTJ8UZaQ7bYrtf3zkO6i+Blf//R/3RmAOWiaMTQwjsryuLpFE8tsa
LqN+yRpLBT2znqYQjaz0uJ/cvpZujYHCAHdXzaxdTCUT7hatFlelOyjmhlSP7RCADJKbynXKdFBp
Of/JWgbfp+v5gUXdB9RiauZoVnnDhNzyC/lUB45yY9UBoOQnNOGqtszAOqInPsaK1SV6KrpZmAA7
JDGyekx847axsic5yiBdMpeU1IiaSY3jfVrCFuxzMwWuTKFXokfx13O/mQHiboWpJYtDBNnHUbzM
q1MmL5Kuj9rYVIOMfsqElyrFf9U+LxNThDsC0bF63mK7FVRamuDxIDvm/3IaLrFGbkosl+z1PABF
7+htEse72ECOEjG9/c6/L/jjNNxmJ0jxMTlo4m/Fc+nR01K3z03cxKgjALHdk7DngTgw5s8uNnft
V5jyjwjV2MNN0Vj+kvRz1D7sEzjN+au+Ep/CY7XcAd+srnzFHhmYIOBRrPs1ZwBMPHQlJ+xTo/Y/
yEVCwzFzOi/fqO1csyibnWiMzlf1DBBGOyNqmUZCbbWN2mYAICPLwcdWdbRAYBes5fxqPDgNMr0g
PHu5Yo49QghkeoO9xeHh2AhvcxtRU3Kl0UYZLySqRbygsC3ihf6rDpMovDbp61BlzLGPCV52Tzd5
CPgioVNr5u+TSM7jl7k2AH5NIKrSCN6uSAwEhh5PLhK2pj5bXOqsX1o8kwUI/xERiILwQ9omOsCj
I2UN07ntlLEUxYFsFQyqc+UHiaWxhSgK8rACB8ZC1ThbsM4fUiS8kLYwb3x20NGd+bNoTs/L/Rbt
aG0IBFmYg8HWXfEZqMHm0OeDadS7818hHFswnkM+Ary1YVJZs4Y9ov9p/z6Y6fvUDZR/L3RR+MbV
OHKjn3RJLAQReQJ+qs2sKGy4uw8myqbSAR7evE7uzr+DTPxUvYszQ6Hsym9tRJV19sEyoyMyhdGt
jUSfvDoCu/nViE2poU1hfYhANJEyuZkYSljqQl2gCQJu0nSMTNFuoyEauK3XHirIEdUze0Kcxp1D
xijKc7G3Fr9F2IvoSc7061ZCVkuhBR9OkJ1+bqZnOVaU5PRkCvRJpKtBWTcjWQ9hhyF7NgNghCw7
O0zf39znP369D5B5gt20gQ+hcFNAUBXqYnpbZTSKik2HvmmKa5n9JwhrcOkfi0I1ZXxI68sVFF1i
+6BnCGG6CUtLIpduu+UlbAUshzw6MT/UFv3iivfcobIF+uOPPBWyz7r9S8XjNEv311YpVXzyiLHb
dVDpsVWxNYxWZIxXfimg/JMoI8lvU9lxIMCEtZDO/JcP1lqS4mIy5Psl12gXw5Pa3xP0Mdv1gAhb
f3nQIkemg26nDIgv6qR2gn1e5/EL7fUvTDmyVSQwYkKzx8aRPjsm2uxznbN5TgkHESzassvMq9PH
t8DVpwU0zsLhfwOZRVmEGwlAAFqkMvCLM8FXHoxgOUlylQHeWWgi/0575S3OHkyAtxavR7AMOEVG
6N6X+emrrkHcIjVL19okroZD4kHiH02HTR4pw0T6v3qiHbtj8dbDY9G3SzVVBq3EkE1Sdqwo2Guy
0VrTQKTwK4ntxeKlaLGNx6iFhk+3Oi71btXig851fGxAzGWqkhBgao3W/KHqoMxe1wgqYP7BAJId
XSqpyT9jl/kLuFA47Ew0jKW7xSdegzljttLxVC78IEmRPnV0wgkJ4/DIhqyGRGakRO/o0G/inlbX
I1ZC+jifqlgpq6eEN6vOe02qJRjo91s0pOAHLpATN+Re96k2EDKWT6TT6Ld3VDcqN2PnFhZNROC6
szAOjW/8zbCcu9wevPqW8rt1nstBlSUHvs8sV+hJ4uixXfuAntW3UwVSVJtaSjOQrg+48ACP2XXl
sd7wOy3MpnCDjzkyuCO6pbrIMa9xvZX1eWPo9a8D0QANM63y88Vo9Kn39AJOQqkd87KJ5BqlYndm
JeeMFUeKXD1Gd+dMgH+efckts/jf9qTZtNztHtP+xtmn7tRJmygL1TQojvXc36wm7InXTh+o53gq
2tz6FBy6XYJZs+mntR7AAPNI7Uwwovnt2a6qy7tG17+DU2EcX6exTjbHEGbXgoVFihCaQW7DT6n/
Bo4LQ0/KKc2Kn51HLccHazDiNW404fm6BryoWn6W9xvIX0cmOt/JDZEr/vDE667u+6yuPeLP3vWx
k1iPKydnhdDq8+6djN4E8k1KvrLNa5wRfMxIFrgquoP6W5IDYgj517AO4X3smf7SzAV3WAo4y26c
fj6hrJQgeDCTLI5XUQSC7cnLFcQea9I7T7pQqOjcckob6OQCst20yLnVfpL9GAM0ithwIdprEi7q
fKd8aMFqicVnJhpmWUv0/eGJ7rPxR9/Bgl+8zDg0i3yTtO8bMouIH08ZtdFQIXSw1DB1gak0B1hz
rRIxd1rf3QDT2sFFVlppEaRpencTQnSOXYB5dDOGWKg9F/4YCm+D1vVpGVaYi8sNAuhMeQ2/vulN
7YCNGXv95bVouOrI0pvq2JspNV/tylYb1+cSdib6HoxMFhnTfiDpv+5vknj4mxUnp56bCnU8jLbR
yDYAJQ7RIhbx5NGZwvu8aB6uNFEAzh1w9yT5m9amBYJokJ2y8OYhH435u2JLQDkowqm1VK69MXKl
/AdSYRpGm3BwURrZrKNTy2GaGQfjL0MWGXQ4fJb1/IIu7fd43YfQ+Qo6u3UL545mJc+nQm6/uF2Z
LloHPm2D3Vao0Ljt82avYcF0o2S9yZCT/s5bd9iVal1RTMA/VjSTTqOMabFeglFz7j6gzezD7qJK
Js15ihN2YCy0ifkfmM5VEAG9N2fLwd088WrtxzU9pdTeZ5L3V58pW1th1EXJxefPSoqnbfIjZcrC
2JucC00nYZExyMMGmGlPLMXlVNJbKNFinr0/CZNUCX5Mgi7bOpOHbSBbfeKS6nrNl1Q5Q5tDWgOm
e4JfpklndnPKK1PKS1NKVm5pRknNUjd7RTzf85KipPU5rdUDEtmbq8tidMROxVRZEZzhbTKNPTr1
eSm+14/8+6731akoE5CvNsoDgDiX1Wnkld9AobucrV1g0k76X/82PXoDjXrzYE98GKfQGE2IyPQ0
fotFUZ9CvJFbtS6g51BnKKk1SUFw1FKmhNg9e1EtikWP+J2oc/2kUwEv0Yt5wT2e94GW2yf7D2VH
6d13DUsD2g/HUt2doTMOoJPlK9lpVkybtWfYmUhEmt07ejfTqm0fRHebD0c0v/o3Qm/enjjViFzw
L5Bpu8DeYJwhBKr/nvRbdn1ad7Fa3KcAH6ZRVUbaWMu6mK5aRkngVfh/hbh6Q+Pcyeas/ZapbS4I
6kSPBfbwcoQP0Ubo35O9roy3k+FrdLbykMRIhvZBqgV3phRk7GzvgvGBtTyA5Q8vvru6f+tPr2LR
YRPp6ecYvZsJrVzyPXyX4+OpV9frEKJ2sRi59giSZcG9JlT5TJm+wUH3UI//EiT4Vab6iNkbXsnK
48XOfDsmkNesYt7Xnvzg9zAulYQzBtlOsxk3qqNf5QPHMl81tZpvJwpzeQpd6iuc1jm56EFkGBJU
2yd2qJ1fsteVuQt7NYQnzqwMyD/3tj44DGeZcXhiO4a/zNc5Dtr+Ezm6hAu9hKHdtDpXzYEHJSYZ
HR1PjZ5ZO6UDNqH6nZ0xpa+95ys/mQGVDtAkvfRnquOByC51W/INkt6tPeFqUxF3jGXivEtYT95w
lzC+9azM3CmkK6LIdudlZ88VrlAnCpMKJd/+dZzwmw+kvy+28N+LoRaWG/g4xBWCSA538tofSVZ4
Hj8uScJm1M11p4zfgF0f26ZIvOHo/jXCEM1Pk3Db+WkA3PYVb2y74zbgXPEgdDF9GyisxBwYM8b4
/OGH/bzLHt8rdaS9sK8FkG02ItkAzAuAavoyrgd2fYZpUiSGgQWjB7Z3P5dMsVUSamv/hwG5Yz8V
4gIXVqTKTyjuyinQiQhvX9S4da5IXKWn8zSoSWSpv9mJsGP584p2zusrvX0wQfwSEpiuv3a+z4O/
ymuFaj9yak1vYJf6zmLD3KbZO3BNHFfMxD3at/sZ9pq3MoB8Ct4I9++kZP7c+ty4j54kiPiNFPP2
LsT4ALz6whqAI3wJpdyk4j6ZD2mFa8qYPwA90Ow7sCjEFiNs1NMGNoHG+iZeT2rpEoX+/PzV7xiq
oLN/mlUuOtlR+ahaggjAxMZMYmZyMN4IJ1qm/ddh0tkxJpvXhDNk9Fh8VSnhcz5tjpcYkR1+ec1N
Rjgewll5NJKNZmqJyBbnz07q2pRHnrCe64xbEEC20Pl5hZFFAkuSfJdSRQtbdEOCKrCwtyWa8tiY
Gei7AJB8iGO62OMC3cDjl/Wu5NcXOJbp8U2a/Y9fj5bSMPigd9CzAfRrup8cCCSQtETpT+IIc07M
3p+6im1TzCr8XfvrwFVHj7sv1wLU/59IX/F4JCF5qBq7qkXh3rSn7x6fNGM99eRdMhxFZZYb5V5A
bxghaz3ag1ImrOjZ+UGLKwpsBEccuvT9E8gFr6i/SbxHGOhINLZ1mHDrSZ5q94Vb9P8oqCrxYdAU
l7TNbKYrmkuyWe1ieDu9tqHasPAQ5zlPlwnZBXOqQsADKwdyR1Q0RVjfvpgt0JNIUzMyINqLcgdw
DnTUJ3WC1I7+smG8D81/dL4WO+3mcrUN5ooHQyGIJj9VPw1Ce1iE0bAZYGMdJYiUImStnEqBFgnb
Ib4kisseBN2v7BteHlnIXJOhBY9eJUvlp5O7opmHhkErzK28isJyLxnkQIeYfhQ6uu2ScTx7cNfu
vKoJmqSSwXcAyYxPZBfEbPkYpp6q2nX2bD74hSUnnK0VaJJfZm3V7XiiX4D47aoIX5gbvewWIEF3
KS/EwQHwQMDaMnrJA10sZVwN/D9xXxz4BhFdC219I+6Up3VMCrXqWrvxBZ2DrCO5QNHpRcy6HHyE
z4nlwG9SjnRuS409zdqupVlIHNd9wr/iU1Absb+sy+OAPuR+GA2CJ35Ndzd4wmdBQFSlElUPX17T
OJn1W2lGEyq9O4DXC5bSMOPpWjyP1ATGLBtYf+sh6l0LV55UQaRqt5G0EaiI4ZzNxqMK73aQLl89
XCG0/v2ohfUDbo5NwA3ZwLBFepbfuTE4CJNqO8bgKOzfblstBOW4LyPqlStWgChzzXMYZPhpn56p
6chJGLG9OPe8vFyDk3X68TmBfX7x9IYmHwgKQ6/v89B3MX4sZPYDvI3/0xOnCcOzhICnHuB/ZWlw
N8TnCpifgyWVjtdy9WNK5IE8j6rc5LvSXPMKpCmzwo2X8IBrYkn4RrJUEaG9b3Sj8pquJg+yUG8N
tfi26NylvfEsgi0Boesre9Qh0aLb+4xBU6UJkZZ5ltZIPScFrWVvMeQcxEfiNSIhNXJwtmbWhDA1
MLSE6d4yOnqp3f8pjUVsUOYiHAeAlgJORyNgY0NrgrxBrw1DtWrfy24zeBCSXpZ6EiD0aPRhdVw7
xc1rcT6XklScQxm0Sn+Fykh5yMx2yNjFFIjpB8t/7Wz0gL6GcFAZiDeW0yo0NI+2Ex2kHQ7cN64j
MN323pncW7CC3GdLJyZuhn91GgZyDH1B3+nq1KRpfeTYL0Iz3/xBtDghN5MSNz0BUzAu+6i1YjRM
sZjH3ClZP5mDh5t71vLaKz13vh0QoOPzorBwoyTf4bed7P+JywtHyVhy+6nxkEUUHpu7+BsrqoHR
R8bbM1VeYKZNq+0GhC0meyiCfy1MnAH2aUe3XSs7EmfSYepU8Ev7S8xxQN9qI+WQWmC001Vlzzyx
T/efCXW0+shbvRkoFdANzpywOEoNIX/Xu1WAYpknklfu3I0G3tJXVOlSwAYQYjYL2B4ER+b8xSbR
YtmCmYe5JzVw2S8oKYIFRuAFg6TIPhuYSRVRl2pVG4PM7o72XS94fE1XdZwjuOt6JgvBHPkIVgiO
dzMqLpPhZH1APBV/HQC+SpTw1DNv/nmbkTyWLsyWQK4utCuPa9Xdn9WBQjbLm+IlIqvkuU1+UFxu
bQsccMhaYEc4wtXxGWf4gbeGeudsz4yVN85skl9cERoXCcfNs3Ou6PxQuju2aPGdFGeZcgT5NDZT
azPckF5cYBcEenShBHAS2ltrRzb5vXttAW/0Cj22zy4ka8Svk/rwco4crv8xMSmdSJJ/IpolEYAd
MvGi5BQCIS+4kEHlXsAsptP2kXpHp7uPI7RhgMWSaTVYf608czqAdbXuMd6wwGpvASDnjVXlLHfc
5sBc2NGiTaoBb3kCAj6ehVJCJ88neVxfogFP4FzZBug8KyhWZXGC32WhAUOCXK0r/5bgsuitAyA9
5Lp2wKxgcJRpFl8rhkBbtzdPUv0FFfsZ05y8mvUCH6Mrfw+NB83dhWG1TMUqKv9WYpNU3p8+3D6E
VfCe3uX9x/PsIAsQ7si3SEDumlvJyqH2NHK/rRMyheE5cSDEAQYtMs4XzcJgYfgpAsFNilel/S5h
0+nIQr3hyHZM8fNT46nHycHVt1m45Egcb4wgZFpcnEuRIXTPDdFSjAc22uHHXW/XowaiW7f103Cc
7U4Wys0UUHijfzxyq+UVQJHKpzFksKuoq5MpncYajrKVTNQpG76Hy8T6432CXgqLQPM7ciNYcSe/
rtVu2JoXOhufvosr6zxL5VZZwe6Nn4UQznnPlh7amVgeX7GJk7DZpqGQuFp1tSQZQhxaxQURD27h
3w3VTP6qA3lUGnB5o3QPNUQ9lOfB0I+QIpXntz8sTDSJyqcvWR6DTpHvuY7JVP8LLVFnec0u6Fmc
56aF8HIEO/ogxCI2yzQ6p/Q7CRgKiyShkod7Q+h78Z7KojxBEA7hfWUYYPlB+utvKsCAIE3YU6Uo
MRKObGjHKryjPHG09cAtcmtUAY1rPNanU0swtutssTEolyE7MXnTH6ivy6x3rkf63IIsmw1hVwCA
Q/3Z3ecy5x5iaKu7351t1SuwSyr6TQdM/IXYxmpWmEEcMv9kPrjzUgQKhLKqsT+tgIrWgkl8Vk6I
B6tN1EJeipaF+LN0f+ajH9Hr/HdUKa2D1Qyxve+EnxgMaXLEM3BcMWwOhCF1PkY02w1ZJG2ZAR11
oXybGs2hWiZmLR6Y8eCzalreKr/QXyyI/QGkm8JXBvYZAZZMU/hDMLmSs1o+tfRoTO4fPNneIL4k
xYrmGqqFIOQ89xkceshjCwk6E3LYHWcHN7cPOv32umYFscZlGqJTC1/5G+C1rF3zAICmvKl0MRTt
/VDSpiGhN1zFpCURSvlHPr1SZXyKAS7Nmj26Fbs2wln/Nnn7+ShCSrCufEspnAVY3QruoK7uwIS3
/8HPlMtd5/ScY+hmtdgVdIUkoISbmyIX62nQNdGIsAso+nqsK4hPXzKkj28WbsCN36egeUQqsmpg
MHL8giq9w0Qu/m43CnQTnPXHoZ8yP8cJoasDbiJ1ep6kaF3qwjuLzqThYB7vpckF+6jBZIa9cd3w
ckKa5rSY9l3n1bc1LObfzdESFmJQe5RKU1fc9EwkcwrGfw4ql1FEF0FdI5VgMK3QB00tEI+RQrNq
5akQ62y8GmDfsT8tCgDw/vUed6Gz4OOYlDBVHN7YZkJcyrIDm52HQK3hpM4DGpE0siw6Xhb8bU6V
TIUk+MP3iV2ZPsWmxBSTDN6mzJBIq15WUOnghu/3+wSEhLvRpdxqCETAq19Ze3V5K/cOSFAmiV08
ch9rC6g4bjBoQgARA/nGkkWeDOPaM6JF3l2oAbMl6waCaRzmO5xP46Prp8a/t5WzdpYXZ84RHE+y
KSK8npu7nPPwRVkikGkcUfbKtKhyhygauGCGflZNrN6mBbS9KIufnIIEkbb5uaHZPOHeTXAEdSpk
Uu0ENbKHBqEM9Eln5x55bb2IKow6IEH4mHHIE/ztGL9pdoOcen0RXaqzyVff2TgAK1hmx2C7z7UY
35jMxIsLxRJbgiqs/jUdgkocFZPClMv/b9Sy04hJPaw2cuTk0dVc7e7lvUXjF8Qpe1P/EhADsMUu
ND1Ft04AUtbLRn8bYf/althOHGqvT0zL9nH4yDS2GCDnIcBencVzT06xwpVkRszNm5wBCpovJeqk
sisLL4Ul/Wg28HsOHEkaAMhf6UCFE/69a701BkkqQAy2gWRbUoqrbnKv5cvZY95X2jN2MpAGwZ0S
KX4Xa0i7omUBIdUDnUGWyWts1th7gnhiB+1f84G0IzVu60coPKf8AslD8FFdZ15IuwgG/Y41TJmE
iDevCHM/SuRM0cNs0CgFLIR3THtbkY99BhD96iC54oKtJMnBxBEMXlBZMBAboSbLm62FemhP31Vp
V2eRumq9dl9Nn8kFQMygOL3GqckZJI6cv3ibCgS+f5TwRLqhz1F2qOHh0XoGAjVXQ+hljwEDFCRR
m8lyBFTvuZD/whRJXPWM65q5me8EyPiIJzcvOnRiK4Yn1BGxD5thYccwFf+WlSOfFZOO7e8AV6Ad
EsX64+oTH2NSdetspMJeJ3hD5PX/6CDdOH40x95Up+GQj+gODbYUPhwaU9SQn07xX6M8NhRrPQob
F24kZ0hpkJsCmAlVz1p9ranFk9vFAEKse7Ood4o3cCefswusYJOxe6XCx6tUE+/2C7eYRpiJwqhN
oGJjLsS7eT8sKG4E07tqNOaIGdVOhRRwHJ9N+KH+cQXX0BYVW/uknC2qBkCKAg5CHcxP4ApNHagr
EfN0lF9bYNyVdqvsheuMYd6RRO0/NTTTPtIQl3IfcYNkHRngiNCaYBE5v9Ojcbhqz6YuZlxUb7C2
GWfJ9hdz7Cx19n+X5x6eFMuGy9m8PR5/N/9Pf3fAh59YHqv63cdPs83NnTE9CQgPTPDf1pjbDjzq
f1oF1InwAtPY6w0GePaU6ndgvmDIWUl0SI86a7KOeJNa0LCNw+OAZUZqNGuZ13Rf60/1P2/Dx0lX
QFxJRkVxrKGfi7vUrMNwgvTsP/sQCA2HBLTDwvQn8LhTmhSTMEc5tiVxZTjU2KGPWyARrYBzhAhW
mOJqmpv7SlEh+zFKAw8czGaGHWCp43h6Wk/LYQ7J2MVlJWsvSi38nXWffA1IbpclzbiYFM4e2TXB
vN6qc2Dtc0MymUmvJ0+5KcbMZhGseuJ6sB9F75mLGrbF5ncUvVGhey3Sy6TrPQZ5Y4ayCXM0lZaw
ObRdgbjDcaFd1HBz2xLPzs96QtPEWbsvDPpWxSqjYQJOCNDPwrmItaGfUSJMql9NqsTrOZdp1krM
4AAPwsOMlBKOJfqtdFYSysyJbbJIn+schUvsDwU1AARjM76Ik65qE6BJHVomUw/7B6z8+n9pFvSp
pK5ZH/8NznwDpGYDWffI+RA+7TB5Y335POS9YYoKk9mVlARxMxhX1zl5Ztw7GhD6CZn0HJbuvzCu
zHxrWnPcEWmIhFIRwBIr8mOi2bGFozwoBBjLXBayqnrsMK/oLVJ0wW7Ww146YnTDGyeWTmI3PtiK
SUlk16+O/mXBEdblzSSJd+hCxBjmI6uAvWs5McYxC/4PAG2N27s2frCy0aWoVbDbTgwkS/H21tkO
1k4BI2SWNmYSDCyRWy9t/PBRCiDXiJ8HEp8eHq/T6nXUSdsVErVHaYn5uj+xi5BPAusOoHL9Y9Wk
QHiuBQZ1GUMV9A8zXIcFFyOys7NUr3oNp/u2TPEs+onLARZe9dKde68IvjBYvf3RvySUiq7PgeST
YzGxdItl2gOuQpCzTIc3Ujb0kSRe9ooQLBi6X+U++iNicYlQfhHGa/IPx8Wa8BND3TP/LJ3dGE2L
s5z/ucs79uiSo8pU2cONyTFJ/t0UV2fD6rCdpMfCT/ID67f/3q4xj1SL3s2v7aq74LT4I9sRWzAK
n+Yor0CGtbc1uf4YJLyZQ4Cy/5rBTK7CINzkXKy+SUmEvMDn2znuhDPeWuGdLDw5GbJJ/MLWEthZ
xczHIUbpLdOnqRQsZw875lwVsEprl+Khd9Nz5MRUXAHnrw/vja7AKbqMDyCnxGoWyQeBILx7GOsQ
rZTSbvJnl2z+ugs+t1efYxVLoNH49c7LQPZNzUwBjfyiqxpY2O+LeXyjTPgBWG324bpNgAHQXovg
8nG4BBDOlEUEGP5Gcl9bwgDUbThqqc3vwCOEDO3/hcfmirfQgmt+vHCifxM+W9TTbXUe8mofc3Gr
8uw4ZtSX12Q9+0FYXWYRfMSDd930nLvLltFxdAG7p0Hc49PVDSEa0j/CVyJgZe/t61CCvTHNn7LP
+I0iHnnA8g/gfL97yjqLkgqTV6in5OwMhagSIxq1a0OcI7D1tinxJxVo+rBGDtNW/tLwBrDUTx2Q
yIqg9fJ5Bks36NZkakklSyIS/3+PGmaWQ4vJRKock7F/fCOfgoXXnIRdlugfNSki8A2OU52tQETL
QKNB5NtbeaVkVe4vh3TfHD52iLpiXCkuiYf/H5ZNyTcfu9pJXXLt0z9+G+RAhouWY5sjeckBz/oR
HdCYitRaYcuuoUZZG7uYDzLzqLUPeQScNXge1UhRhgVa4Fxm69e0gzuXROwtFSfXa0xGz4a+9C3R
ITK8sWCP4foLWdvOQOQwLmaqAmtSNEZDgZOK7+Yt7IWTPe71AqQ9Dw79KvPeltk4xt723sXEBpxg
zH2zRnd4MGQC9Thh/adQP3i57nMM0c15Xe+78F60KCtXJKOV+81BHElcvYyIOfLrvXYlUvDaNhRU
26PE3IicdQq/SWX6jvVQFjk6bTizqRBrxkENTlZ+20xIfqFA+sPEMoW3WE6QRbKWryWPTmaphGGx
3DYb2ejLbBPsk38c7hN0InviBBAMaC9PQfdTBMqgdTbY8zqtllpZ0jd2Z23+3ujz4R3MQTKflcB9
SrkzyosZe+fXoo66t0UbzRWJ6a95tianHC+sdK5SyoicGrEcZKN01g5oNe4mq+zIaLgZRA0IKvgb
yjtv5M5a3zlHlj397FkA13kZRCwznaLvW1EWRp5rj3+uQtYGn+KI/+yucRTtdtz4vvrgmJtOb7E6
hMSlALPHuDFXR1wyNeyYKBLvpJYw0Ds7tQFOtbxiMTAXPSMyL4znPn8G2zlYFFk1MUyCbfXDZ+4w
coVZZLycb27NEJUx/kilnk1Z+lMp/ObUjjK+fzYYkS41t1PhI0wNFRS+PAGLY9t5tV0Ipe+BXhym
E3IIg4EmVDic9uXYi03AktmJFYiykaCOd819SckrxXNnqS7ztt3kNwaBWoWGvL6eTpGbjf/zoM3S
OngZAbrTM27v/PUqDN4xpDxgocbGuMqHMG9vSpslGqw0o0Tijz2GMG1Dowixeve0G2jQCKxt+yRg
aSaDngrrGoVVlN1G+fhmljBNs7rJRcUChaXJPkRq69H8NmvX15AKqKWEOR0/j9JmYV8aL7Ynnw4U
QUqGo7EepGPbzKE5Bi4AP8cLxh/yeyaBHKuGqPm+OyRUxgHI/CsIhgroEkqcQey7rCmjufIRvo/X
26Udcp1gVDYWdjih4kOPjXYo5xERdCRqCsmSgaDWLT9Gz33VfMl58t6RHJwhZa0O2BO8nExJe4w1
X4yvZ8sCFH4bp9uUDram89WcclJFWfw8jX93Sp/3OQR5/GFmP6UdKVZ1aKor62NFJL91u6d0ui8H
jW046tuD6sqil5AoOhBsKyrRyxb7LBJ/nT/xAf4RBpo3ESQPvKmEEZBALQe7bUhEANtpGxbxbQl9
nnYkK5hXVUV6L92EzC47XpjaQDeiu1+y6Z63YGSuP+MK+zIBwzcDmgrROMeMryzQ1MTGIgUrXmHU
4/laUALDOEJ4sk9CB5G/gfivwPjIvC1f01j0OF2BIP2qFRH8U8c++vqOsSLdLdwGMAY3fwn9Yi9Q
gupX00hYGuD7TKCy1nXRT7sBtTqUcQfz4QfiTnit4CuS8sf4Ei0D3vdY4Z9n9upytQ5PGeeMrtYY
XiWpIRqO+HCsse45WnEAuJGc0mBvLjHSM3AMHaiJC/OTbjK0By+U9s7m2pVe+xKUBh85WE72fPYF
l+rokN352A9rlr0Xk0Q1Yhgg4KkVWdMaSfoOeAoffje3uOJH5LwyIa2JGv2Otf9t9XaUUSrx1kpO
9OPN81+XGmReyF8rKovmhRvZ+IkdzoNOKg+plkF3eY5w2MA/J33lN5MwcJD75l0P0/ZwfRq6hvn3
FbsMD5TJdwBEUmWL/SAKo2CorjFtfDxHCUbG1iMw+9Hg5sUso3WKhEvcqmdAkg8mPEEy7uaSNC1G
izSbEuc4XiSpzSUGTq1tDv5+fXICkgyxuvgCeiO2nRaMclNPW+6I/LPlWDvc1ghHq+uqpZzH1Hnl
+io9ZnJ0isI+KfKlJ7MJlp81kGJcgJ6za7kTKc7dRTWJEuAUq5xO0hfYJ/rKDj8TzQCz4plmWQTM
VBgPppCyX9RctigI6Noq+h17MscoKD5fZwu6KXexZemsjeAxzxrEOo7qRsRz1oxEzQgeEKMXBPLi
hdgoJGMkIP4pZgzWmlsgOs2FJaYwToAmkZX66G27CFCVxTFjLC/aj+7V5z1qGXqjH/ReRU8Uj0ye
KIdQbAoZXcM+8lohwop1/iPK6RV7fbvX7JrR4uyQnK2kXfPtPKTkivUbguqNG7WA73ke76cm9cRZ
CVe9ro+W2zbogawN6+TwKSYnla9mTrDqmC83sKO5rJaUMgv6+pjAJXmCMK//7TfHBiImTgMAcQDc
WX40B86PPsICv7kjccemdbskp4lfRx8dJnbzsn3H6pD2j/0xG0v0oGwRsyJGmLDq2apt/G3gcr47
2/XTFSW4hkUkx5zSdFZxLDWm0hvvHsybFBSKddSPw6tk5KG6oOLAdh0Vv/q+WC+RjWCXlWRXfM3A
gd3d2qVj8E/V4XVPp6a4mGHnnzdgsLirTCIyHdbbPfDK1KlfJsVVSdjWhYtFw2m3UjbFePgRtF2j
IJv3VL7Trtpf10hmUS4UsgAwQ0+7l5i4eMvlnfZG0TYIMV07ktNURX60r9TnILzk/O6OCLkJ65OX
zA1ymj/+aDW/srsKetCmW2kNcJgDJzowT/VWZ8/hzJzJEU0vEl2HuU/KvjHBLfPVDegmyx6i/Q0P
HvjsqJES9IdJXNBMWfZzxSo8fKQHukrC2h7DHO5MYK/e1vIQfd2QVfcHZa0oHI2IuN+BjRueJ15H
kWD188lPKL+ISAq+hic2Tr4AymRNCMVORilyVToYtIMvAySjyu+kK2hIZtyuhdx3dLZi0QojTNEp
VWq4c4fDFUpX/8MlNxKFvKPcyGomgZHj+KS2pOau2Tm1upz5UIRVaNo48RsAY+fbd5mXq9L0Y+ur
Xnve9fY42gAKe2YOaAbHUPp+PRd4Vl/GJ+0s7nBUeQ9TpgsRivLmvPxZusmvcmQJMRQVv3SZHjA+
CcpF/nptm+6mCyRjSxi0wKlmS/e3eJ9Q3VT9Yx+a9411nn6WoR1xpqwE+yxHCNHb7StNogjG9cE2
o55/Nf7sgJTvE7baQlnrRQvYAAQSTAkGq4IOpycWZIxFtrBbBgkINVNrNlwKhOrkw2LH+4JnPitt
lbbio20YVs+kCPP0BUXtUKOucnp1O60QJPAvYVs427TEKZsORk7QxlqKp+P/WhJzbs0KLAlOIt5A
mSGhl4FhR7MnqxAZc9hVkqmDhD1DgZiRLwmn4rFRH6VLvWh0Yi0wmRIWhXzJc2Wvnv24zAVKZegp
A5W/pfrV/Q9dpZsP4YY/ioCRq8TOVALPQKWOcbUhQtSdXtE2UOJWiWoz7NyHO6K5S+WKzk7dke8T
7aCgC/UqJLIWfpA1WORxzPQku0mPQpBlaLvZYy4/YXXLgcodaPTLoqzWLCHQg8EDPVCPblnjivuj
yKJcxKfTulryWhzjYnpimAdoDYn+FRKGNMgg7N7wgtp49EoqxTrdgssoKB3n+joyQIMSGbd+8LXo
wI9dAqvNcAbPPUpBjUNoW5ndGQk6ZN5YZSJOme4gAeSH74AY0i3rTvBXd85JPqwH4LZ1VjxeSb56
PUoHbJDdbZ6p+T9IyhWBkS4ciBgm8Z7i3IwCER6Ypk1g5mVZUXKALGg5fUBeAxZU6oWvFFLLvGkl
QSlIwtGXjwYk0nlO2uegoPZtTROsrmEqXnj1RgTlzlSLSQKw6d0aThuRJt8paspyM1L2X7S9N5Gg
83/vwlfrdqqB0bIw8nTbXdyK4SgJkYrxVDKQHMLKrYA2JsxXEgnlrM34Ac9W0FDJNNQTZrT/PG6T
4naek84paRKiaOdum488irbKlINdQYJCwREO6N16oem7kin6saEvjb617DlEVnjGeX3GbaLD9+Fe
lyZaH0JsPSFNAjJ61cUr2qzWa0V9WmgY4BI9cSpGqkOJKOnRAyKiZy95oxuj8oq46Mukiyshk1v1
XbJsvkOKeL1cjcHh6ASnfTEpQTTkXNog5FsaiLvSvy0lZDa4Wioboi2iUqknrL1P/uFT0qUfk1c4
BFZKsXBR3zDVjylQhG98dgTVhFRvrdI1uTmSjsL8tm4lnMJ4u4aDoYHPOAqggbWprgim5OYPdcFV
V/1byWWBZxg4KPdMFq+LE8cKT7AOB6VTmqDVrQNYqqTjYOLDOXMfWWKhYi6064SQQwBiiSChnrro
Yhbhp3NXiGPhcx7QnsY3j7pbQJ3p5o9e0CeWRTHoAiRQouZSIRmCBvmaZACKimje+2bKOiDTnEMj
7qfX/deOzzUqcKoKCPd1w7O0wMJAUuq46xvizcmFSoQruq5zp15XHX2haP9SMhtyg7OCX9SsMeTJ
VxNpcH6VNuz73k/mrGQN1bDUz7pSoev6FeDopCEEJj6nLI13H0teMVOamVGsQ1BdqrXWDbOvEK7P
JjZiQ+zYAJHk2DT8c4KEJRdxvfuNq1X/k93NSxsMcAeUp2rqgDv71kTum9IF6b+BUz23TW3bXfyJ
BWumze6vEjdxjLeQbVvEdJz2wBN9MJoQaJj4to/AIZ0mMJOUQSJ9Se7zUXu3KIyZ4e7iV6j01EYu
wXL3ST0VfeFId9DlxEhLYDVTdAmb+LaSewUHMIZapI2t5pFE9WIuiR2twYr7MbDww/mIkgR4qy90
ZEY068h2Bz2AAczvUw+da8nL4Q+kcH2WWlerl1eV7EGNDpAd1ZXraaBq471hru38nHCUAp1zFfA8
854c6uM2m0TYh/0Z/6quvwEuudIxgq2tQVNvVZmcOCGgYiu2xuS9cmKUacHBIqfRtIvYW2CIrsnl
7cO6yV6KiszOCaWXNcSDNef72dYmiGNHwupZMe7ZcXhQ2rKLELynfhKPxGL/nbWWs1Li2UqEzrpq
j5qCNwNCj53W9TjEOwjmZQExMn/RrdLUzA1UyOdj8yAxDUsNCAJJoU9imJggZxjho5FjzTirrgHU
Jz+A2QR4TDUnf0am1C2+Kjx6W8yacQprhKByzWZ1ZW9jS259dwIbvCIigehpmJJuezSLS3mLCx2f
rC2UEeI94fqJ+ORHWhHMYzd/J+eLcq7kqL1dZnA31+uf7oCPb7jUC4nKrjVRR4cvDB/S9y+0Sfy7
v+Sv06XSXANAYEEqs4vpBCybZ6eZKmmjnS2jj69WL5TvosrYAOIMk6YqoS+pEpQGZa2ZY8JEjD+S
YjCvaHTDFMpSjK5z7TveRyQpOa33L4tWS34eDa5T5wi0kcKZ9/2tHFljtvTEgU8cYLcp9G4wBmEy
Gw36BA/uWHJ9EpkMlANrXrFNwqRmbhlsaQFO6DUdkoA6+tqMCOnAFkfO9eEB5OpszxuCkv5eSTWc
Z5e72khtWITz+S02W7ikizLnV50DUsuUlS080SKeaUIIjv0hx/HkMkkO7noIW2gPqVPnZecbEM0q
xHm9JbSveJay1gXixj30Ekjw+hxUjphZqZe8Zkpr85HavrF/wgPddrMz/fQ+06d8NAQ0YeWjuDz2
fBKGtVr0r3HM1NROFAvcphlFHuqV+xvE0PmWqGr6624il2rwi7bUsJRTsiI229YC6C1s1XLD75Se
RP9/UY/hU0g251FV+urVc5RfmUBFxRJnboqSJ1ZKsOAhJ28Ll50DtHgb9FplDYJOQxgdvf4i73VH
Y1EoHgCmkikJi4aEq6ACk0pJ3M0rOsQ61DVhApzC26+tET1EcrAGuGE61PgJz+yr5F4glIgqSOz8
qqcrHSMVVnOZ17iuhLujs4evu5B90nPDtWEXSHijxFsRAEpAZDxZP/VLWE2kvRYbBUcRpeKigByK
SirHo3iMnVsgT3Ct9gKwY3KHk1jFCXBaxFxUQl5Bk5+zGgC2Jl4ucFI6OmLXEcYBMLXDKGPpIBv3
Xp1CHcwp3wgb6ZKRiKorVGe8C3m511lBb+EcCHz9Lwel5FOdP+jU+hWQmKSQV0DlGY9AAJD1FY0C
itPsDwl79XsN/A//8Wr9CeCJ4nslXLDTJfr3fqAyyZSeVn+dgZYKXZyqbWuKbkGVgKBJPrXe/KHN
hRbEcei06DAIjrtAKQC5e52jxA7vh3ABB+BIP9lWahBh/UcLHdCtAhLGS3CZVdYqBRb/IS27V+07
8OmulmMOxmxsbbCVg9yx2q3GAiMX+VcAPLTBQARpIZzF8nExt483lOhRJU2Em/a63iJWSF2hdDlc
+h9R2E0x47uAMUhCn2zh9t9GYXm4DpGcghATZNP6Kqr8SlpjwARAtf+eXKGdwkp2yjOaCbhEsNml
BXs1uqQLbyhJ6zKKZ0CfdbjSK1bmZv6RScBXm2JyR4dga3DBPCDwzA0FXPWBhrO7ED0f74HFWT62
pqICp2CPIycM6g9UVfX8T344JdPQRHUVxx2rfnj0TfuYkQJKX4FamdUlgmKk8pmiw99o8AvIPNcg
JOK2OJgEeUx0oK6lHFf73dhRgqumKmGjkeU0Tay0gWAS9PYfLVN1/YRAX0Jor8wiiCSpJoPJXEZf
jvNvXQoqpOrpJ2u1vACYfTyxz7VRKLuSTRLd5dQgwGCOvhNmjyIy9Qd1QkT9c24oFy5K6wNbqiAX
aEi7bImcSuyU+tK0THS/jrGMLMQelsYPWL9O3HfVbD7X/5HlFlDib5eg/zU4CvpSwcOf+ntKewvC
p+RtHSxUiFBgb6UA53G0QKzAiZ2kHFKE9SBVve/dAXHoXL+cxzMz6/itr2le9rUOHuhtgWBBUAtD
hGsO56gOkiShf/zEQVF+zVNVdBJ8gSkw6TtZyR2KV33E771BaxYvAf+3b+YQ4ClxLYuutGqfhT+I
G4HUR6vKedsJN2KqEGj2XMDAnDWmsYDq2EoI5oDJCqA8EjY2TsrSJwJw+wLghMYpdOIhsk4T+LFs
krdIeWvMdMjaVelEXveGGmxSXnKmlQ1ujtql56W+uXSNyrYxcSfOyuqJukGR16TQ8JUzsbwN7ZDk
EKT6Xp2Oo9YfJ6cLKOHgDYQZ4DD2n+YD60ZjdT6w/uKX1krbwSpFeRJUZYDOM2ZDlWUoYr8wr69p
EcDZo68HQ654Y8ZioqTr2GifdF12jvbJMYML5UwZCS2bYlv6yO5MWOogYuR1yqnOH9zhC3zllWov
06Hbnpa0coHImIXGvrVVU1dej9cS9rL1G+z+r9voRKpuuvPFUA5Xy0Oqg9vHxzJMrg1oIkHt4C9h
bQLiAotXuCY/K39CIrrSyrV/pruxwfkBT2Kg0fLsIcKhMPHgKpPqE7KYimLO4xQcMO/yE9jl6pCQ
2qoqIhgHh76y853HOLjdd5j8IpKZX5SM+XJCZKSNvPYm/7nxqhClISKIINGO4KHnaon+UYhDWoCD
ccewxesBCqSgcQKZOzqNWTkQ+MXLZz6jKOxFZuHcnTbSIW9IvcCbTzLgR+PxBnOEtjHTGgC4iUa7
BxahbLR0vCX8BqlsF0YNlWjwKujSvJl+gWay5psd7MY1adCe8GtCtKPB2dHAziQuT90eInf9hm2p
nbdLTlMXH4DCcdJu9RfzxshfJjtCluT4ygsPWZoUkUARsIg4d617/16sik+jG4cLD67zlK3pc6Qq
NzKxg+/TRSZLPVWcMHApqogW/dX0nW16JLrRq9c0CzMwOPK7XFWlGTJsQUpBdNbXuBFhqALE2lt+
2TqbW/fCetVvbb0mPixBZVNVKrGQIek0Q05yHDnBR4lkLzv9SbtqGdLDilK6cWhl592CTXfk/qYQ
54kTVyHQWSjPUnNwnSZkk7nuHGhPZMzjqOn4fWGy2xp83d5qfr7rAA8aspFbrGZW5UpzO9+YClee
FzSjc/H7BYsmtB0KcXRJ3aOLTmBWwxJSmENCrSx7eNb41xEkvYyQZvj1HNt5k3VO9ZMF1T/MgW6A
plxVww25Avc+HsOnQV+pTFdd+1nlcAomDhbAtpDYTFIRjMk6mM4KQDolOel4bclJIHoLb8+FXruk
AGCSfxztht9M0SnRQ+0+5kRaNtBrAx7iIJ3vJfDPsA62jDoUhrnkFmI8X7Uy1A8luYkTJnZYR/3M
RDYn2/BdqQ9UVp8i/Yjgo1brSyfVyn8qxndZ7qH06TTxeGgfZQsbtIlg0G13HyGdREcftzQ8jGFj
N0WwB3pv5reNPUFrdbx27O7rO9yvCiY6W7K6fQzdiR8Fl35+KBaR4Fp3aUYhzspLE7E5rukGkEG/
YegoOxQwcW+IuQZixSSgPyBPp4bCkErZWiASJTmlg+cl8thYSvdLeR5Dn5tsAcmg7m5s9uN40bTF
Ai89jpKSt3zPSjoOKGfSh3n/4FYL+UCnJcjrpq/+k2N5N1KbsD67eHz8w07sSF/4f+tNXaqbEEFJ
DKWUNd1a4B3b/jLA2h/DCxNlcNXer1fbHnYtrHGCmFO9qgnybBcN6FaAPnC7n1E1W1tMKN4rOaGv
SeZb2CKRxKoCy/AtsaW+u4Gmaz0BG7pvnYLMAS9yeY8Z9WBqyy7r4mjezcRvxHgEQ5KsOJrs4fmE
xKdaQN+aei69jZLu4dn8RMuNVd7AT2/k/dfYHW5numIw9UjF4eamkFmiI+pCZ8ULTGxI6a7wEUT8
hlKhNRlwHPGNDUDzgrv7RP3iLx+5/1RKDif6vj8dV+l1QBUo8LKadxQykeLQg/D0K61vwJZKrHap
9LU9xPrftaV0XcgWlXyF9jKsxmB4zYCT9g8JG0C8p4DPLIwMTfWEZvb+y/g0mg3mQfiKvBvY3JVu
trdIeW9E4xrlHQKVH8HbAVkX3k+ERo3sHpHAgTi31i4EPdm2F8maqjgoNqPzUmZjfxOc+6aIpDli
mgxt/v2YIdVPdUF0axFu7CAZBMWcdlcUM//2zDItGtcYmKjxWShsHhocI+cPjqZ0XGW3qS9SUzOO
65KcYxIC44WUWw5Xi20O9YvIJ9gCV9HEWlSDmtlj/RwYwLS3T/deFzWlOr4YzQMcRA7LWYtT/NfU
Cu75huRKWFkp6AOqRoS8ltfmaldcPuBQmTf+0fXaFBtstfuIRuQDf6yz/lI4p1Yuy2zUAElhqG5D
s3QMbKIivUZmlEioO0wtM6Y4gr228JuuDTZ5PjbO7rUUrFtnR4pdstjuStlbic83LlBM/RFhAig8
2B/mhrkonVroW4B5qbH93MkAkZB4CbTyE6JxItdFUrFGIKoEmUsvhUccy7l890d96MzDMVqz4qOL
skFv8akQqctunRouXH77iaox8R0XIXNstaxHD6fwLs5SH5oN/CfB3JMtgWxaphYlzqO7WSzil90Y
4npw5/e+x9JKcRgRLJx6S8JeSq/BK5Y9iF79j1fCzhVDnyG/dCCF3cK9k5twlYtF3f7Wg6dk4h9q
EMszRzZ9iEqAk0U4jFXY5t9B+Y8KxVDHKHesJxwY8iiXGgoreTVJV2jl5uYIYgVYaWGsRc4n3mVn
uHdtfQPjuDJ19u6rfSIHCEaIr4La6e4B0fBGvqjlWpcbyulDxEDZJWLqfzdTAjoWxxHArSj2gNVv
cbHOQjHw65S9AFxQHS03N4AsWrAY9fkY4GeKcneELyKU7PGoyIhtDL3X/ossBuwcnuzA9DgFqTJK
3owvi0qv1g7hIyetpiwOuSm4akTqi1FlK8Bo98w3LQVlOYbAiRYToJP7hD6hX3l3BRWRSHhT5Br5
SOAN6A3Zm26T1nu9guLMBE/LNEPjoKvlW1VXw6cEHj+kJbO9dZkieFPi57di9Tr2/+e37ZMZTbZ7
5rdp+xIswYzEsz0ntlRfMkfeLihyeqNthLICfpeQ4FgFdrwzmoHme7fBg3TJ3cc/vvOIWJr1gsa6
CRklCmUTb3ADNpMrsFebgjV8uqmy3Vk+LLmV85DzNaE4FVbJAtUgDvNA1O+pDuufXMsgVb164Jmt
+oUZ121B2mou9q68tE4t1cqEG/vSkO/zttnoov1A1dTuskfwdL5o4JJgkahjAzVrogLrFJcYkroe
xQLo9BYGb5ZxATChp6/J/GD9EH6oA+ZgOgQS26noYd5LQ9nHwQsFBL19UUKE+5b40luYJ+Q24R6/
wMKTha9zgMMlucdQdzb6CpFU/vivwXflJSId2PzBeMnOeedzSbOoBLKPz7tHgJ5SvIuT0BUDh1FL
VQHHLIkOg4bdRx0RtloDszED6897ih8ss6gtVCanCQyqT6pfqPjykTZbfuniYqWWwun0FEZ1YgrM
zZsBLjCBTRPSwNohJJ4WND5/pxq+crMDfAzYvaxxaZ1+xR7pEKMKx8sEjOyTElgPsB9L1+v8KhCR
3UNIF98W1lQMFejx3sKMwrKBgWLWki0egNAm6Xk9aLPINXyEW0rDCwR4IgZPtaYPSsAaFM1tqV4L
TnjUjbSG6AOMzNiQ1r7QKQVmF6QpS+xrlITpjNI1n9BQJVqgo4J26+rwM6iujtUPo+vkLAqzucZG
ByI80YiQ09sZTsuiZWDv54oabz6DtgLcS2IF6piBBWc8J/XOV/bHpu1/3pXZm/qlY7+8/dng/Rr+
rxiMJmi1fZQT7YcHkU2coOEw1M3pnm4EWd38kNrLW4Qa5mpeLFKx0tMDPzPNntQ131iWQoyZXLsE
XK7Er05IpluX6noWukwMvIxDp3VYLdGDhNaFbdA0cHj1PiTCxpnhEDo6YcWHuObXq5xCVkAfLmZ/
4njfaN+8OBF18VFWbdrOut5GaErPycSc3+kywwRomxOg6wT7Xd3HN0n/1k2AQ0T8Kb3Hi8yZX5n1
pATVux+Ffy73cFkq21jehjkxqLQb0D0RmuLtsrSnqFPhLxz12aPLJRCcOQrjQpWZPMUagMq+k79k
9USAReVB0KNq7ApKB5c3alLwXPIkfLJg4plMEy6XAprJ9vEs9xpZ4JMqU3N5X2SB4UFuHmo63kKg
0Wv5Sc4eu+NJCiTuTms+ooks4uwBDi0QKVy5SperUT+qGOWYda7mTafCeq+OlyGp/HnoKU2/kbtE
2qI0OTMv1Gq4NbIYYodauTB/XWM630/vl1aLgTVj9LqH3jn+wM5V7aHAynOJ+T1xy4Uh6TfUsXrC
7PsiLYgNJKhSm8pIdlF/tBeH+U//FWPCTZcU67lCh2TAI4UBz94n464+M3+GXd0B5ApWHGLA0tvf
QQzwyck+1McD10l1+F+YLqCe608OxIxPk7ONYg8TiPML6EZBWR0DcgppkFpNF2JbpE/c9uNygfb8
IwF6DaQmjyYOthwG5lSUg19mK8nY8XfRKh3y/z7SdIOQWBL0KB12yYPF+S5DNYt0EjmHzAAdr89u
BgX70IeByYdA5VD+nefvzG5araqtPBl51S+52z1rugwKdkLXWt5MLIJI3jDyh4vyAQou6+3fTpqw
UD+fGWOUPYFhTo1Ytmg7WuYtl729pD9TJIx7vLZR6SLyG3yW8TPj+ffsduPRqywfvyF9YdT0RAx6
d/ZlikVYSAlDH3FSLaG/DNJ6enkWnF9kkfjLqWdnIykKDQFnvdhxENsgcED3bB9qrPmJ/qcqOH0h
vyMT7axVZQnXuyvqbQ+lof9LiFhpt3HbQVY+9JtW4fLI75DC7R6d1rH7U70B6u6t3vwYikD/Q7xO
IEZgleOgPnbc+SoeR0IFbBccq5061u2N9mbFSgJE68MptL2q5s/ZWCwiJPG672bJkGBh0mtBtXbF
H8Q/xaO/5HNu10w0+dvUqtJK+6DFCFFnQfZvApDpwZqrbY5KEHuSH7ZfWajdkdqJY/C4Zmdd8WEJ
pUZXYoUD/0Jbh+Sjdj2jCFIyhBXxapIy9OnlvuMUVlXNKVmv328K3WG0rXtkx8O/dh3axn77cYKZ
3NPXxW0VBrc8KeczqwlGy4LOHoWfEKK/T8F4Q2oqR9ow0Qpd2++QH5meLhTKg3NQ1tFGrGXS0EkW
gyiMz3zHBryWRz2d8Tofj8UAHpS7g/7oJDHVvyCQyJn8WoUYgq+PZQHx5njbNGPqJB59Y7SGLAyE
IZyU6dsUKd4fvnxF4xfUBVgJueZGVeBJb8UgQ6np6ltIb2gDUUlWdPwSYynMosdMFn+F+gLdCIr7
mFs2AiSpiBQ5uwTZQ97xrAwpnh9vpdOJyqemVM2ajJqUjiTN+FVXFo/UhZy4j4vcet7A36jS+wUY
piH6T86lD1hOFcpSXafeGIIQ+5jMiQmHmQgvix8oPWKB7cyHq0qkWPPIEC3KK5oy/pazTXlMEKy8
7IDjQNxAwMnhsuLRK3CXjw4RBwyw92qpnU6oJBfjNjVzc5+tmCZUpmjUKQYjOIlmIf2WJLETpAFG
U+0wQFvC6mvF77MZeHugbH7D5bRL7oM63IkvkB6e8vPE56D9ckOADJRpAdMdBN35k+STLfygEVJK
YloYjAKwjrcLplCtHXdQGBVKW9ognDKGu6OTTPG/iUh8YNi+st3OyrjZPX3Az1zVAiPHyiBAtrP8
PhHXroJ3PCLHj9CFu3hZpHxwGWllwlU0CnUnahvwvAvcKkzUEvJDtxnOEKCF11zDh+ieO2cBSjtk
mQmb0itmK/yNQmNGvDWbIj1sxjZGBPzn48mG5S4KSujGXn6+d6sK3tMOcsRL/oqwtjILtr2XtM1G
jWKuLDMo4xOC/QamjskLHxWPmEJNFoK8/SwytLmihfJ9CsViP1MTlrSwDImLRXF0u89T6IDQ8PB3
kVX6T76HjISGOMU+/nnWUeTHRQMC57EGThLMYhYPVyrtxZEBtVVw2IyHiYFoTK4SdD+yu3poUloD
jvlevVcAczbgqtACxldyPXc/9MZIxImAAM6mow141X6vXS6gHGSHrDrU9Q8+bo2H6S6u72aDY1fC
L9DXu8B9iQuAVB84HIwE1lYKPP5uz0FwoXwndo3MqdZlDfNF0iW5IIf8SPa44NtGXlVYyBEsgZW3
8vqgCAIxvmTkdSqBUCYtH7CsT5FiJxzSUkqSqH9kfn/lMY/bWHYWGf0hEslU5ktXjX7HAnSL9/i/
R5eAp+wUj/0vagzJJXV/BJNN0kn47EUwpveByfHzolSwE9j5pil6zW1BJ5EqJtJdj2p+SbXf4eZ8
GoxYwhjVct3V0dIeqVrO3YUQs1xpFlvTwtc1ee+rvEP8fs4O5Er0zo3tGoSe9s+h6oQSKCus/nUM
9weWiEYV6veLRIK1yPa3gIgBHucJC1xG4LpsMjHTKTxj6+VDUBs6x4woKLMZ1irCOrvcV38200WK
AlklzkXyu7wbPsb4yb4qckkmoNiaW9MCvhdVVgLuu13+6yIeJLMlrs8bzQgN3eFXVzbmb9eF82dR
tE4CM4vDFQWycOAZp+JVynlWei8mu2zYsZwrBBwwIIhrGeZRxwflJHuE+kVNYB/KHdiUhGLfO0L3
l4e77BHe84wwJ1Pi663wCCufFUJfM52NNQQ1vR2KQbfDhm7GDDz6FGKDEM3Hz92pVcQ5GG9srnOq
k5vHyvZuTJW77Ma/lDPsOimq4R9YnqSNmhux1JCEsamVSDf138Hf1VMU47iVFl9GnLDiPv1VbsbD
R59pEweH/MGY5qYLbOQo17yMFhXL79qgs2c1StXauWJqDMSc6Ft/A0kBjgHZfbRUCKxcXNykMa2/
pzQNxr5pn12TEVtutwsRn2YLB1jHA/vC/kipolxiL/Hxl9uOk1p+ZFUwg/gxnt7IE+JOZL3cAUck
hFxkWmOPvJu4Wpx2KHhURkQU7oIBTSrqT3XxW4+OOB0Wpj11MfKji/h3jsRxXbBU4mtEtf7B4EhT
pTx+KE9Ob2Hv6Q9aVF3sL4WYBN1wERlu6EFW3QTcKAWpYGJa7qCST0BuOTT2l67U9srcuHRn6ED+
0BrN5NQZLEH+F/8ioNiLLCjpN1H9QKQolCN7Y7Q7vRHc9Nq/UIYFg74W89V60cUkjACgblUMVLUS
wImJ9LJfAQzQ5wibGoy1iW3aC2U0Q85Rq67ly6crlCFPJtUnJbU8xNI6syPqppUX75utDaMAGg88
OppibCtQ6ffQu72qPP8oqgVnz6JeK4t8JHIUPhOkpydOrxmaWfRDpar6AcDm9rwoISmw4gvkOJph
W3SNbfgwNKwSGjkhpSziYIb5KXKaeb2HXtShB4hm0YkBfw2TWaTJknJCZL2P8By4pNpGS59JTcxB
yHPOxg99BWOiE17d495TDa0NbSF5b9j8Ynaor4X57GfHdTVk/TIBEl201T+kzxtAwJ9rDUPfV6za
ij+aA75cpDCgmzWkceozC8vSPyBIm73DQq3C7brnXKN+FBXv/dmM1AUziO4OPB3epBT9Q0LMsz2X
n1HmA1Odl8JZQQaVH8TAodygRPbL7E8/bMCZh5C8Y16g3y6TFamH70b+05KoB6qxwB3wHU++OQcZ
QjKbJ+Q5pUfonOUX9aNQ0Aum6+lmEHx1VArNUAIoq/DCLbHCw0gHPgf9PvkEHAt7HfWOHRzMqrjz
BQ0Pb+SN3WWg3q1eDc4qpFgZdf7mSwHHalOyVOAcnnOSqkfexK6DWpxYn8lQDZeE46fjCYHKxRBv
8MU9lbpX3nfQJN/eeAa9VxYMZ9AGxh/4tvYj+B6XfGzC47hLofar0EOMMb0WJZKFhHHXiuz0dZEo
bWLfG+FsbB4tphxq4yeSHCbyrI3Zy+oO43KQMiK01hDu8oBJeje8+7MZZ4rL00bBCARncN+78V93
1EPH+O2KkygiOM5pEHZb4uSfdfbU+rEBwCD4r5qPb+7Wt5HB4bsJrXgXNQz4OE1mOjJ3I+Wee/Fs
B43usfTyJR8YfepoiwH30+EE7g4HE7I/WDkVNDVhArFOdVlKya1+jlGN6U2G8ilfkEafQu2TxckB
Myt+pkbT5S496vVOgtmTDSFZdm7dO3HUE62k0WKdZ4kgVqwuU1NIF0RBx6UfGKcdyawBO9nyyxe7
FnyOWZHMHZLJu7G+SVz1dXHTkXv0xc/mjY5Fgbr8dqmkJnoktpQ+sm1WLarBfd3stW5zny8vlXak
OkcYK0aI5CpeWodKnohfH/i55PmwBWi/FbQj4ST2/p+J5JkHt46AiPHS91BYB6N+7FlMHB2GxyNx
KtCKrKi6TN6s3MmgDvYezFxsUmL6fhEHTuaYDEHcTkWBHI0FV0/Mj5JdytTxI0nUC+uXRibpFMVE
jJfxWx8e9kqfraPe4cGRGw+vrRgmz6KAvDyPayIeNopw5MmqwVQ8zgtY9528ENo8U5f+E/ZnX9QO
yV0k0a1wCSANKM1BWXjpe7IjtVAgMXR1N36dpmHOLPvJSyBB7GkUSF+IYUnoDrGp+rUGypH03M+A
Jgw6aUu/4LdC+L/CM0VtFpaXGXSMSnPJPQh1rgVMIYQynyGJpjsDmLMGgtT+DV2qym7oTvFHshTK
p0HAerE4O/V1cPp8fKL/H94bDtOBqQyGJDve/JdpY1JLcIFdjQKt9wAEAceoSvTTyJ7Q1dthzU0p
qakIFcGlGETnIEwxLTxGwKf4JNR9OaOLGiVv6+pCP05F5MQ5o55/hLAW7HiphpumnavZ1AmSCcQz
EuEzBFeXUvRagrhDkgZ7pYhD1wcZYhkiFrZzki+449S2/quiJf9KndvrdGLLX4lqFxhfDPxr2mgz
cAEEZAlZ5JBtmE2kO7aA3MiFked74FqO2hGBfn7ugBzVk09z/ErSm45dpko/mkTYmaZv6Od9zFFY
wdlSelASooKRIUbuCe/AGJYMrGJWr5ICWFPoucKBHbKVjt2nchXA2ntefCTWqAmVqT9XVdVEWMoy
iIyFkwM4urs9XdA8UUzId6vQIm8a+e6wwCqr6W/M27zyklOkxWdMzUbcMg3VEIsi0BtXS54HRRyr
jT3frzFRY2WPih7OYjzNw8zG7RTIayEcX45RQwaqa+FAp36PVHTliEAGMzigku/WM+Od7Mt1SbWB
lvS0Ch5qP/a+iFB8SoOiD4AOkIshppdVQ+mGRF2QvvDGJ2r9tt8Hu8+3RaQWkBQt3hGFsRT+xcpE
nxSkfvu5kD5k7EAC15yZsWoSk/LrZafiA2tXFQ5myvmNrBsjCsuTXzGDY51DjynwmeoVPZtQQFYj
CPuGkSglGSiPdGnzLw2fx7g8ODCkzaWDBBlpIPnyciyBRzG/13VDGQlKGXAI4OnyEWQ0XIkYBmFl
ViLcdRAJAFzVLAuzPgjJ0SjAKl2SGRjCzqoCPzycwcuy4RlvChCVq5acj7aO0+bbhqRxbVeDvt/C
O3qN74tcs7+77eru1MD8JpoNca+tyyTxCocfd/oQ5tgRJFRl0wQXMRH+4mJyueiqhHdiO9sav8r8
P3RpyDT5uuDkR+7BG+8jNkskt7GJDwK7TZpuGUlUQcFnysqUr2Z+QiUiTyaJ+AKb1UidSf5cqQtX
gTpvid8p5maJvONV3puHT29yRcLPDQu06qTbgyemq/tKQsGE+2VeFYqwwzek77gWZ2Ljqy2MHejg
SwNP+r081xs4TaCukt7CDawEqj8wVTx8jhKivoKwXW75HDARcvTcZNjy9bxDcDPo/wxdF6Jc8gOI
S4/KQSeIei8Ff1foPYgvs1a0Pv58330cp+v8XMFSAFdzCFWLGDX4d8frlBO8pi8+amjN2rzIN+n4
/4Xidvq+/gv+hOV/ICeOhwDOaJjpJvWatTo74MjH1YYfL42pMEIst2j/bzUlYdkpxvf2wRS8Hjmt
CwZ8/LarXIxRUtxvCstymqXx80MGwqvwCw3ahUiiMuMgABlt48K9jr/KnV2jbM86Ij6cBCVUYcPO
YnjqVd8T0r9rREbesAEer5B0dYZKA463DhBAzqxS6txBRNDxdQBd3FPcA1UIeEoOiY+c5jzPGBfR
9TZQRo7puS0w5zv0zgbLCkzOC36iscd7DppkY3MfgSsmJ9i4g+ev9i+upA8z6e2tepAoJNx31QMR
6AXV48j0b5TkF6TQ/sEzBkcd3AXnvyr0A6ZfiirJbJYXHb7TB606EJK39Pvinw11tgDzjIe3RHWf
o21IpcKv0Vvl4hczWgKmqkiArZ0csw3prS7YNUsJY6lNFWdh7+03yABxnoHm8D3kdb5208q9PpWu
t/jFVM8V1x+Jb/g9TLyhj5zjEYmzJ8EbMpKqp6wIJVV/umIs08OGbbSeITi3pKLP2Rl66GEwYXuu
l/s4K8yUE6l8F58x1YrZ4wooHvq15db8BflT0eqi6Hy8npZDUXQrPe6CuZRf6JGidZYIU+WqyfGU
vK9mGP5stwWXXsUnqdH1AnGHug3qremJ0zYgdGX7gmfpfFm6aMUPMaugFjLYKnnf4sgVywYc7fYe
wTKXKWgYsA2waX/vA4udg4wCe9hgprb5+NvDPudpuEWXO9wz8paJZTFCP7G0VLWM6852dEf8HqQw
mRkmwv2e85RWkC6WoMg4nhpHvUs0yJEdMmyi3Y8Iz3SYE7h8RcdPdeFcfHZ0Hq044Tf/L8OM/y7M
N+1eVOEiOU6wFeMtJJIg7Nf3LQpntiYMbYjOWqVfrzj4XUWThO/rvlufdFYFBxeT4TzXk9KZyeod
FYmDIu1Xv7yZtuq/jU78xIebgflHopRlciYWSlJ5n2GbZQGDth6vx83U3FhgGURtKUlkcPGczC+a
Y+LTQgTrYwmc8IdSxWtzSW1zA67t1BHAc7w9RnMVkELfza7v7Ge80eO4TxFD03q0dOAyHJVxovRe
YvYvN4rV9qEVoa04YguxzROWc94DSclZF1hRjY3kKyqCNcO6enZF/8gpTBZxDkhF9ANiup4EjahX
JcLRDTYbwPYg01kJ7ukIk87fJrblraOsOnS0rQUhXm9+IsLlr8iZvV21mZXdXM2nLBbEbNynWzvj
Jwt8GqKVrnefTh1Ei7w2gLL6i/xotbw41qzeepjGv1iKkoheVQnmNqGKpLPkmOwgPXKx2ZSuqS+9
utmYOMKphBM7mEt5lLAakxYaQIeRRlhWnxxAJ4pIOC8ydrJ8Pwxcn8AOIFrzMnPse6LsniM6aK50
JkPy7yHO7/6+TmynARXwLUANcPUbx0LU1WRKHhwEKh+CzPlIsAser2SBJ1po7X2+3bJRsLfqac1z
IhLhu9X77eJPho4ulsFICd3e3tvFm0756vGGqQnye0JIHQrYctqg2EeFqoLe8Y7w+/xSXeZ7jsPA
mvET4YP1Ge/WnUXg+5LUmS7bxrAcFbIoGtfjWBQANXkiZhxS1LwzvC6HwER84u1mHSnY0yoS0xsM
XAxZlz3M4KYmYcj3C9ESrLsZnr4WDrx3mtPuBvQMRWzJMtcw1Ioeir4cO4mYIKjsn876oDe1W25V
pq1pOGSHxBFOedBWYPtnPbB5VV7EoLG6Jj0j21oko9w72eg9TmdH+dHZ4AAqX9ism120NgIdukmN
nbd94Q9KPA29dRdwo+nkbzh+iE49E7wsCTKY0NOqQsrTyHfLDtafef0Y4/8hbhxZ1km2DQzjGWz8
oSGcjnCpScNV19JUmXGYURD8ZO0lMyBKfS5jeqKMDn6l+OE5PY6Fm4v8prvDAFKNfJRo9AvBAsM1
STsMGhVF0ZO92bAAhs/mO6cpIAsOMiC3hwbKuMqTry8/eMFexrPjSaioBVIxYLkNsSbj9VKr8bWf
JxmNvyFfZWQ2KrnbDzb+wLDMZ4+LNI/7JA7caY/Zl/MNbJ6ypdIxVX02qfXvrhs62IxO87JYPc2P
IW8xp1rRjmw0giaEcevsqsbt8yp6vbX6fyW8WFuy8mYb6CjpQMoI8pRwCQ+4WqUhsplglUUHm042
UqiAsWM607xt9Lopso3QZkYYwJPZsWHJWOl6JaRFRzfaZ1kg0TfmFLrhe0XJdAAtCgzOyM9vuRCC
WYIkfSAt3LwytqltzpUKPgJGXsOiKwQzivAB23F91uXhZ2TGGuADj52w9LmUHwvwzY02qwzWWNu3
UyDDarW0UHfwTXpjyTdKvKItYRzAoATht15urEHVTzOwOSyz+UYu8UiUOm4895BsKRubi1dQ5aSl
+e2jxyKZgfUqiFy/P6WRD+8axlIsggTPLfB65pL8I+E8CDdxiR02EYtqF8sLQLV25VEbLxGBUJbJ
Frn+1sS2PATL9BepJku4OYD1hEml3/BpfSHR30fh/9rXX1L6rUXkYMYOJ3x9Xms+++zF4E9Cl3LI
pvV83aOlV6I9Lx+lk/HF/FG7EgcOooKnqgFsCCL/13MAqmle+BBC8kclcieExVZs8AZEMmxEE9SS
GU6U7y2zXqFEs+vu+Z6PwZy3Hr9p9YTuIlbnfP8Y0CGm8Qafkm2W3cSpKpZtB20nROhyNBw65x5k
cjgVec8UwgVk5oyw38nbJP8gV1R9/93cOgT8iXBu9ZLVMDz/oeNS6/0MfoREBV/9zDLR5Me15J+g
MH/SRI1NHwl1Bmrfhclu/h5z+tmW2NSnc9JNv7fApAYb87tLViA9Ff9fhXKaUpTiwmNts9Sng2IW
vPSdM0U+Qebu+RgKrH30nl9hC0n181HjF9veq7Zqi4O3KbwPuBbfK+nRJr1EcbMc9EwXiLlxgzHS
DRYHsGzGOTHsMRMyE7mtjHP4uUEvmHARj/P22JtpmRdkz2+3wbj3dQDZ22Z8riqohjwZngQysd+o
2QlIxuzqKgyxpt3s7hdTzZ+9bA/bgQQPiFe1yYLrjXeEMdkBvRwGXYXFRfyEF510hv15SK2GKjuw
Zc8e4YbSIN7XxyjMPDfaeiktg+YeN7DmwU4PAnaFD8Qotot5pZNEsy1892+/SGgYeCwnbuqwz4oD
g0ziI319ZaQtjRVxmt4vTO5ZQy5XNnjz4kCGzhKdem9uiOMkZ8O7OLXaDi7xNgkHHPs9Ou+L8l7M
HSvBGdXIgbdsUvUnwpgb2hUp803A74k/FTXtv8T50pUeNbK7FXXuOGTSnq4Mt1Q0z+RBajbPGTw5
C/GGKzaJujigNsUt8Y+Mrk0aUzewQGCyrwZ9J8plPngRSkmSpIpw4NP3rjU0NSsvPBv4zekrqsbi
R90xxvokwLtpiERPcbLiOIMkLKiOLIGS+qmvleHmaGctFE0oHEFqHCMXxL+ru73wG4qNQMSYfYq7
xwUKaRsUp52n1RrQl2C8KbmYVhnEc91A75OBBlRQlXZf72q1dQ3SWOhiQekAWMKbICM8EyH1//h9
sTH91rPAqORc6x6PS3aNBJGrBnP/ZII83v3yReV5BvGhY1zWiNFAbMGU6AdXbAI2DQOFlDqvhZ1X
4pjg1NkHh4JwZjXnTH9SIMXbNvNizsLT3+nuvLL+SNJh2o+Wz4K9dhjQP3abeaf7mRiqKwIFWyQy
3l2MlfSnKCzDtnp2RPqrACFPVPn2IBOSCDjYpSGxsxwHwuHoZQ/iaobO4r3V7eRLNSOyoF9DRj3l
7I2hCqA+1oJ9QNYE8MdJ1yyq3Btrb4JmWS4XH/Y+pM+FcsE0z2cjaFeVyIcKGxTZcfoSMRvMb2TS
7TseNW/EZqou5p/lKepgTzLgdzfdhpdOpOLNU8VLSOJdBQRmGzcc9k2CrszASYVW8Vc3hdrS+CWz
XdLy9BDTO/qMs1v33skPKdDg60OdyjCoVfAZ/37Ocwv13y98gRLHQQhSW1Te1VYVYfR9hkmPXChW
roUkF6yvvztc06Vh+PXVSHJWe0Rhrps17+OyDjv2shkpF9pP1d5/VzQzLS+EaPDiiSMJuUqKnFXh
DddHtmAe/nWWsAPnQYj2uO0xR+/EWz5RGXx66zz7Vt8/0SuAc4ZQ+eDyERkJExJUfMw8AJ7yufFK
oQ1bMLsHudsNETo5Y+64dAFlsHKlUoFKImUsUFuXsvNXzWAcuDCHNZrg+dCefVfCZCvppvgMCV4Y
QJHpPGkJ6pioDOIQKZLcSDUAHxF02/rNgoGaA13om6ib1GNg3M7d0gHJnnjFdhT85/GM7MxHeBUj
5+HyPAnasZv+N0//iLse0FVsmRYdtDVpRnfLhKB/tWs+E4CY9V/oVjWEJFBAcKWCsqYFVWopDLpb
oMdNSsVbKNbD6KR9OlrMtuZIZ3m+jO5mibCB8ubMDsKnQeobNmlf9HyzIvKCz7mi69Y+JZujCxFW
GoDKQh8Smip5Zb9NJIiwBTREgYzeWc7i+17kXrMEmheUrdEPv3PEJ8/Gw8l6Mf9d1B7UUzXoCssd
HFyToAVkn9njBM8aPQ77GEiYXNhcbJn3HQq+UZIYrjwXFRJTiJCWmoPbfD1qxYB9DKZuMvk+K7c3
Kst8mCPNcwrV6hW+6RjZBsEcYSt5sg26xQReotIU893qZ2lqhUYXCvGT2V9tY4i94vpmQ8FLPCbA
q8vfMvjhyHULk+2WhoLQ8HYd6hXZspoBOxSMgMA6BmFRGgSeK4C7Nz1KRSGvwJlzWSVPXvk9KF24
qNwTQSpjRjIrLmFGr/U6dvlBSFhd0heOkbnaOB7aGs1aBpWqU0AperzYvEl5BtjbWkKV2iIzCSIg
yIgxHl/SKu4CBouHB+nETU6AT05WWkJS1pzJ3d308LzhauzhE/TWI0xM/OBKmyfnwVwfjj3TEptw
YXiVaNVYwmt0GvtSt2m/v8oe/a7N8kslF7e7qMP1FthwYzNIrq8zCAsr2XU4/sSHdJhIko/DqmXG
KQZ1En8Ifu6falw35EP46isoesu2tcP2bu7rj5lEAlbqokyqD17ANxXPF6PBKI6hEsCBnKJFBV6Y
SrSt9DxxjGIUyY7N8eqOVOw74F550/99we3MXxbz0/ElwF6B+1nJGtDIepHAZtUCSM9B7k2IqsE8
+YoZAXzCTWacN6y/A93VroaBDK2UqIztEbUbO8QQ/7+b2jr1te5/jVw51GKb7lCb29uDxA2wzbN3
W4ZULn4ho7b5Rbva+5wR0sHQnjzXjpH4HzDnrq490BXcxBt2D0ln0FrVpOspE5vz8Vmx6O9Aeaf/
es7k43WbZzuleMZxQ3ZkJGlmhFOCj/QY6WR45BubztL9olTU2Dg6ME2k3CuPmt4KiNyZqS3zho2F
opFOrOxpoDZBlyA44GdQ7nnIL28co1ZiS8RwLiE94V7FoPYI53j+ZSabylolSuyB8lKemRmUuxof
ELdIALU32f6NshZkG9nJ+3yh6xHpohJyWGAA8gZ4vBp2Lg3UDzz8F+eC7Sxa/I2tlw+VZPCFs8Lf
mfrVncFBawA3Zht27YPSaCN7ndBOB5ipQoCJmfq2FgnHq6Wk3tPB2SUbPzXcjyPukJPFwWmKNIFV
7KEn/l4i6IFe+UnTsDxG6nHb76ewIra+3Zl9XI+oFdUFIwFOLMINAhCOjCYTDLWY7lDnzXJ54ULR
2jbgkUyr5NR57Wl+65dZog9sbZem3ZQO3iKGREq/SIEZXvouvFS+5F6ZaqTc/DADxdPt7/2/E+BR
5vqdl2MrNjYuDvfdmWUQCsymsZ+R40xJdrhLIKOFxJlijz3mHUYw4JRpEAJspAUv6BepDRYKotnV
MZ2dTnT4cMahFjeXrJw5uLNb/u3ofBw56kmo1TdAN2jynT/AGlSMiEMFc4uYvJ0QcVT4HRIy305v
a3/AubIdFwmEcfZ7qbo4tz/6uHLEH7tLpCv3r1uTz5CAd0XALcdD4+tiEf3JumPvwP+dtzLNME89
szX6ybfmnThHfrNBPUYot4D7zMjv+BzilLNifvM4TrVVsWzPs5nviIssmgJa6xNLgSfNQvNpWdid
BEZbnCdpDOptDbNgEjnGPICDn419s+TzqbtAPg0iT7RY/rEaofhWGiph/aWtZDuHJfUSXhP134Bb
Dvt6TOf18OWt359o+fFajSk5qpeBWOgkj5dR49euTVwXVB09FUEWMOX5KB8Q11a3HYdwfIbxj1KX
LI1+z97b8bY7XYZ4HclqXCoZzL0jFrsNSfWtdhAmIpNllfFjUmDhN91QPaCo1eYiS5G/fxF7abl0
l5nQxRuskO32GsF4yIKD6pNzYYFCsIWnzmXEbQXOfso4iFM9wp3JiHEa2NliOWiyQLcalngdVWLl
UiK9gogAKMv0pWvKiJzg4AqBf9rJL1BV/BJueQtP/c89VKBKj6n+ywoqZWBbl1uDtx41n6vVW8nQ
fQOqxuQJcOYswqmeE5HiOWnV33rz2MecQgHmfChX7vPY+tXiq4ifS8ZA0NVdDqU5ZPkK/fACLNVT
VsqoYP2OIeFZaJMkaIWI8N76zl4t/287a+RYLQ/UN0/MavpZzkTSjhEJFci570/5VDrsSUoxPl7I
K5ierL56S9FaYo2W7JV7UAdMDDd2p5lG/9zKj8Hyj76NH1NKxdyXWmT+QHgeUOvmiuQFMG6aazl7
DALjpS+amFDaIHiu3l7ddn5vjOo1p0SilVKnJgruI67ZxaeGUGADjMsGntAkN3wqJEVZdsGTtTL5
EUL/kyKrGQHTwxPEa6c1ufDwsFa+UfD9UwlbbXI9AzZX7getmElTswHsUmbwvpgdKoM+nLKWY1Ig
ozW3zODKiNtRdNNIFKg7OEWDL4ubgJMQm7VfHoZDMdDnWKXP8uhtVO1fLBnZFH9VyCxPY1Kjms6v
FZXgqdekparB70ktJV/jI9RTy1NUFTqZWpHJd/6cbJpV93gSuzMrMhiG3gs+9/vcXYxFs2wjF+YA
ivRT+RlrFeyhiLruBDIRKSJ/pJ6XB1YQC7tjIWDoAh4VgvDqpJfGcooOrjfjSxZRiJcSwkZClucq
6dgy7L519ArkxVyc5kZnOO2bNZg0KvVa2XEyCFfmBmDeTV7Qi1EiGIN0wZ+NmHeCSXQjKt2eparH
QW+BOSCVVKNjScshzuj87ISPsX5Gjfd+qFLpfqFY47lu+ePqZzcLmDc0PLQWY21ImbZXSiYhGxCC
ZrtD4KBuZxHpwG9MsjA7hYZcEjdufcfsxKGwCXHz+o9iPkn0xe9NXcDlMQkVkIMpsp5e8M7aGN3l
RvBBwwcl5JJBBwzGP9xMr5hiA9ugFBT5JDaZIN+G7WPeSIr4RpoQJ5UO/11kHlqaL0eOQrHdQ6ca
prVkOkQbRvOSayNvVfPU4lbTS8LACaic1opq21ZAt6pSfHiKRGgJItqkcFvLh90YdLna4TpLCwyK
rGsk+LF5CdgbrD0Y82CO7vGW2Pd4DvrRR8sWvPV9+VKhngsmb3Jzshn6hatGy4w7k08gKlRExVvG
nCdfvWR30xkf+2fIm9r9NnEcRZPdKqfI0C9c9iviz+s0xaMLJw1uX8qFyManr1gx0OLJqtAoK/Z8
G9u0hF8Kq+PWSgVTJ12sxsziKOxZ5QOA12CJ+LUO8R1PIwWDgh9U4tTTDLC1N26iETrtCdPlYbTp
173c0hDeFXQRJQChx1/7b3YEgmuLUE/Tb0Y6r/L046NOTAge7CVkNCbqHtqVqBBXmQP/1DOKaFVg
3Msztk3POVD9CefdTG4h1Blo7rlDoTg1QixhZyGms5RwTs1k92O4ZQhBTf9TJ/9hJRrDaNflALou
F1TqyACQxhwrOOrXB0M9maudAaJOlBGf83UMUQIiZ7ZXQ5DrtmE+StfGE8G0JRbHik2yDDvrP6cQ
YlNnA3HPArU22V/2Sm1SoMsjlp8WfcnMggjuG1+vxGev98T772lGhJ+1itV16ERitGBPkLNzrgDA
DwfSeFd0aATdDbqIYnS93/nq/587rLUnIAFnaHP4PWW9Xu1KXGygYkCAFlswTNWfWwSaPoOBi88/
SKd90Bz7g89OSrd4nHj4yAeoZdQFEFt+iHUkgVccJHaWPe62zMumWVJWBt1Sd1pfRFV34cxmSWNc
w2YhXVvV52umE8u4K1PjCQhCZrjICXL0P27KR5P4dBxRB/ozx6gGw9StRtEKVbrplJ4AVyhaX5nn
MhDJzy42if6ANsxsTordiYZ/LarI6A8MztHHU2dYDu9Pfnc1cudkimvnHGq7m2jtUxU0WmO7drL4
FR5EgiAXmDdNlY5Q/m83/KWwvHmfvCK48GT6Fj7LIWwtltaoPt27+Hug2PPqr0xgwWwqPiNhzteh
Yedv9XhRikKOW5EvoHrT3Ys4VKqK2KJzLa0Rys7VSR5pAJgSu48B4gU1u7warVKJcEyRDEHrVkJA
G92abc4tA2G35LfPqrQ1t7aET4J29sVOxmWsUEAw5OLxgdp+1sNLO60ni4yfudcBV3JHJ146ff8P
1i1N4O7zr/IdVyvIln34ZOanjbaDY2zgUTqEOVqK4F46I23xVABnuF1PfZlZvx1CcyZF2ZQZ6AP4
6dktoNKo7/tfR0umnbnx/A+p9JBa2L5TesuBTQLD7+F3Kc1/jDkMKHhK4t16md3Mh6O4jANwEMli
hbLg0S1IEHImbdFIO4ZLKnY7LW06M26+0YnAcxXqqXUXl/9+C9EZyaZUg4dE3ELbg2N3iVGPRsLz
UEaczhokFLJgiCOOkV8cSn4YzF3xQqZTamYHempYu1I+i96QMjPFbkYqAJJIjEoVDcrJHzMFwKd+
HSeauyIl35HyHEhk9PxjYsLCThgF1tZfvIqfNnz8sM/fZJIQhnmAXZwQj0GJJ+GotynJ7tHVcNLs
yj5Hpuq9veXPmUZjg0LIi2xdxABN0BrF58f09/T0xkEmyWja4Qv9lD6aD/0FDLsbfptsvIxVgx3P
o4VHnkNOA/n3UpwvDm+NPeCsrYHYH2zq66ghnUe2c49ZJ8JVkxo6Ati8rw82UKSKZsNyU/YwwtLm
1dO4jvm/WwgYa8Vk0BCItWgV9hwGlbSZGwnTlBnlYuJn2pxfAj/bmccTAzaSPGvKgkh6Litv5K3V
WNmngP5eGVTSLFBJTZoA2aiqmMB6v1EU65nRNS3JlrDD8nyhABsXh8RoarEM/1j/MrvAve3zzDqH
Qtf0ufQwk6beQU6VI+MN62OSElr3afc8dEUacdQ5SDkJoplPUmtfECfCqt6UNGyNaNr3P0snCzdc
Ulv20WviNQ+1v7yBxw1NcESen8VKO1ACTRUY3w4otO1hZfbQEq1iTAQE65c2c19BdWOQs3wwXdQM
XaO5Og4VNGAtdhx9+Xfz9QcR7GQYioK9qxsnvFiI2qmIbfj9e3IbdvdpgkT7zAFR07nPIimgfesH
3WA2scw8XyQPcHvryKuxOR6oglSfbtrCjdpCCZabElUd37mPzgptTuYHEbHHOAxPvvz7NYCo5PTW
ypAaVL9Il4HuutpVfk4H3x7MuGIZ/fmF78Bjr9sTZ85qSe0QvZNuzbYkZE6E3f+lkCcuaOWbfzFn
9Un6N168GuGeb7KSsqXGssR9LOrqzv7F1uPxl6r44e4ly6af0XNDFXXFmIylRJ8Cpv3asLiUPXLl
3YexpGxtvJa02FptrGdPndp+c3en3+pf8vvFzMWzEeWo41SxYKE2+U4yUnv6uoo1i7vOsjuCF31e
UpKRK7qe+Xnth9NFZy8JDKBmfrUIQAKkmQ6f81jaPzKghGr79geudtvUNgZlJthGYzJ1y5Bsidu4
lXsWBo6IL4c6lBk2UUJz4Uw4V2TeTXL1NyXyiJ14LGehYQvmTBz34Q77/XuDfTsurzcYW9YIn+BE
NegTCXQW4twBy0Ww7IDD+8Sk9cUoLYwiWNJYQs+TeX/hXte03NoLIrT0nt1VulfPVJeqi8RTjYee
rlXA2ZPCHkAgB1CaY6XxS7HiAyDyW7hkCPw8EQtd7ytqJrYKx/H5OKwvP3dyPcKeXh/qtWAeV1L7
qfPWVRvw5Onijtd1O5h8WMjPxUn2zJEyDtbUPCWbsHImngO6FQnPDU9DjNYeeVcm7ezlCq9xwKXW
b/qtIuiiOnGN7q/4W9TWPrgjnl2rVdshWDRZe/N2gtsbgVcyDMO0ysoI7E6XDYAqI9WCY8iDza/x
Sm4bFb2iYYlTDz4dnccoIVAF8mVs/1r5LEZWe07wo3w5ps/ntoVvmyGjLC+Vxkn1OQCP7hSGQmDm
FNfCgbUlJsYBRzYWBs0BfXjHFXrewQXgcp1LIYJFpD5ie+va6HFtxSwu1J1+Er7aooc7AtAu7NKi
HKrNOy+ZrQoiZ5/d1s9RLpED6pb9o7lvpGXFA2wZQCzRPlNke6/Derxr58wLhiBLb71WpKXU8fXw
UtTmMjbbSEsiwCAaLUfWmf9U9wZXsRqKL8LcF7JHCys0Wu/JeRhB8GOzEpvOej1Zghaluh4Wis8q
+JBAMFjqQSgDOa285sQaTmpPLmhPMYpB30C2H8C0Du7v7ZU4LAdkGgUih5obqKuBws3UQ0p415WZ
2NxhhG/TK90R8P8vjZuEvwxL+IA1BE+8Bagd2xMpqVYywvUEH4CCbvCT0UQDzZzv8wkIeKLh2Z0p
obhgpZmye8JHVK/z0orIdGvLI36+upi9MuWHnDj8r/mPOtQOtdltGUi7rOBkkHDawkFQzN1c/XnI
1Oq3kAuje3we8H6hzLyjGdxDfK3i2qFHidI6KfV2I2EXpYKQjZTc/+qUaoiS1UIqYOYaY6G1Akai
6RPbMU0iKbL4aN8dF61babAas6N8CUZ2GV+I4oN+iz9HB9eCUWPIeg9iif4htTX8NQur5Y8givuk
1cb+LNqDWk5XR9MDWXg6HkUAYXTuLnk4Oica6PfdCb3rJJL2U4Haw7zKkzzPDXF8scvX0yyYouMt
yu7TexWSX72oFO+PqVky6W75kBRrLgK2Jc6bkmplvriLfE1TUHvJQUE6QsGRaxU8fuvOUklQ+Hew
M3rmVZZ1t9rnTEaLqe0qb3qIbDTN+nTKnZLNtJUxAayCRIvkL+q3BfBVfBe4yshfmfpxDvKWvB65
XY6pdQ30KdT2ctScs0o/YY0nM8fpUIjXh6wdcYXF1uxsHWzacsDfIzGJMQ22UYbe0WQUnhEFFJxW
X8Wtl7NGuC/A70adYVSSjgc2CSnZX9zgfil5k2qNv3rYBdCvhQzMOE8Ai+Nl1mfhg6DE7bA73ZsJ
S3+P+FO7dQ2nAaD10OFSHC7y8glIwlV7RhTWQJmcNo2KoEhL41aHF1O+rGIQC4otCkRTWgz3WHGh
WCdlzZOWktKgQLFc/N/bsQ1NirQRHzCJLr5ixSEQtuNxY8i5elaUJtqOtHnFCDj0Fj8U6EJVrd1j
Z7aywQyG8U57yCTfRZOkB8Aj6BraixK87uC6v4Lybqqt6NkcwHX16UjFjTC1cxVNaLIYwH79jWLS
THdh6Bi+QtHjZ5kEZmcz+yyFI949k0DA17QBahwaGJTR1J2Go3Y2CB7iXZaQE6HLO/C0OKRzZ77i
ZGllY/SLH35Sqcquv6bn7cbwyUd8b5pRyvOg/wiRQ1mzcFYoxIH9S7GfTCnUWSaWb+vLjRCIaADE
cmGEn5BadDhFvJ66hSYc9h3Rc45UrQYU9iqIV5ctDdr/U4iW8RuTL7YKgP8l5YEqkD3B1xueJr1h
OI0z3xNlpqyuw8dnyklMpZywLKbCig3a907pwxcnsx6dazuMuaurqxWw7LY194L3gpftAXS8e91i
2Kmyyiy1iqV4yBsMkvqk/2qOqPFXM6MccTqvTak/xaD4wkVFK7hlauWCh+sMs9RJNYqpt6Rkv9nH
NQOpKsFiWs/NZ0HS55doN77VpcXQDmNizY4UzQ9j4Dls8uIy9/IqvR6T/zuRlL8b+hqAmJNOPN9a
0UIMgERzD4dzdgmwKjxV8k4MJ9z6JpCI6GEV9pAP9lEwbiWM2cDfgnPVQ3mp5dut9vVoi9FugfvP
PBM2teWpBo4Cf04zeAp/30aLWvalucyM035Csn8VG7H69zMZzhRjy+M50JS9Xx9e6frcCxR/G1Or
SctfgI/poobUw5uTgyYLSgq/r/HcytbwHzCJe9VqBJdqG/E7smgUagFciPDMHxfLOyKFipuMPUWL
3HqqQKAzB/HHB5uIjamJQac9tPvKVewIhJlJhWQY+XLGz2+21SWbXV01Nob58qe6oFK9JEe1Ixnc
4sefXKjJAWzW2n2PlJXEintrDhNu5fW9z6nTisjW+zQkgU5hMSB5IlywF9+MSwXLGwWKvsUNtL7U
QumQ/C9eQg2Qt5tJ0tflPAC+qYJURva3ffe4Y7z13CiI3DiEAuJDDEJCaJ6nAXFX+yG5KMho9hXL
pPVa5YAoQCTCJ8iUlqVvx8OU4699oQOjBx1YbIsWXlxEGY0zcO2f7GkDuh2TsxbDj3sayEH3RBjA
0WxlWOXQ451ChA+mQSC/MtUitxOZBl0mDKf3fy2Lmo85/tVPEWZ1G8iQoFZBwquMCw7w20VTI35z
b0gIcWrbhJ1cidct3rElYvHnZJdNshGzBHZusHNlBvlFHY64mkscw83yXOPz5uqmSvfNufqMyt9N
MSfo83g8xToUSsILJyJ9d7SNjaSZDT9gQKY5jNtVis4dECFJ6zqQw8Eb6H7GtK38LHbpY2Gs7fRG
CEiNWA44hO8197XLH/+2j2+mn3sXEpoYbIxWGWIyufq20IQ9qPUY8dQy4Gdo3O9KLtWEUe/qTm72
V8/GIRbcV4hKaD3egsTXNmSipwKI0j0UJEL84m+koWQyglKQF6GucfKsxcbqeWWLIqgx0AY9QSap
syxzQ64leQjpRONx01+IrIJBE9EydUy3iaiZP601J9WGuHXBxtodVFJ27R8/hDOQLRpFkcrfZCr/
ky9j8clhQvO1EDrqi1xeKt0o0mR1dbrKt2clRrVbhADutC7i3NWzXcSlVXO0kaKT+aY9dMDGhB4r
Pzpboe00AD8JMVH2ZkCKgBKepJRN/xtBhdopedGhb/SQJuLM8MJGBPbv6EU/PFT80HyRYwJxfvS4
N8+u4y1bdBM5sKLOm00oMIP3WUBVWuCd7VG1Qzoj/cI7zy1arINwepGyUTBnF5WoPYY8dlUZ701Q
U5zDmFkBed5rrFKfdtFOBuOzA+R4pcOkKdUeHPuYi/kaW6piEpK9JWkhvXBh1MUSkyG49Tv4KNCo
xyDpCQNydxzaS4UTnzv07mU5fC7X1H4EMqUbuETNz+LqIwFoB45IyvVIFreEzwytSmZkgq2YY6N9
zOjf4H2AjVWRd2nuH6C4ZXueOyYpotFaskqgvrXDj5XH0qcdojjRTbo0qZZGVABmYfI0XXSbDzm2
V33i+XvuqfJ1zw+JS3ymZA/JEkhoTL5F0f6CzpIOpSvq3uup5u7K5WBhR4pgq8pbYFtap1/w/lem
lhRKOO6kuOEG6Dgex5dcNKI5zGxc+yA3ErYlSTBSATNRMRqMcjklOpGHCn2po/xk4R1E/XaU2e7+
MZ/jlxKS8dl6YbKumREG2Wejv5zWvBW6HkjQtFyjGOj21mjLSOJsPyNocOTG3kzRIWsu8t2KMzKv
tRnCwidLphlq/XdIDji6S8ABK8s+gfEhkhE+4OVHrCg9vjdCnRWkOYGk5qE0BfcUP6Pvu7tHR2o2
6RJj0S0iRZqtfRpP9uuP9GXCVrb84dzbrj1JB/kHndpWOXNKi63XFWXQmHknpiAiu6eG/4VUyxKA
vKMq0xLCu6LM6R2zVO4R5pGMIIkbAHoYpeTgjQRSdOrXeGTo/DMaX2hsgNV4HuLKsC4R7UZvWbgg
k7/+UkZA6xNbRZ25SN6pTQD2djkaLu1DazUiJGQHmx62hiciyJTHwTBYiJNYZh8ZFqbzCkJ9Z3q/
C6PLEn8BCs9rh9M4TqJ9vKESuV5rFGpm4uGwfZX5DEYW+0acU6Nje7XWv/pTWF9qsBClgs4mWCKX
V69Clw+2c/Ve7MYKvQIz3yrhjMnw0Gk9t5r+kKW26pbsAgAVVkEZaoW2nBI96LcVwBjtmNNtsnio
YDR2em9z9Vo2pF/pboAIZyiOPLODaGqCNhiUsQT33A9T2/n1DQjXs3JJR1s44Kx7LWoEkWYGsXds
TSmVJHvpZFZ0y7WZ6vxm+cdMbJm820WB1btqcAiIWim/MvTHhBii1OjV/lmfuAXTDlbAvj8IpkVz
0EFmpq+Fz7WeYd9hQVMzM+uwmqmXlcjsFnPA1QTTVtMyL7e1OAP1O1QsHtkpAVnec+xfcPvRv1gu
JqjHHBWDOmDutoliEqdJ5xXDlBRN8lxQ5md18b5lkztpLQamoT/C97ZXCazqxOlq4c/JKVIimjfd
aGlfNatWDIncx9qV3DkNcvbaDM05HbfsRiX1puDtV0Z0LCdtKfhm2GZUgbVbVMbz+xxXhe4+qoLC
VzVp+fGBeJOaZUdEOaSWvl7+VxrYJTLhqB6U1tmkJrAQvcH1mt3dys1MaEdY95XPlDQTAF2sc3M8
pbwCLtPhGtEmyUmGflWCC8KKEkiMXXjCDazI8nX2TprEBGum8fE0L/6u/xUX0N5mDGHMpeI0BTQq
/605dQ/Wa+Z8ZEWR22ONiZ2wD6wtKybNF7Yc++B21vyXJVaiGlhBGcCfPYQHij768ijgaatPttIF
IHxLKdqy/biraG6y4ljQ7vHeA7knRL/eTFSaDY8TFaI8yKtKcLcpCPBEie7eg08PQxXmeSf4h4U3
MVikEtVHg0UmhjnvExn8BZut4FbhPmpfN1pFXdrsYzDmQhJs6VflREbFvfIWLfLmJLMiX59uQ12b
5D7MQakbtENPFFpaoleqnLIvWfQCg8EZdth4XxzonxFUNCU0rAGh9IR798IMkBmjWKsesfn8soVD
JTau7twsxQmrRrRizBvR0e8YWBp7brKr8SqyNMXXu4wzagkEQaJar/cksav2SyHvCvwSz0LnxzAF
B0SdiJhAqOBisG9hp5NPcTVHrD7MwxEcV7+59n75uRpl/tNEyDCLbW3otKYJ1mTogCNyoZoUfqVb
D2jLmGmrAaSqufJTrcPMoRf/0iWZpOm4KO/I5FqJWLCZXe1ZZXIz2zog2SLCFXSJfqqtqsVaIPB/
PXXYFWAPLZ/LpVP7UhEtv6w5up44PGmdmpKOftVK6SmwoBeLavaKVYdV584tLspthoInhu02+GNy
62cenTXyijW3YXeYT2PiPun51nVD5WORZj18KX/OTTTdsc9uNUZXbYe1u4Xd+ZLHoAK//wGMUYRl
BTB7vQctwHQQNrkZmUdggO//TVf07z7GrKHDauo7aSdv5R6cB93LR43pWIrOL7dL+HP9NX7CXkRA
piVnyCQU0/Sl6KuEbAM78R7j2eGQ8iD9ZaEdIwJWyUDxzbieZKGkznac1cDyPiQ4w3ADexHhu+1e
Hj8uCNDT5DWpc8FNXRMG40UWbsbA6iK2y1Abt1WbtZLqmH+DSzFPYEIJu5cxctLbKliLaBKPir0s
QJLMbRwFZW/wBOjLdVLlWlgTGOHcpLkeinrP7MHMsDh80PSptoRQLGASk8Do1lFkcnjA/jaUDHAF
FT7ZmuGDesBzMEzfGv6AN8fFFrtSGF0GZCd5Brp3qYWdUkcMiHZEA4JonKvGvvXBxsdB8rCRPNeO
YFtVR69essPW6jeAvAvQskxaJ2inhtO8CS5dNGf250MrfI6qU6xf2Fn9uAk4V1lm6iVN8Wy1QCm7
giKrlyElyBXbIAdVr1SLcTKRJNdcBTzUnUBKymcQfyz4OfjJIS9jAG83zv3NlXEIAsJENfnpqQCo
UTuMtFQovYS/aMFz+eT3CDzU6wce/VChvYAzqDcU19CKQzL7StREiLj3zqL1B96jcfJZhvoqHrcF
tJimI78OJEOuMzdL3vpGCQjJpWdkYmzMFdI+bt9ozqgi85njOpSBmKJtp+1+XWmCcKWiebDzPss6
U1NEvmFiCQ+O7TZifABvM0hBfktNhAhEFkUE8yetZEa2DeDWaNojSvhQU5qJTz3ULBdejB2zLS/M
cvVyLQfJrxvg7DsVT0929uvaP8uhLdE2jmgtgLeHZg6ZV0dxVZlL61vkvDnrvKGkiDE4qmEVp4M5
cDjw7R9VaRdXHaUF77RiNcTPeZgHqiB10cPmUXpW1Ls+UY8oqqu0YFxJF5vTmli5D6umfguM5awS
lQJdRbq/ijmAKSRl+vxbxDrob+W910FkXAZ62tbTEJe9OCDEjVX6i+jt/jsP3zLhBROOKO7V5O2V
Oxg3PvPfsQK7ZMcjX3gl9Y/r8RG/RTCK+w3ugNhlPCAAZn8g+Q+0Y89WLnyWBHwj6BMrDg8Xaf8J
q0wTgiuVNyRyV3nqfn4Zp9KExelStwJ1LGjHvOx5m3eqDjOAAwdc7Bh4M2FByJOWcOmK32hPKZ5W
nKOUyiK8vaxGzXMyZQr+HbYDhAi34Z70tWokn9OaubzCQ/iW+mLlknv37qfyKhz8gmJIWhpXj6eP
asK2P0gz/Wq2zUJeYoKTOJ/IKxxS973iP45kKuhwEuojO9jK0cKSMVswGMKEC/7XR+3RXq5LgLxt
+Zkg65BVaSKppMg7nD5cLeQFOJ3nMREPFKcXFv4bU7bAyOnLYDAnb85E3TEBQvn53TMdcMrJTRBk
7TgxGP6GtpJgpw3o3nLHHf0Y6h9WH1ZQA1HCWBD2268p6SIxAuV791fGL+UUl9vuNWMOpMbEEXNE
KVOSjnoX6DOy8v7ZTlEQXc/MeaF8VH8rIM6YJj5gsfTvIrWF4HRlWt7bCuYLqnfdXvNsTTXMEbkN
HPBMU2OgugErgRV6hxOa48f0qRMwxlto0lxsFU4D4QneGgP5OphgJN0s9ctFmpTpJtfpVjRy97oW
BSWaDf75uOa4eRfMX7GWYyjVxxg3h/dm7CB69/Y/KgydQMJfly78PXMPItAq8MKN7cfSQK0VY//k
YltJ7Iuz3hQTiJ7pTnEpX9iZRGF3sXK8+FkLHN/Zjj5FWhDCVOH5EUDjX9zFlkdMykrG6h4ejS2x
m2dybW88CsRHHGjJW+NcUXMPonWm+S7UF/yXD7dcHdDfvZJHRnIHo7P18p0aIow7tpbc0UqSXTCk
zaLoQtcpGVcUVSVFD0uFaujUlsQlv7IAVUGFmq/XDUgR+orJLcXM3KO9kV8ZjhGv4VVMj9c0WNmY
hiMJYv+93pspoKab8Rf8w+9N05ZvObqJCW3uIlqLcUMh/V6EiiXHdsHPEJwchBS1LVsZpccOdj+m
K3R7HTawUbsJsCWRTAJsrFyEkCNtcEP5BhmxY249nxsAjxPgbsdlGE/8lO1I6IluQ3oRm5N+HJVd
6YboDghDqZZzW5OQ1Ab3uEy/6rZO6cg2j6H9G/pYcJOYw5C+9Iu+3uNVs7JmaMVU2GANZ9cJADwa
l8F0qaDxHMCHSEEsZJSkXDpkHngWPVUyVQthjoAOB/Cj5EeITTghCLb+BjHW/mCSLTqFhii8f1Oj
AisjcFtvweOR1x75MsB0DfvoDybPX1x6knvdeN+BCLi52XaTua7tRC24CtnNxqbnax1GpsgwlI/x
NVkAowzGoA9V+bhS7Q3j0UWgB5Kum8iM/jTItgxuW59maSzky6duaZ9J4Mb0GyEeJzMnxGO/MhrY
jims/YskDeG3zQKe2XjpdxWaPwRShejJSaQM5FMGTVAKGL42OB9SkAGtcknxr6/mW1AJxLqCt8PO
9pceHcfrCJfVvbtit3wPo1G/HhQpek5AazjJJbjhOJ0akwOUmWH+yelOOMOKaWbrvDanMMTr+mbK
a4SKvtuZ24w5wWtOW7lIZH1+wt80vfcJ5Yr0x99IQzy/SD50JW3YXY41Xcfk6ZcvhcuZqqvEwWxK
Q3kQ3qYhY0aNOwl0josaE5llPA5otZ9b6zk4PbAviIj7th+7NrtS1Sr2SLCeE1h53WNUTrE34A02
eLvcPK8HFiwu/+hGj1p1w8VOVg7gfmkHunc+8226KtznkRyGbq5x5iR50bB+ka/nEdUBKNbcnbm0
3+uAgjZaMPisH79Nk/A3bVsnTiU7C5FfRGoGR+5BN11uM1jVtcfpURPkDIj6W1bzA8Lcq3NO2rJy
wNrxiQy2mA2Rs9aJ7KJr4in1zL2tulSWWr9P3Z2IjPJOPOSQ3/U+1QWhZtBywfVlq1cwFXTYABHR
FyTHpM/7aggpZk6e6zBnd9WrqHauJ6y1kn61NTmvbEUqvyY+L+TAiqMr7YzyU24Bc3pGUwq0BIN4
gky6PwV2W9OS9bTfCAqGkEfc5t26ew0Wqlwt3dpec7u4rb0sAikBHzNKtOoNVicspc/xzs3TkTdZ
v2PW28kHykOmKmuwbMrj/gNBtPVpXNjMFHc1+r4ENH5MzjtgZ8Z+ixsE0fRkGfpkQ8DTpNT7RAeh
By8zDtY43XchcGasyPa/l5bF2dChhpolQd036Bzb5pPF84wmloMzy360xmGdTlTXvxXfF5mZTTvx
7tXoexZxFgBPeHK53I4uKOphyYoOnqTrSAxeskGgrqWbhnrLGWLqIu6NQNU2wfwR9h/chYuGQHmB
09q7j/fbwai4yUEH2PDcrel0ffi1lSjC17WVl/Rgd+3ru7Y5IKo/fQRDC3eW8Wsh7j4HfFUNkS8u
vQlkFljjx9ctTgVna9L98CT+QGm+kyHz8Thtv3tzNJ/hNQmzh2HwWOh/h+TqrxD0hehhu0jcN2Qj
lYghVjnEvVLALljgWIIfN73qmZkfSugLpvhAwCHAUNc6CCI/OgKcVdlJs48ppAqaXhZUmtSlW+A9
tURwdxMi2Aqxt5clb2id5H+fgLEA/Vz+fPd7nJObCJu4EAa8UthxLMrOGGvexwq8sFlv5adffkOs
EwXarFKwPXE+WwCyTdlUvb8TZ5lltpP1YXE5a2S36eLKEy9xtfr3NHZazz2MXYf+BcOnRG1IHjGu
bFiwcBvJ0557vdHZwvloP0r7/J9ZUpIK/YXw+ouRRpuE46V6H9soUdND7oja1WfZkC4oU1964OKB
5N1jIjJYS+mja5ZMH+LeURO2//T1pK5NSbGc3l34JlkbgW7Y4Dde7A4eTEUXn8MC3UcDG2CDzNL2
BygTZ1O3qgqOg4R8cBFHcrZfsgSUZw/gWaonzS5+b+PRoa5g/CwCmYjkB13DzRmcFhDmxMD4cxck
x9Y7/QOGidB824jY9gq4OkK7LPuKI4Afkkjyjamc1VbQVmHeHOIHmexWTadmKNYSfYH2ldzWiQe9
Cx72kEJITKQq85SymqvsvBLz5Aq//O1wizTJChu4THm2+kzQhAwiZC9Q8VYbO1ZNq/FJ1JoRe764
Xu7KrjHb4j3AXYelOBs3Zm4ciCY4h5SfnmjikNvwap6bfYD6GdntRSYEyzX8f4GWAhEGhdh5rCkE
nG1bo0xk1AJSakM4pm3Usbg+wGwIsrz6FOEw4UxoXHkNKQIpoD83OQVkFd2KmiTIJBpzftYVul0Z
HKU9yZj72+x6NLNT08YMC2piIOlC++FlFZN97/Gj+erGMifqp15vOcpJeepzUzHLMKtVZMQ/QMR1
ftBO945/pBh39wwx1UqOAfUs20dRqmZXCzzO6GhFPXrUzcQLBSrfJj4jWasequJmaZ890jd3PWFL
u3ipPzQUIOH68IblHBJTAF9GZ4n+MAfLsd0JmF6QgO08wl8ci1WGHjU+kLSMcihGFhMYaRqpx2/M
L4Jk3oMcpm8LO/mgLfW2Em/sgeS/G+RwHTfmPYwdxOXo6I5AHxRKq1zdeDEgKjiNfVSIo8et+YND
jbcX64je4JgaJE4i24Lun/Q8oeHQqPitHAjhiy3drUH+V1ZdNG34CfNFA0ww/zhaNXzRS/43mJPw
XcO2UAdg72h1k+czCBEIJ0KBzr7wN9jaoIRgbQ9UmDNB+fG+uczCqaxXB9iuVS6YCRmeh8eyCYLg
EMBWbwmoofKaBuxDFwUr50SpVHLfITCIfaOY4C8XR5nZzHdv2lzxXbCkyD1CQxT5lC7tPTC7zFcX
yTDTE8VUsU4qsJ7bve6SwRI/zueV++5cHoUkak4boRIyzw+J0j8WQYbdmUJK4CEkfJB0IMMPCfwt
kYMYofnIjvKaa0CQRv19OYdvHZB10gXJ9CmeKGl8hjvQoVJWH5w5d08O/InydUvNS5vzEWoIO2Rk
9/Oxn7Ot1J/5NSxoGkRgaRWB1cKi6/Hsfif2PGzKcySdiZmft0TQbktzOrDzGqpUg1WEU5AvBXJV
5sAFb56XH7QSKgyDSqFlgxOr3MmARwv1tASZj0h1n/L/QdqppZz0yXN/oBHAKBtNYuH6ou4OfWwr
YoWnO82hE4ksCKG43XSwtPdubhDbK+YvTpadlnu5v8kEm/iDujtZvdlWM7NsycjE7CbkI3piSjkp
sR2TU/k2wgOsGSLDdfEzwlW1F//mJU/w5ot5wBKQNq6rylWJYorQBgMLQiEEInENE2IPuXnh0Yab
8q0vrRoH6U9wU/XCCq04RaafmzsW8EXb4cfiOyGZ5X6J6RrG7cjEbrzmCV2hYl4aJPwjXN60ms7y
2qb5qLkJdwEvrc0kDE6tnUhr9I/6mFCAnHow8GDK4RE2EiZUFKhrll0TH68a1ErdpdaXUV3pLcUS
tuY4Lh+eOkGu6X4ZdtI41yCNRjNcxrvqjvjBo9W9tY5pCfFSY5w/VQw7PrOXW5MLeAKB+tJ0k3VW
zfzaEkmNvPtvjfyJbuTMpq1L1iEEWwHWLgzI4wfFw9fC821pO3/AMxXFFx3eBjrZs9m6mMyaArHe
mjgWibCUAyLt1N2KmppeWcA0y+4WUGsGA71h09UAnHSJ1YHG6C6P1Yzwe5p2inzSGp1UiycP1YNo
ZLWgEUAOhxOy5oZR6q73/X9H0/HxoEn/V2STD/bk8ESWEn5wfXh0Kj0gIv7HrQnau26wk6BvdtFW
VunYIiD10Hh/6DELd7N6oJ/eN3/39S5uTURfU+GKjr9t7H94kpzEME8KZAzxMenFmDov0cU2FIAt
4jKwqCQ5vfqYeuqH5by1Jh1R29DfxJQU6JCKAUhkwXhsuM1Xpv/vKdGvM7Cy2MmW8HzUVXLCdo+B
zC5BdsoOiclrfZvNXCE9Wre5nbuzxwmx3QOW7ZnU9LmACemW6N0rJNsQH4ePP4mwS38NL8IXXHpN
xySP18Sc8fjcombhr4/6nGVUVTdqdG+5qpjl4qjhlFRFDuAG8xfTD7KFnjs1Qq195oAjkMXkyeYW
tMx/KSL/bqD+20KUi8YzUzou/2BWSaXuGzDGVUxsgmSKVsRqN1ojwSjpRnApHwelJvSqCf3wMbpT
wo9gOYuuNAHjI2DIEhxvmgz5/7sRKinAQoTUXr87FtITIteeWRzzinjEC/PJmzuytYz84LSfQNlt
tqqIlxnjFmC+L6oyhcb6w9IF3f+u+ke7e4VDWykhOt3mIs1B9j10DY1cwfXnD7hj1KegpnrX4hGy
U0hBwInDXmc5lRK52lP8LkVlz+K7mvI0TIYlxsZ/S7TocdehjH7GSVYjuNnU2jzBHoUUovU0lA8v
oHKyFce1hCwuLyu8+dh2O/oEyCNwssU/qUBslkJ2WH0C+EFV1V1eIRWomRe/Z9TCQKz8fOu+Tb+Q
GpnqPOkGor+Tm2tZUjMIRpqfe5OV469A2BUCIq/YVkQwm5WQeM+Trlv8hANy/Ei1IBDIYq3j7kQh
0X1jV7hJI1XUuBZomM4OAiVTCRx73BiaRdhFBpDGHenemnXuWer3e2s3EzIyZ9JOoiKiviBkzJPs
bEDunI3Ys7G4big65gTVYqM1i6AGGPdHrPpIoTI6Od6txzmyf+1fkz3CbO4qEn4+o3AdAj8rnuP9
gPsXaq44wsOmjn82rsO8J3tj9yBBb3hT8weRO8QDrSY25hSnlMRvV4/46f0Roobf4pYES2oJS2sE
l3Ojx+ja45sW3YVcVHPNZ4W7OW8XZYyBm5P31P9ffwxb160va7aYmiJEaNAL8Q6gK/1aXi9PN/3j
N7d42gF/sWO4H4woJsPhyHGra5+xeA0mO0xrZUP3ikGdJlgwA6sXGayFwY59sMZdX5ys24puuGYM
ntNFiTw3h7M/ytf34N5LceKylQ9Gdko7yc86M9giMc5f9NueqnfqaYkop0D7MChIsPAdNGUNpS+M
thUzLGhOAttUiLaN3Y457XDCfTtwan7RnNvt1dciazAO2H29f5Ams5xzhWzZZ81NiNqYCfkQQQ7i
Q229CfopfkeC8rbAkaae9zC0vyAixf1AwR7SnUBhiIHTBkyPMIaHBCGgyVkRD2QbWhep7BBR0z5j
NkjVETbhkfKBDTod/51Z64IO7YUNoSIoIxV3X6I2+QtlvgpICQi6n+hOLHTy0EMyr+9RfuQmAowJ
5f0vdz7HJqhbu6ET4/uGVAs/ZhyHfARavEFzPbL9hnwAIWPRVjj6hQttwOUwEJInXR/PbYN5mJFX
8fpiQh9YsPBjH2O/c9TJ1DhtHF8FkpEjsztwqXNudSSvQZ90Cg3OMi5rmHlVS/njz/B/nMD+sWg2
cVbd+2GR35Rd07ElLRrFeOvFsMpURJk3FkjvREkqsVmFWDph4Zzf/6xVVlaBWv3rOWLWvESBMtdZ
1YgzNR5S/zacT2U6hq+g13AYwYA3JrMWACfRNZ7PgfqAsW2eS9M0l2uEBJ5fsD38FVif2U7NHgKq
5D/pcHqMC+raTJjN0p/DtLTlVQP/n6nHu9QBRp4TU3ts+trbtum7zrLNKzd12Y7ivZt8sfvN/Jq8
tvv4izXGU+O/q4+YVyQJtKbQpOICvNVe6CyqM4+QkeSP64MvMua7cQuJHR1l8Toy2xabPfLudPRK
nO7vP3g+wFf4tP5p3IODy5g9E4XJ9cmwjl3ybJhz+wn8thvU8m/b0DdcgWKEUkbgxXN7V0RJGUux
XWFLRy7Zlol72UviCx0A7EOxN+D48wdadVCio1TbrIi8EIuPOsWUvf5JY80A628SmWqFh5MdCs6r
yz3ayneGta4eNmIGVXvlyFdgFK2EZRgvmaRXkoj05pryfgqT+Qrh6CxCBvzAa/2UnCq6H/x2OKl7
dGdUwNPVmjJ+Pa0aapuhXAWVni+oZ6BerZZ+Ab8p59Pnykiq+nbd1FNQumYWw8gR+5/tKODmvGlM
dLV1IXhBl3AozmKiCcqHCRWZ58mTyEr65oixpgxPxnVRnXY4iSEJanJ1reaXOcerke5ppBM1rRrI
AaYE15fJSTyuzdEvH5mBYrHGDUIKsf/MF+n9eHDI4ugIzPzQcGEAIuIozLv3t50uJOwsweqnTHMg
XJsJNmrHzEmQwutWy/gjg9aia5n9rCWem1fQtdpsR6UYIr2WLcyHMbjVVV0zS2e9iEEyNzeCHFTs
gixqaP132LF7Wh+xm/ELoK8D5vyGisKOcttrnbfa2uZ5TRFe8/f2t6bQMZvC7yTUK7sOT/RzFAy1
fIR9/01rUvHVvzu4PtU+a5GlJRA3zAL8e0NMPU6h2lb47hQk0Xdrl28/p5zy+xNYQM18QrX47+at
rFABK/ErA4IWOJQymih0MLiaSWJpxnVMaawNTEcofoGul/ufH1vbDs1iKykrcX3YP4s0BO3lUEhc
3yBGhpLp4l53R56FR4+z0UbTQvDnnhan4t3ZX8yCjdPhYk4xAFeHhLGXOpBNxeVxJI/kIWMheMMn
2FSDdJ0gjgMS4iQ7YrDDrtS2OCC1eSpEm2kRmlgeL38ij7wa+BKu0Yw8BCZ1m3BgXxo6AHNhxA+5
WveNPSYd/cPiYQlLy5hPqDVbpUnkpW4RmfNK1Qd6HL5DupNbat+M06+jC6/zJ31Rr4Mv8DC40i1u
bn7Q8QUMHQz8RD5ANwXlAFUfJ1S+tv0G4BbIWtIGNSUSwQtAX2/+qA9vSSzxGqzQitq/vjOA9Tcw
ujO3REg9mugxASaXoyyYbNIdn8O3ygD2CZzXFTpDjnQc4LEqcmCNIMH0mYYPVwo3uIzFBLxV5tQx
xDT0nOkBfXzoVc9n/PIMqjvar+It2fHR8JywHPOApoCvXJCPJYrz8FRe/TUIa2WYoRXOAfSue6hd
ixo9MruhCfITGAjRftTGisUQ6J7Hvv9rDYEenRAABsBb9MAJn9Rw93mFYKggcZOUCX1e2nqvpr7i
euAIpHTbJuxG/FVBXny84Jslh8Zu2J0c6HelG9OcqaMRf+KEhjA8phd1vrULW63k6LiYU4O9E2pr
CrQuVIDdwQFVG5l/b0N/N60e5FoG72iCH4u9Abv/dz1g1XqloINN+cO/CbABlnubLdILLAYAGq3W
KDlLXMktcT6yWKIloPnrGywJnGb+KxRb45XU2xHn/aivIO8oUJ8JH5XM/duOZNsuLC1Fyj3MTN3H
5UQv+FBdE0FWS1yjSN7ugZRWAkX9ysNZU8R1MhMizpnlcpJHLWh0ZBxqKhOobx4R7JjLHIMJv4LX
mqVNuDrI283R4ANrF0Mg8BvqoDMbK3zAs3KLxSEtGTrQ+hQmeozyNR1xQjL7w2jcU7DqU+517iuz
h5+E373VnJgNDluKzsNHX8BXTmtz/ucujNjNSwHz5XTs76R6zMgCL+C3Af6ds5jqbmfee5ZRyHIv
5HrFqeCCmTuoGeh4qDkbCqlkUvlvT0xETmWxGzXsFL+BNXRgUMZX8FQ5CEv/FmCMDPJRL+/Tnvq9
f11PiUaFuWTktdZ7Bcv6/2aM77uKnHXrkKfiaDzj2axtlq4jpAdgG/InfcwUEZ3LdWwaiUW1UDNP
SrD9LjHryivk07Bg0Rqmq7J/6I7lAxgS1bFmLmSHGVZsWFqrIAYO85A1I4r3/KtkZvlgfg2HZM28
GiRyQTeNs/UBKkYLrZjlAYoUjdap/2JAIfPQ1jf5x4Zz2TstjtqSAD9hPq5padV+JPnOaf03eR3M
yuwt6KYB2+qgv2gmuP7FQ7Yuk1KIIZRMz1G1Bnes3Pwi+93AnYHvFARF2nQxxbBLySZQDaewrD9u
5UCOiKexpd+1C1tDseYZktxvxBvzok3qNaGp2cBfU2z3vGfbhL0AiGcqF+YRHxqdLKFyDDBmXn8R
Z+zXUPlLn84qs9GeVlfwrhCoEMhb99bSr3HtdxYhFA/xEUvPd0yBqcoLaMxlD2aPNOyZynwmp+mr
6dm7ae2sx5ze6SGr5Z3FeB+HIXkHHfEJdonBU2prpyo8fkkCKieWq5vdNcBSrJJ/Q4lsJPP2fB9e
PQDQN0U+rLtOgFO0I9SPu8fIRhoWwb5rT3bcegkby5yw+7nxuZhnYavdmKXsUlLTePoiYlxpGcaf
RxuasjzHWFel0FDV/HJgg/qdhkVIIFw/FL292WYnAPx9Z5lWXabZ/Wd4/3cGcf34ZH1W3gnsnHwS
M5zlUwWuDKyzxe8VRSf8l8ovOwZWXFK43le1Pr/VJfmAgxo1t78053mHjQUHX9U6htGyGmzCuFXW
pbzYEt39HECoMmxh+A6iG7Q+bydSHdQyv32zQFbE8IWMkZ6yR2XeRn753Q7HcmHEs1IZ4TpzL3vv
QuFYAyaah2yxRrKeevVcxPhEa9yHDSYq8cMevB5wilWe0BIFwR/ol8Gwqke7g3RBf7UYwzfN3zsq
ceSy9ZYi5xvkmD1eM8yBs6NU+SlOnWnaqaRcpckYpTe6ZzvpfSlZGJqdcRhzK5SrYcKX5GIpSnfe
KUK1Xk6jg8Lf/RlrybjOztzlQQZ/LwwusnXXw756ukM1nyxFJTqDtcbL9AMZr/o5EEpTLF5vv/yW
OSdl5r0ztypBORxS43RQV7EDObDOdirNN34xQL6O7JlREdMsh2aPHdnDUV4awt6+DUzpzdPqUKo/
dqp14lP6aJO0nAGQuROoSyxmnX5OVMjBPJUQJZSWYumzE2KThZWTZy640bO9RcMUdT06weksjB1Q
59W+H/dqiAdUepdCsK1aBwrxU5SqWsxf7fhx6RCw1lMZcQYfZ6eWrjrVBTudUd30xxi8GXYcx4SC
z1tnqDoWy2wbqrsNupAexNTxO6GJSZEwmlxyf8HZff0aK2EYhHYP9pjV0Eucq0NP512aGJSExeAU
Wq+YX8O1gnGcQEN4e1rwk+JQFKeaQMWdQe126I6y8Jxs+Ikf1zBZGeLHOL6CrCldCuZlXLf52lWM
ltGml+QMznjTwWi6nLfSWdyYMW8DbTOhEfs66bUDmAQrQB9JGbuZ5tQ88j6uQBuiFHzHE1J2D9G7
7xI2DsT9dyaVMT8qjvh+k83e/d3FXYqfyAiRqxxB8ub+2xPOmJ5UrsVEYoi0luKjptvX47kA7LbR
EMnxyDyVy7YHRDRsvNVLZt7PmcYG7Nifxr261nDelc1xeAc3YOyiHaFjTphBIR1B5B03uZeo01pM
9ktqTd9lJdYdxjheowA9Eqz4ML6QUqdjrI7cAYFRw7v3EXeMV90E2I+C9+rpk0qnWEQ4YYZQvq65
QB+Z8MoMw+mJani4Qw7rj9pNb6YkokmjpmZmXc03olFL/L9oym7b3NlSJ7o0HYPiXxZAyOrKB0fN
E/jMvklp51mLo39GQYaxK+k2HqFK0dDUKV3AVu9ycHUta3FdHlYXh4HEEhlP+YAy5lFygC6naWgb
vy+UBYj0Dq2UPEP147LpiQwWKdmVJRfbTOs+9n0qIJGqiF5DLHPU+Bw8pHBhurF2UMyVK4VsH0MB
qnkIPGd/gq1zJY6B/lDcjxPEkwsIregjEKQ0JTjzu0eBV1c60Zank8s1c0q2mO19mVLD7drwaSEw
D07vqdTCeJZLpI9NzmZ4xKIQb1MZ9FdN4DIDeX7OWYisSwPkhWqreWs4sBnBGNZ1V0oFNS144DSN
/RzxUfAFfuRQNaBw3qq2p3nUYqGGMZwnusVoh2HI4alxiOa1L0vK2tisVvn5oukTCCdsqskIB8Rt
wsGSqYRGTs5cgLT1l1FxY92kW5bS/uv5Rw7QBB8cZ3F8g/glQ8Upi+UT5pIZwF1RSl0IMfNWwo31
sGP4bMtkkd9dS71vkOIFjAldR/ac+2QHEaNEHudbEMKCIKSUSSHCsuzDSrusBQMxf+d7qbUOG7sl
KfzoAufE6OMz5Kz4r6Ed0aIQXcsydCvwwzeighAUBlD0URAcEwwtGYZxQiEZVUGpgFa3oXHTRBWk
7ijTeh/FxPq2Uy7uuzZx5btM3MPwsEwc93ehySzcu7Uc9qauFspP3oU+nznZ5opv2It5LVBIIyWa
jKA+u7thLYEldBBIVARLB4yidYiNaOKnMVLsStYOS46v80IwLcCWGm5qZsQtbSneFXShsEyhOJcY
zS2xNKUzQac/I8EallG6WG/1KpWLdt87fYTTnkLgBWiXE15mz/w5vbnvI8iOFP+tB8Q9A4h0BmCm
wOiIqNLRZOuwCh3FUgYH/bl0ryVBH+BgUz+XrXCbB7mugZDUfn01lQUPkHynBFf1rkTVwEJdQtMK
t94Jbzq+rDJUT0Fp+O4CLur3YZItbDnuRgp/DcfWUTUzQ/HBZZj33nJoXyhlvoasvX4DPuG6+HWU
1ovmmoCCaGLK5ES70Jaca+20Y9eNTD6ifm3H6PFw/SmuzCrsqgpNTga/MDAXsacb5B0wxmDrR+Jl
NqcDyvdXUmKGVzRchssT0yKv5zlSsbOv8nq9VAR86vqSwqJMLKJ0wKLAyAH+6O3Fbm24kkkho/kx
r1YIiG67nwK/wnBDBHIgvZTmcv6S53l9wEU+KGd9eBoS98czS9sm+ahOr3loGfkFobKKtJxPfRJu
OmnHpyviGqvgQ0X9AxW4yU4b51V2ozB3kkqsgq8uAr23GOu/ofIfJH4G/sjq3a7zGmnIZ23OBmLv
1QHGFXtV11yFf+/Os2dThi0kNELM63I49dHJegbEgaCPmk69oo2G6do8W2lRbVmVFJmrPDMwu3ct
ooMs6KrDExnWFEvg3CLbvthzAQnOtSfQWwKH9TVRk5EVPbUn+6WI/7hyIW/xdnc07Set6OaHajSZ
BCx7UCyt6dkpz71bKzG/U+gCVmEy2o7wLoXk2EArg+H7bAYjyevniVfilKDiiddKgEF0GSN61d31
E62cyoQG8t4xyvEjEXIoIMhZK0NGkYAsnpkM+zkNCthOQxi06hPEtZ8jiePqNcGfYZ8zCOrBpRhw
Izo8ZFNp7a1ilJ/DpLFdP5vzhkhyVps1oqIIbn0+NG+FOI8J7TP7Yciuvd22Eql/9fVwrs8zfC8A
vVu1bVlv+TtExGS738513iJrMuLnSBHCnKtj36QMVcJ9QsLHxehznerrfrs6dfj3kw5kztTXsXLv
JyLeu8WMhCa1Hc7NtInDi0y+moD7SzJuJWR7BZtx+B2KV7DR1DMnHt5N7s9fC2M+NorBlkhtfcYc
nUZRuLJeJl1Qp5m5HMIAj/2gN4cAvTotNpokpajHOmhjK5O90bHn1LYg/5mVodepdM2i6BFxHNZb
qXLwoSgV9cwZE1FlClr1l39LzUgFFT1FXz3tgMXJiEXucq+VYH/v/sXki0oJy5UqcbjeHyuc8oRp
bm29XJZmn0MD/aFUC4mRI7Ap4+b7/kykd+qJlTlRLYR9UxW32ANsVjo/RvooHwK1CvGZguSCuPX9
8zTYKx2fpHALzCsaFl/0M9WBG5jfMTtzeuKtQhVqsqT3WShc48zxn4UkJT9ARWmCA9FjNcsirvZD
JjucKxzVYFbPdwumpHEsF5cGHotFrAKwOwYdl1vDtaCbG9wUS/X2mr5Jv0noEH5B2LY5Qf0oq4DX
Zi9H5JWFAgiv6dhQWSjo0Eu7Ig88ZgvaCwEBQBkQwWGKJzMMTQAAYHbJ1LrGVRpRKq6kziNU8y7H
93ld6UUKNhAuGPskMN3aaziY/7QDXw08a9lUp7Pu1XluXPV7XjQ0w3lXEkJGOXgglqlqykxpOhYR
j5+0HHpnNTXym61PhkizWCX0U9j/1bYoBS35sJh3uH7vgShxRfvHeGyKlEA/1eaUs7qHe8gmiopx
qu3LsGR9XNKhai34jVBsmiVKolREM2leeuk+Nj1asP18iAXxJ54OtpfjF86KUAxsRerQSCQQKgZz
aOO36EodZQK6mThBuS0yavcPw0iyoe33tIE94Hme2zDDWf5CW7gs+iI8yX90UBbeXQ4u+jmFf+Ue
PN22+rPYeLIlSPkbHq7VTl4f9QMMicVDBMHb2kboBr6qCIornMucJKeJQhOsOL2pa78LvM4F3iIH
/81Ea05IaV/Aj3EeibUgBx/grhNrOHtzJTBnVLjLp5/xojTEnPFL16aC8DKbHDIkoS+TgNgJ2rOn
LYA4pvEY4p/9UtYi8g8KEc8AXPSLaRsgdLJiq902CucMHV5TT3CRoVshpQ2N+NX0S2wcQ28mqV/L
IAyC0ZrbcMvitgzg6i/8/ivOQaHTTcboRnbmxYVqT/F8xrycgckiO6jIAhonsnWsMWCusRRxYApV
DBs1rd9LrjUfTsZrPcyX0I2ZoQUoI36v8BWWKBc9pvt76nDl10Go5GV6EQMKD+i4XN+DVQUSKu1V
c6Jhfs9t6tTALyPlBiEt4Mv1Zkr+4B5SPqLIiLQF3qOvnjAKRTVROtCK0ZuBsDhOWF3Y3tofZCH9
y+tu592didwyfcmSzNTAQRT2d0Dffb+kOee0POMBcE3pCQXPnYJG9rgrz86Ycfw1b/pCK10KAf7q
yTKHDzZzbdypVT5eQgNNWa5Xeq2TZNjmZp9hkfhN3vxIQzVspFe4J98zAOM3uET+ZiYxvm3VKhmG
jEJU2AP/7Y150O/STdRIXArxDQXm+4xFSyR2g4KwiA3+75Uh/a8Q9rndlbhut3ATUVD3JEqhFq6i
1ZeW2Ywob+u+Lnfvw0jIzEO++5GAU5DvRJ9clQoDFO2xrPrh/cjc+VXAr4AVNxesTPyg5z2ZhzJe
/rxLrYfkZmWsjgth7yeLrl14Vx05sWQQapGAM8UdE0caAQ/GvEXDh8KXQQlAWqCc8wibWDhR7b5o
S8+qnsTstEHPgx2q4Ceq08bh1XYEcKHdgPfRluSVAPGcwbiUDs7vS7fFtsSWj11ZpHSB8e6kwy1M
I4W5NuA3u5vK4hKw/UYmgyptQ5DOi9A7ER1+NOoMMfqGE18pFLM6CGdZ3dYEp33v5NdwkrchxxDG
pj7CuP//MCIei1H6iHRsITRb/xuMNUCocqLA9FMjYHPHYcqI4xdqE7pqupsNnSZ+10Qre3BwG/f8
mR3f/8pw3hpFHhkpb3uN8jI1UGkHU9+OgtO/fsY0oO8LFP3lLHeWOvAgi+dit31ZEAfmIM0fT9PU
yzrZq1L4g0DhTqsJE0kV9wYVobdsw89/2RmrZCeYiBWY8zKq8xO6mAcPtGodDenbfY10KspKeUH4
hyWFjNhTdGx03e1ZzInejM7Qggy8fxNc6ODDbv7wpHsRr/Sq33UPI8W084chAalroMTe4rH0H90y
MuvgnWx9wsJNOC31KuHjLSNLhaFnXqDJSN4MznoWtwLcNITJmc73ohsrv5VA7JTNP9GI07FwyWdS
3e3pVM3+h1s3Qu+o0EG7UlksUA5+5Gte4PPpnUn50SHCKaM4i3sasWWOQ2ooAiMoB3Z5LN30Qeiy
rZsbHYwAG+7jgQCyHjU6weG5ooQsLXOHLOKRYvmxPwVhWW0xr+8431ORswjwuQdWzs+h2iXn5V5t
+VQbIxCODBQt2v8J7BMx7YrZX+GuJWiI7hR9Op2gNe7qrCn1c0KMp4VsyAonhnRVv1/0+oI34JDw
4rbRZA9UuuRUusyYnYwBmiHHerI+xWW3wzH4uFKcrJWP7KxIqeXw56hiCtCdMP9/n+H8ok5N9UYH
kpbdR5X2DrljDiAvUJGOzMbJB6ETGW8lWn8c0O8W/yHtVvfsrXSY/r+sMplmQb3+dhStqE6z/lXa
JhUg+ClqDasYFbXb90OrfSuKlL2QNzJclhKAZ/z8096WvdSx4XUbxjwSSeSjO2ZfkdhFRplVnBDy
9x09mUSoemaG368dg++UrlCYufvLVooMcP/7Np/BMz75uacZ30Ztg5JAM5v8+GmTdlAPaIjDZg2j
VQZeko0PRF3k3kHQwZlVf8MbmXd58kBLqFC8v+TSzliwoD3PgZnec5VA2VN5kzPOmxMdxSU+aTDm
2LFq278a2S35qIR++v2QrxwakxuM9EIGdkSfThw6v+nB7uMLLAIEgKD5pAS6hg/zywj+qo4432ai
6TQ7+XMCDIQJpt6RcznnqSHasK75fMxrlk/Hru657yTvnheOK+wfzq+762EO9c4fGzEA0305Ixk4
y3qqzh37djrv/NpAJW19g1nBp3EAu0Tf+yOLjq6vh1FV+2nFu7p8LyRI2OGIr6oKSfw5laku/03v
R2r8PHg0BetbjMFfZa0jBpGcOXHauVtyJoHBFh7+L/A02nO5vHiW4N+ltOUdxp1HGuBwfJv+rsWQ
ZHUGtL6Z05xnJgett+55ON7tMEUeVB8Jqqxo0BYq1+pYMlpWgKX0Vy9y2rQ3Svq1ZN4EdpMo/34X
n/9eeIbEnW46hRnKwmo8U//rwm+J0/7+KrodWjRLy5JYts1OhRvqzp/K5zBOj+mu/N7ST8OikTi1
meg+DA1wQDwKcRZI0lBOCT/NouHuLGGGQJscGEBxXXhnGJ+Xe89zaPrL3Jl9wqrMw9GXnwazonsS
MgOakwdbepnxGs42PJoH5wT+1F3sCJkZXaWsZ52zlubBH5WgYILIzuJvUn5yaxrXJyWfgTpFYONm
C8e1NXvMSVZ7prSXDuXg9I/BptBGqeeB3md5krT4r78JYalVU4pZJ+W+p7EU6Q7lmuPKB/Ry5Vhf
kgFVVuIOa+ahbklEct1+IRmq7hl001JVnp5+FSUQ2SEE93CsBPdSwxKFoXrfEOTjzYCftweQlQhz
467sf+Ln2gUFGa/BabFs/1PLEGnI7aQt7sj0xc49leLQYAVBe9IMjZb5eF2BNsGOPAN35JMP90o5
YcvGg3NkePuy+raTxd7PtoDHxF95KSC8MnkT17m1hoVzZubBl6laBzzkuW47XKjdKL/7rLVV27eS
ppP1j/8F/Bt3Tro/zDMdY7nAtH8CsKHM4Fl7u4rzXa1/fDdN0eWyGhJdybGwmerVRAOukOM0XMG7
hESZQBmtORpr73o0uJ1pDf0S3iumXqcyyWudAqky6FNtGxxZNHzdgZRNAd0/fEvnLycaxTVTkwKr
PfI0j+skxeczlkV7ptQwqwIGfnglc+uhmjVufyv9pwWRqCq5ggaoajYiMsigL24dStJHTJdu0uLs
dcnKs+fI6p23WjfNupUHwCnNIY950doIwmkQcrQMBn3CxhMh+Q/uQAr1xHrytYVlOLTW20pi4hN9
JeHIXqXlDdNDMSxF8WISMPXs6hFgmy6P2VHdJXOct024YAm97WW+0jMmCZzbj0aGiYe0q7/MmEv+
Mq77YtfuVFT7y/Ia0qi2KNDVQj+Uwkb9r9HrGCdh2zO3ZbEZmj70MjCeoIyR53wB17ITFTFCkXzU
LcngpUZEsZk2+pW/Gx4z1S5mTcQ4sI0xFdPZdiFzd8BgRIo8zAtmmu60nteSngzWooznEyJb6nPV
mGs6xLfE/aRijRcNuOVPatcnjYA0KTVeIR3+aCRCtvaHFuTnFWJVaF94fY0R0e2eUM0WWEC3fflB
HYFmmh0U9b/+EBjiBlqKDSido8FPlS+eg6KawwPnlP6+n1606yGPvond8p0+ovb6UK3j8Kzgv373
qJQOKUnEQa70SqBbkadwENifBWt9dZk/tCM67vlF0mZR/w95XR5cs+IFRB4hEnEZ5F4EGlEMC1Po
sumeWs01aMZExsCM2edu9Wu7sLDSgv9VySjasE0as2WY82j0/0opNcz0Y8bIh6qo91p9CQ9V2eo2
J4ZRr/jBuAMMozyWRE2tyMEVPzyoX42Es2zu0FL/QO0rN3J6f75AemWNj4mQ6Upv5WMkwb+/MKrC
eli4V2TQ9DZoJDb0Q5Q6D9ELJYYwJkua61HxFq5OdIuMHEJfCUVvEXgD7k5qGkSjyVGUZW6rA1h+
MK+cWp1ghE93Qsr3F1m3TIFyswU+RAxUaYqQgOlcqxR5aY+tEgDcyQocnEZNdHHLL8gYJL9ETNcl
ZUJ/pV5haKFGgNMoR3fx99wqoCW6ZDwXGB4w2AYJ8kC4emrqvbw619SiFB74DG7NhU3kLLr/0eJa
2ThnREdIhCER94mTjQDt+pqqLpVHD6yScCP0XncvFropbKee3SWhgLeOZHkwly8lPmC+/LSR2xcj
siDjPJvyGd9jNNYjSbsDvP68AKSTpLYrjLHhUEPrGZDyad3Rhm906XPpxnGYB0n0SJWpOajBUAlt
hu5s+xC3nJm3RJN9ARo5Q29ZZ8MrCEIdq0Ny+FdLJM4hHm2Ky/dWo9cJ6F/ABcOmATl68nMbmuN8
CQ+GojlAUavVXcJvFtaSZ7P9MnjGLgWeVOztXCOVfPvaGcyMo1EDVRyk13bgkVWI0ZHplRYtT2Rw
AlNQUr2x4dRSd+eQOf+myqIWrKCFH0kjQvPa/JRJhRYa2zxsVtyeTB3eZ0JUIfJAlyCnu2JpML5u
+ZOV0BJF1/dVslsQWiaLwxfid8Z4RxXwBo0X7pe2VUINVA26cyxUUi1SuJVgko9gTlqdZJnbKEpy
u5V4qEE2I5E0/GCwROX7sQlUBsfzQjufKh2ifcUbmDRpIf+hc3UBXbeb0GGwQj8oY2Av+yANUnsY
vjx5Lc8LxiP7tYjkW2R2xVs+MezYJK5t1yGgFSY8988MmUMDNhFcn1WTHh+3z0AugdtVEmBaEl/f
3U4ODJ4D3+P5MyXGZav993tt2B5MZxknBZMhr6WzgQjRbsFaRnoNvnWKUxjF4gr1ozbF/x/xpKqw
XxVtVtf9q7RPVFXdAs4wnRzi4yi655/jcj4lUqZP92Qp3BQ8zQWW/i91XMN9rktqqytHXSnexyXN
NpCXPmkPWu5S7nPSn9XSQsk0X6jZp3/lx2RRIseb2066e6PWV94G0qgrtXa934U3Dx3KMjP2HikU
yx0EaVZIdQoU8gTeTtMZMD+YCu3dG9e7x2rLsc0hJ4qfUuPgKEwU8+g5ogepbkZKf4hbgdMci64C
w39X3chdL6D0zX/ZS9HkdL9KLeFjJQcnV74x6r9AaLuCfhAk/FBP7z4o/gKGaeDcvhTj0bU8bSJE
A41vafwppf6jSMVT+rMnNd8q5Xy29xZPUveCDrnWk58aP1tbRXmc+nNTdpecDCukKhUZv8lzOZVL
0zJyY4KKquBkhP9s+JBQJE6zfEOiUYqdFv6LXLz9OnX0sTIcGHjHC9+u2cG1QiquL/d6WMWJlkIE
Xlj/JaYgrCLeCvykcTC+Rpj8i56rcev1/fYAZ4b6FOh1uTbeEhViVuu4HQB76/4R37oDgH0OC1gY
+F2Ag0C6FdwJZjwfPbL5LF8/OgH1xY8YIydyu2pQST1g9uKDr6U9M3cp/i6R3dP5Atou3xFwimLi
Fc2B4BLziXcJDawDpCTWbvBOUBWEcuKsB5xjQmL/sE7MEqv3WS8MtHlbdC4gkO8NNmeMCjysWOVM
muUg84FhzJYh7+D9+ZU/eQDpGJM3SFpaRT+AmAmhVFbgzKXDcOBEOMfGgXm+UK/TBDMVG8lr1qfT
YHrUVdD1ol4/ITgecOo7NxtggoAGfFBcLk3JPa0Zx10/ZQdkG6eASRU9mHBTf/62gSkXpnC7rks/
wX8529BkzZIz1Yr4a9YqO59bbDMwYYBDzKewUzEJDkMOo2/FPy1XixOjWnlw2bntufgk6keWau7P
5o1gDREfQIIwWLGW03+/RVL569CTLIU4eTBCyJLXKfle3x/WJf+1vLcwacO/lrOBuTrXALLkk5Ou
fAae46FKmeRiaIeLt2dOyOwBIDiWHeC2ghOJIe/9wemBZaXSVefbbUbGuYIbYxut2YSqPvy/iuoo
OlU9uLx2vmH1j7x7TLwmGbOK1V8XJCgj22roTsWiynYqq5NWGNec0O+r/jXMVY37/0JpqS2tV1eN
W8k4JQd7a/Qyih1mZOe1JakjjGXSYb90F6Z0IhWIz+OH+qgVju4PYD550559+S3o5uJ3RoetxsEc
XBuOQ20xQqs3Uma1FYuORwUo26VNLw+kEjb2tdD+9Umva8Hcy1ECHSkSB72Qw9tEAgImD9trhfvG
v/dCVjS/yOG2Do+7VKnN70T9QrFw8ph7McsJ9xNntRhDpbAvEJILOyWCrSt7vstUwJ9TOKx9t2Rv
ESNfMDED7oVWlAiLFwafEp0tWhnfjzh6vLtZlvaqde4CV2xg+NmtJ9ah/e8+0pPWYItCB85jrt+P
PmFm5tJMPmq4ABN3SE3f0vC9Fb7RJYlVYtNRH9xaR8hiagrKnRYU6z7+YezBt7lnYaxxHBaZNOCo
FIvixPQcu4cJBUsH4XpZwndXRPC0HT+ITDVs3eO4tGr2nkwT+YAYQjlQdKxmF8xJFU6jvPv9UsbY
67ScSxgkVYBArrW+UbDD6AwTE2xMT0IiMaxbIXD8vMMdWNHoUgIVqraV1jqSlR8f5cjGI0zcgChw
R/6470mIAgU5zuEEbNrOn2r4J4rkno5puM0FOeulN3XqS/oBYQfNQJgsyWTcSSOnYHMFhHKOjtnO
cMeImblfbIOmg77pAsYft5tuUN9AS0mwv5Ofr0ZMhiJwQm+sJm7knkoXnLeNDrOg4iD8s7kVA/Fl
B7uRzhrOx8XAJ9Dz7emnee5jZKh2eRf4rU9NUvM91agWcqaxsYoW9dv81/QDIpkKG0z0gwYuy4CG
Pnl+5hkczp3ThsyfHEwyTIxDwB85zfC+Yw0N/ezAo1rfkNAe3uydphdvgVnToMZFRDFPhU3XYpwS
7WTZkJz6RNoTy5xQU/mj9Y8202MOS9DpGUNHKGitUSciPCBoL/tnPIQpmH254YLexudUn4A+uNiI
6kcdNQeGJFdbFT4BBNCDQRb+ipmN//QGrY/x9IJWAb3t8LXpECO+UrFkk08j6kbj1lTisLaWDBa5
0SKP/g08XbuyoKf6CipzMHR+pSfbWYXUKxhw03tflUhdyqosldM5j657yyAQ0ZsWvYehlwAiUudK
lPAZdam09iDqEf9fD3tiAwVVKshNz9FJ0TIDHM0OVh2yA/4ChVwaV95jLTLxlPCp/TVJsr5AOJyC
WUdujHSSWGNwQVGaS+v/qV41YcSpqRPQZ8MrOCOm5RFAsxVTx6zLqe/wvrrICHww0RFKyPZbU5GZ
XTvOsE9XXj9WTBFpu3nv8Y0OHlLM247Cm7YT+2DSvw58PWoVmmXVuIRUTC8jKKz45kSZxAtEQ6vD
QRoTCKGQ3dC5y1O9hcD5/+HFmFizZpE18gi7WAvbHlw24+pEpEVJkfRA/rpC6iLJwSwlrXlENfIj
m203zyXKArkB9mwnyUJsunqxJdAbLKO1f1UVrjCmVrx1Qq2BvLDgKBdadue7PlzTfEx69DW566JG
8iUVbdLkJdC85ZRPT+KZhXCgAOEdX2bdbA7VVEjTRnzavSd4uAwJBnfif1p1+sNN1BLxsMVwHSKl
qQZn4H7CMUI+IBluhCSsduQvRzg6CA+GJB/ALqHg7vIyl5fEBIUTpGB2GjrrCEN3i4linpyoMx7L
xoNr9hy/PTND4ojLDt7ZoSR4eb2XflbfI9jYxCkbq48e+ucc5xZL313Q9V4KJQ4LietwV1W19xU/
8+QI0towJywaVAtw3U0StrRpV9T7BpBt+EqymGQveqDEnPWqdN8U47AEHVd+Jun4Yxgt4/98sg6r
owGq2cHzdArNNjaCm0byRv5DGGkHodVmaRfDHqPapXeozxnXqc6UQ8SGAHi7i9MEYPGjs9UhXy6t
If/9hXCfHakA5FTMw0w6DtQ46ZhE5pBKJFPgzGsujNpHhAEgmguZPZJQHZo6yK/Jnu3YbqGsKChl
gccX9UrklB06mJLKwjYH8TYzCHmh61skGnVUX3Y4I2JVtreY3SI4OLw9B2tG7qCgUrSRh9AgZVlT
Rio9C6YpwL5d8EcY1ixiz6/fzJXdbChp6YtVcAz5c/WfCl9dPp9BCVpHgdRH9zAReRa+sc0NmPb6
v7PQ+fNHMpKXKNp69tfvtRCqj0eYZdgzKnRJNYQdtTttlbmaW+lc1ShRjLIfanyypWWnkwstY7X2
+WbtEB02zHNyxSI2JZAxtpwgbhoOOWhn5LRjZXsi7+SfVPQtQ3aJWTzpA9uMLBb1lFJHHk6EYcqr
e5Qz4UEcN0ZeH1bDvd8TDbjmsy99f7E4r4xUme6YV49nh32BAzGUdVWju67GEi8BtfSwIBui+MDF
IvvUX9ZgOKSycnwW+aKFrr4oVgPimFij/2iIipr1kHrw9+3X3puVrtNWVRY0/pGP4AJQD6d3pva7
TWIqc81Ajdcfqgc1YUK3GSFJ48dnt8AtYMoVEBTH3puWK6uPRVwe59L+OCVdkxMWGEA8sklig43E
V7jz9oDtfUQkzTvHdTtXtF24o/hfzqavPsaUGE4+oTHRGb8OYfgu2ln/CljqAI+21+oaci46Y10d
ridHAK+nEpQ80796UK2r0poM+N+5S+8JP+AI+iu0QYDt4K3fS6vg/4xXo4L8O9ZjhFXVFk6IpJpV
wweyXrJzq+7JLV+WO3RpslxSlsiv97bSpSZygoB0VGbMclpZYXF9vEHcE01qa28ZG43EDSTjQShs
VgIDaYP0KqixXRoNNAsSCOeKXGFdbggma8xQ1w0U+k4JmULhiC+LI/0W2cCZAuy0kkTSAv6HByy5
xNYw9xRFTckVTS6v5xQjMJXsyZFdRtjFX7mcHQSB/gukqNXY45ObWVZf8SPvyLaRiLGDbu8ug6U7
w/POY66YaUHDcF2eb581Aj525AhS7Ok0m59ezAhi+bpR55oudndNcdoswJW0x/5V5eqxG7dBbDjP
26gBP9y6V9E1N+vUIUWyztZirgUtIUyktuoFvud9FhWoko63mzTBTr1YIUYFgja094/voZvAB9DC
OCMmF70/bpPUJjkg6cx4mnkPpgltXm2CVEcD5KYgrLQorvJTlMCDHOzuvuWiTQ/NquFfRWCNCFg0
M8Zxy6w9jt9ld+hrc8QbGpHRFZvwVtbn8FZ5o3HRvFo5cHD2a9s5gx6WIoatVTPoCgtiFM5goyw4
39eFZUojrHLJdbNP93AnXSq/MmqFQGEaM2Lj9ofuYqwaEiVrG0aXRqW/1VaG0gxvEUzr6fOGnOf9
cEbemz6djgnf9RPANl7Fi5gU7hmZ7mt1tXWXMgekNTT5Ag03vcrYZMVJVFGeIk/ntHhX0WLVZ/7c
0b8NK3dJzV1BqmAJCGo8UHCTEWcsAUs2w+5+azVKHJm8H24dUlGQBvVwne67OQPSod/E41rTmi5f
wC3s2yWjiswBDlKw0YWkd9e0J81PLa6FS0tkBcryAorLUo+Xe4xhfBzxBMl2MizdzCS3kb6a1Ydg
q+MlMzJiU+DZpNlECtJ9xCo1qmlFITYx8cb9DM45T4pO6E775BzCowkUydXbFTSfgqMX9dBr0gmR
9Tp7kbCV1VX3VjEMFNePYuASIdpiDF0cn53AgbneOv/eZTnaTeGOYaalTKiu7AmaHz4epm4bwptK
bKT5ZiYgizYgpm30kgDmiaSPeXIj8SYuQg0G9utx/42+9A3fhmnUwyo5UcnaMhPA6CfktVGYWIVh
/mYkqZvMvkMgpNrbhg6y3Ym9IsfIs2pZcL3s7qgI7OVwkQOszsYAwqIAz3V9MFoITg7GGbdjiZXf
aKozIOUbgqN74XnHQlpIdi3U8hUkkoDCP1W5VVqkbqqCFz1W4VwB74EK0MEs3MhJjloYQClDE5nO
xMJJDYLvdOdqK0yGjqAyHpPfwTJGInHEj10BlAsIchPfaHNy17sibiPBcAa/qNCPaEGVjyw0dnl5
CQbXlIC3CRvyXsm2iXADD0RTw7wAfNyn/E4ycyRqwsTvPYt6FGhwEBUqEtX/LP0+7QOwEeEVDjbS
te2SbcAChQbmzOPRYGlEwFbHwQIizbG43lAbhnqi3c/DdraahXKx/WF+JCxfw8QzVQalA14x7FI0
TXwFUgFL1UFEtADzZtUAt9WsFSUJTvbesqI2ABmP+4XgLRlLSEG9Xterv/MLG2YThN22dafXuPJT
LwUxmq+VHXTPe8kf3IdvUZdxE4WLx2sRRhETwaOhD5DSXEKxDze1k4Aaupr8Zqjp9pvdLa3ZJqkk
lVRS402bF50YI07TfSkcso7HOEZL/ubkSS3pMYYzXPmREXoFwO6qFJnujrUudJRhCp4UPyaKLbK+
HaL2OmLyOmVWEEIOLaUBQTLghL4Axj3SgF7IBCSpSB+aa/cUsGuTScJ6Rx/+1P8u2sSjdR7fNkBz
2shdQQdzZ+VPHMwW4dkNo9zqlrVIrSp3Y+L12fCPPl1pwqsE3FBlrD1KPoPhwtPb8E+FBrbXTgD8
TaSLaFFdSAsfG1Mj1FjNyChe5sIYKo5e7fkSJ4vSKmNEQQBlx9uXWVmxfq2rWJJNC3mDpSAbLAb+
ULadKmaO9ez0kIufyHG0MSc3lLYdgH3NeSL5Icup3dIeBc/M9Ga9PvAocLqjEqtRI21FClJ42I+I
0KZz8V118hi3wK1dVSZvEo4bwfHjtKG0CctReNOSdDt2btfdzAPpvhx6raJJ/xgIlt0tPYayds3w
vJ+RMiIipDRMtGnESNnz6iyRsXzYza48eGuCwrK5mTrigEKvKWER0FnsYqqAIFgFvemkAEK8Y0sK
rmuktpmvdzexoCr3cg9wOvXqPUILkhSrlD0HEGNxHo/S0CVJlTOVGsdamC3XHTnNDFdiVc77flO6
ok3vnueWjY3Vxc+kRlpG4D5Rnu66oxpvaVNfIeL1vEW4BWdJ+0XtPTSC5q9+/wlHnRa0OzDmiopm
DKgmAX/MFmADgsnMOoGjB9iIBjvChCHts1KZwI7SduH9JByVUzkgrDufhG04X6ySQJkhd6qsAHDE
OTWlL8oFuvK4m9iPLf6ZIovopD8HKDfJpcl2z0hybxBxf3/KLwv5p1b81gWlsnVsyx7RU4xB3oJx
Slg9UDZxkYYyF9Jg0VE7HlHdJMZ5miebejvyhkUamgkN5kRWSx1yRQx6AbjXb5HSj82UH4ksmrPJ
8yLAnvac2AWB4vg920ETggiU3/6/iOqxeF/LHae2pHhqb39EcLrgXm3z2Ved5MSpy8AZigCn5amP
YVXbqzDIwln+4x5RnUAhyq1VJJr6OY7K2tvV9dl+JOcy0PC5DX1t96TdS1OlNTUae6KMd9O3Mzdz
OwGc+4QH1YxrEORg11xoILXDKDF1/2B4Bz/RdDhvIU5BSsewRICJTM0LuFeWNBMP/vof/V4VcF5c
DpJiGtPE8SOvv7Dog8e7FK+xW+slAAVI0EpaeRSSi8T/Giq6s0irDO8PGCggQAyHnYoW1oMd2aGH
cN/qP8H/hXR1fL6uUfifokFr9Mf/t3SqeA3y/xkNxHx2NotqbDQ6rW5GensZYFAkuGKcmjhCQOJq
5fkxaE8GmJ9Wqb2ohAkPbzpZD0bJ0s6opxNBtxPuqOGrRGV7HX4ASe9QjuECAbrha7umTQsSUQL9
JSNML3XBID6gVSC5YQWY7ktPhG3M1HfrHyzAQKunfW0o139Hk60OB03TyInIQD8p3Z5XmeKrU22s
gKSWVjXW0F4m3DWkPUyf9W1Q87YyBwVrDiXOaYtR3pUww4zSP8aex/JJX2pnFrvNZ+Fbo/BR2FP8
9z+u+ciYdLubfbr8+OabEskaupeEBvIyFGZPpVRxy4+I7QKTzw5T+sO5+lQ+pKLF5xACZko2yU4p
bHTJV7U0CkMK4YzcXv872OhfU5IVKfqVGekJSmmcGzNEMF09wKHyHXAPcLyo9OmhISXTLy8wIFJV
4OE8VWaC4Q9IZ7NY0kJPco4p0wdr2ADUSkWzXWNdQR4xhNmM+OqahADHZfTUg6e4EwSdTjihc2EB
T3bfnJpPHOgPkb9dXc3Bs+MsLE/RpXd3cO5Wwnaa4ungTRXF+q00SK6G60P4LyIJcXpRYhde0VAF
axvlN4WzRuoOYHOvNJEhbMXc9DG0Q512ZZYi/BUNi8M7ZulS9BSO7kFVxKlXMztt/0MAVuoeK6P8
wvl0C7RjGGgTVTivzREvGjxhrodiyy9GmH7ZoOkwF6CL1AQOgYNH0xnB5tPmDTOtOjhjiw/uzkYY
LT7tWohq3qRr8OGWR6MtbnhZpNn2GT3BA8LLHdsq2YLtN7VfH8rw1b1fN8F+jzDNDQo7p3qDSYNg
bEDr+cWtm/jlrDkUuulLNHpeJSkoB/LxZDKth2XoXGiCs9HWR28Sf+DezZUBt8OlQH6rJc0lEJi6
S6nCkfwF+3xo0Fk9nipls+6C/Pj4HLVkGbchHEOvahesq7aJ7MuosoFFkLTL96wvqE1DfwY9LXDe
IrrnrhqSuLI+ReoU4LBzvSMTi4+DQ7Q6vPjfXBnNB3sMZMAbn3S0PL0MPFJs8g/M6nY+5LPBHRev
SlUS6OVWdEbw85de0oP9spEimfJ8acNXegC7mAoIWd6uy08E9iFcqeSCc8Ge/1zfjZ3PIAKbrpy7
T6fnbzOLWNAuzbtRmk7rN4M16SDBiF8lir/xpHF8oWrCxBHkrN96zzWzts8GmKXIbDN+hqIpL421
IIo/CTCM5oX/QKUXFeb+gsyzmoRHOZyTmDohZwU27ZKdTBxocX8At2MyJNfP+xYQf/Nlib0azz7X
jiluQo2pf8s68PxztXIns3mV2rCZpsGjmTZiBj54OQqujP9J7+o3z5gAaADaOx1k98xJf8sRKFnF
R4F/RZiiCgv1UyENUaUihaGjRYhawuHDQpyJmGwqoDZxKDqjDJ3yP9bW3nh5aoIg/X+4xZ8iJr+d
soln2oEABiyUGwFUAlVlWoVvmQLdbtIPh/AwNutHo/++0s2vlCrBtbo3czqUZV0d8FD19k099LNq
mt9unxZ/Z+aPhC1J3FVYhGbEeK/eC2d3+Hgb/h3wniN8m3+Qc2P7pH7VykaSJ/jbizK8ghXUKY0H
zWgOngseLWtyYkHfCk/xgmMq76EufoUf+kVDPs1DGSx8q/MOJnsU2l46f7oVcwyV6G2NOvqgNt+z
IaSutk7lbEJzYgtkWC2d4LFhmIUr1azkTWnB0aynBECARFHdiCW7064W2k8AblZ/n3XtIwUFFGDR
W1Ga70nY1XEtgAlVtRpfo/Kopcp8EONyVW/qUniVAJokOV5tdMUtbdT3KHn0S5OHjVkGgwOALRd4
W6SRS0UfdzKu6oPd1v3Ij3Kg96XnXWy+vPpk7N6ElkqpM3TVU1I/EoLZZ3msbWqHO5WwKFNcPR1b
usRW7qMewOUBa6WuhHh+0pX5q+zn1JE/KG5hOQE9+3UD69BJRMUCTLOSqGWqVOnzIquQTaCnE8ks
3vlYUErIltCuQnq5zrIExjWQUVYfFz/+Wh4d81eJOV5/yerfFs6xjMb1n3Gxw+Lg6pwKdPc2JTUV
6Xa7jY2NotkmxNRnznTTnaBJ9StBylr7GMr7RxQpDKngKyswHSnmaWiGLjAa1PD/MhWd+hSh2BHK
xftmBcUAKBMhqKgjBZBnMmiL3d62hJSIhUcEFiWIiWgeoLIrztfqxbIV2fsFXVaiGRUKk2xpVF6j
XgxFw3PvM5n3/e+IMgCDWtfUVnU7Qa5AzY2H0vuHUlrLnkAhjsLrFszOBweb8VHBiUyI9JuYa136
Z22EyhDyNce1iQkXVK/WVfmjU481WLv8vLtoYr8c4jwtN55ageSEqwMLeoeNIcEIQgDP9gl5TzGS
v2zukJ5NXOQ2imuRWFBgSXkFSmTJuuCXaviBiHbjBVIMFFhlPCYehExCufsHz1KiymrLbhHgoreo
WltwJPekxeNprzLnHs3oI2jcWyjx9WyEM6JRypl7YM4szEP+7mej/O5GRJ7OO4g5ps4+E9feLp/w
dWZWm6xB4OeLqoycgFq0dBuXBEmEUwojgtA0XRIPF+vP0ixMV/j+SCfD7PGtdxniUC1h6SoiqdPc
T7+si97CVRs9djiNl5PikTvxuuf5UCEl5YTytZA7lHv6fiVXUm2RjzQy/QFUGtxP5xbDlvXI9Lss
EbFEMEB2dm0KypXIptCvlWkalsQ1Rl8y6u4PnL2bKJ5/8NyGfOZXs8AJN3yUpfxdCvjJ60qeX7YA
xM1TFP2Wa03NhR3rkoVGUpYUUkhCfXN8sl0Du9+9gpzmDFQa0cn8tbKblJvoP2XBbeP20tAsfjB3
+BeYE1UUQLpOo4jddU8gsbDzI2RuNTv6inDa/Fb+tpJVKEv53WVZBRoUs3WgFv/LnEcYSqsd9ndA
87VipQ5y3yUgAd9fVPSA3d7DxbeSs96BYH3EvkxPvjZhgAUWAq+HqzMUi7IMCiyMTU5Jl32wXOk/
abTGAYQsVGjU6o6yg5vFHcgs1m5e5cAQTOmMLEbzUZTXKcYL8JQwbvR196VGmCg3QSePUYVsU4EN
vx2PozYUHnmaahX/ZyNpuJpAQVwEVAA504A6NMzt2D5NmD8D4KqjQPtm5A+in8LudwrtOQRBwaD/
eQfwXBHyRNERkFg7WHyqDxpzNRfiJV+FiuDZfpdr7zos/xnwRUAvQqFpF/Dw/UgYAUhIyt3aiaTH
ElknCREk17YnRIzIr5VSoVStQN80K01Equa4Igs5IIameQn5Xhf6g6t5rmCJ6z7/HWXx/EjOIk9m
kFkvnL5qiLE1ohJ6rSmpMbOmPSZ064NP2ekOEQZGPMf9H1YlPc0QmfcoEKP2x+IJPs56Rw5KkHGW
XJQHEl0O6sGNlSFbrrX8cN6Ik3vDmf4vpFderJCeAvrhTb9Bq0CFyM7qQD2oqgmRnV3XFqOHVT6H
Hj73U5ViLVYsjiTueN+cRa7D4/TvpZOkfB17ubIyrlBgrSP7K4u1Pn5/dlNoR80GCVqXa2KXfb4k
2nKevQPXd0UBEXu4DzFQSFun/IBmvcoi1IKsbsuWDP2lRFLaR5pecB1r31URRz7cZy504gMtnDMb
OOZUxZ8ialPYCjL8RkZow6jVu3ZiC1aNuKBZI2mt7pYXKxg7yZ8NzMQ8oDVbpcXRg81sSgqB5b6T
Zv78tdq7tqJQEkZ1Zrr1VNpZ457Av21yItlOnzghCHeqDMy5BxZGEfmCInue3zcmuIpc2LrIOTuk
iloH1nF09n6cwcltucFDeMBm2vgYXfBXJkpKhqPI2qJzQG42UxUEtdzTy4qHuxzybi6CwowBLa65
FpRCWr8oznju2GcBh1sQ2cLqdmuVYX9JmePJQcid/lDeK53BBZIq8vW6bNo2cyzgeLXX4no6V9kC
snUNW+enolDl98siFPfsssCBpu3W3aaqd4OQcukpsX3crrdLffF0kNsEQ2bDgH3epPyVt9ioSCT6
MV3Ui2aTjiocrVIa8IfS5/8GsMEUF6G/ZLuIPW4ryyuPjG45VRkfYFTJJRvyJyKJ0+YYB7ELDqu4
VhDPMFH4bX/w/BFLf9Dk+MO0SCeMf7+z4a4aouQ/m3Djh61STysbf8F+1ENlBew9t5F2H5JW+1gV
0sM1JfOcIcI9HMQGtUw3AT3jm8mglb1GWEA8uJY+s8D41UVoCcCYJvJ/JX55dFUbdsCZtwDFDNoy
+zuSXi/dJ1AJ/6UJvx8I2FqQM8yrSHGAwHf3ZOQ1qvg0d+ljR7rtUzs22CWS5jvtnHLYFtOaIHgg
YlA/K9jArKKSidNIYuW00Y+Sus1UnPqcLXVxjF1uXhXqb+npezPNKaK19FTLHRZQI4i6hA8h0LOO
vuLV4mkRQKy58GdzPNUbHW4J4ior58H1x7V/iHGLOkkIdyZGn6SUs7YDD0gRFPpVMZjgK6ANHqB8
gr4sJiS2jFra1N7k0adwK1G2cYQ1ylWyE1OHKXZCVlyIKxPs/HU3wzZ4+Rq+l6OK5kazaa2VAGMC
x7lmN2HGBJqaGjUUKHM0zURGbkZMvP4b8bdidsc9AuCpgJyV6kiDVMq3nLVLJFVtY0U7B1dR1bdP
zF+jtfJjP/RqBResBP89ICVWx+Fy/PmZXhogvDPTXcIaFQ74W/bSbj+D6lp41TyHb/8cDo+B9tie
8Ow0RNcet9LJyUwRAtvdY7cDBkSM+7fFb82CJnRnKHxPZlzoq7cMqET7uadsd7urgQFMeX6+cTqb
ziuNqnzVVi4nmbyTYV/gkXsRgEO0kGuceNUKYoZDIlABzYmvFpukv6Rl71N+HKeo6+5PgPrWcPO3
Kl+CKbHlV4G86RApioTBuVvBxTALos4wzmjy/YIqG9o0506HdRH7dBMLnTX41RxSHiqd8WyYgkIF
9TnqzlbPEeGUWejgmVjyU3pHm8aBArgohi4OFkl9aqLlcwCD5aLisdoL6bQlJS3m+iB6/MuMLkgN
IJC5kLL/bAcSbO7YsCO5Gt55gUk/ADGtTZ//6ETdZkgItU3jSabl1TnzRHHAnB+0lLHNhByF31aN
sZhxa2rjAibVNp7vpuVfq58e7C/3m4GXTSllmi650PYfIDlpsOr90UQPlOzjtDQHTQjy3+ZPq9sx
poa7Pc7UzK/aS8gO6+0YUTvTTo7A/t1T5C4HoKs4b51dACJKhm6UUE5B/3I4iud75vWAlOe5ysVJ
zvpw4wzxnHL5Z0sjxS8qpnsAVAdOwY2/0+Qw/8jIq6wSWF4W4vmhIVnyvixGp9sFfFr8AaVHbiYo
6cfWrZpdx9nOX1Ho1JAu/72nyxSLUWN1ZlPCMRH6ec72jX4j7SQ+uTG1AHGlsNSO4UaJNwV4cTgu
LtjGuZdJNnm7ZSHbinbRPmZHxTvKBuAIOQ6yuHwkDn2mKNm7UsnYHp42M8H3UekAGF5c23ERx8MD
4LCmn5IFaVT/E2hBqz+2/bF7b6DH+5+bwVyMbqaALdE6QrUnDgbzSCdE8k9AJR46wXcRWo/CTlht
pbQdgDD1LW2C/deMZjs43BTxOrRsp2UbGc9jXuQGM4L6bb0HR7p0ZQTMiNpjx2nHqfelSOx78mbg
soN3pwJ9m2SPYwPUh4R1mr2a9n1LlE6HQNYFdBNpwI1Ny+fpTwcWa0l1jiaZrfjbfrg9daZ7Jvpg
FioQjM2F4UzG3kEa1AmSRiWnv/YkAKSnCepnTNhMtbcb/WcjKynNnajy1qm362gwleo0BnYB5OaS
blvZcgpnPjWDT2/pU3FjNjcAdECEGLscg6DToTLKXbfHY1/54NdRWXUcoVdHPIdeeANJOOo9EVDU
PTpq7CSClWzuVFSJHQzlBz5vDgiEm8cmRx6JroWxSqB1HP2ULBTGah/dgVan/7eOeAHdN0pHfTAI
MPRJlIHymQZ0ig01UvTGmf/zJ4NU9z86PE/aOBVG6xCZl5kFqMyajXAU83XZtweSVs2Q/LSfcVIm
aSc2p/weA1MbLrmGxAdgGOgwvPp/jQGfa/9VWjkdRKhVMRLQ4TaAsPPyVNKOvQgRn9BehVjEpxKS
o6Qb9cWrf03572hA0H5wq4B4iArqCHiDYdzoKpo6OheXQgdLoAlFOmF7UbxYLgFDRT4WdkOvw4sT
WWVFy74kWVNg/9r7J7A9wTobN3SlCwMN7HhDy39qxE5y7FQOyYszgFtokp9vrHRWWXh7Y0zBs7HE
VZEV0kWFZM7p9ZGLPDJ52TW+81ICyBt2EJV3QWwN00CRxKMDMTsFaVYRpU4BW+0JtIX/Ap/X9hBn
/1HPZjaB83F5oKL83r22tOnn19h1icfof1elAB2u2CSo3sPjTESmGo2anWE+TAb+wm9izjfJTMmS
JHBNRGqhGYECE4sEPjGnMfpThFOSJ9H6tcM28mv9fmKvKDv0gjo3gS/C4o16aDpl6cPBv49J3HXH
taVGLJY6l75RL3Lgmn7kFDd0vTj4yZUuLk8JCJUn6Et7SPoi4TIheAwkHy1dl19n1O+xxacAk8LL
VAgkrf7mBscwALJDiFR+BRaiJoWSdTpSmZdqNs3xetqt1/MMrHRv8q0nQ/3QkyPJi4JZfSE30C1V
m0y0mn+5+K4RxILVrx6cz3reg1rQVZ4rIoBFEIKkB4bZ67xS7ogFFJQuIcRSebOMr4KCsjVgAHJx
yycX+ehWrEZaXvls7BDRbRfs5rWagD6IpCI3DXriGqBQXhfsYTKaZwkqxCOAwp445boutHcJPdfh
oy771EeFHeg0WPuZta0SP9qJksPrtKtECS1QyF1rJme9RI4dPjlsV1PFRy9w7AAR2sqoLRTGnsAu
H1xQTKCa++FAzqpdgob+BBhk/KNwxcRFarjNLj1c3i79uW73cEkHgrqIxawWxolYX03IuzwsgiHO
7555ZpbcWfAVKTuemDQZ5I7avTbeMd5ZMt7laYfZiYafVoAs39Wwrux07qidItMV6flNrEA/cn+z
BwF9TQJpmk9cyAWjYNqd5aRBcWagj3RvIb44SCmwIOPV2GP+upYvKNo3V79/XG5rOhY7a008wRP6
W9/Eui8nVqo/U5uODwObzemtrqDbOCqyK4njEw9wZhLFGYmb1HSpvJqWsu79zVcnEeUSvE77xNQY
6qmMd4a8+2g/aYQBsB0nu1HbrXiIzdokLcTKbeQ0ts/PTA4jEOYguqy6PJmYN+pQmxNBmzNDG2Ix
0UOM4Zi6sk06dHJGRNIMpfEmOIbuostoBT7HzNM+aHb7lQJaFPLMu73BBnpf3H5lWHMQFy0P8feZ
D0jglItGI9OKkIreSNcNNCg+6JgZxTEwCMVyYRoOGeXGt5GV9GogklVA533TmklAlJvp6tAQFP+G
4wMiYQSRc+WPdKxWkAHhcqMlgi6JEDwgfTzuPT5r+sfUqd0rzCLOPoVzPUA8Zu4KlMgLzjHn6Iiy
p5SXbkcODznpEBNcyHf36zMV36IU5FouVvb5aebq4892KVntBfxx5EnkxVwjHFm5avrD3fO0pAHh
7UwKyKcZUEwFcszyD8nVVw3dwf1nAISBR2lNZQy2Z1JZAgW3iUdvqU7qOgA8GqQuvn345ha0zunv
a+kCtDmLGtT19otNyB7NzSwiy6lgJ80bWvMGug0Xs+vxCevSVobjTMgz1SggGSD3QP8SH4jAZbCV
U9OxFSUJ3Oxur2nIgZsvFdYhiRuIhfZ0RAsU3NOAnjf4sLYz/8bX5UQoq61TpwiRtSvugU/IHfnE
b8COnTCDqlRqQj/txwgd27+cVjIr5Agg9iDRHUtXuXtufOoxjKvTGSRFle9Vq7SPd6yCEX+yBhN4
qWRfA4H4IOASkB26fighUQWiyKevgBQ+9/oQDiEsUZCS7MT7vLvBWy/AOpMMVsVYDy9sr4zWf8eI
ayfSHtDBmOpNhg/XqwxMjyZpXd+W1yaQczXnfBI2T6PQHbE8AvOOpgaisseab/IhJIDNrB4InW57
7D7vktPIwHDPbib2Azp1SLwHWEPojupFLNqo9hDvq1at4LWQwLWJEVlIT8t8YGpI4wtXOxc40vy5
MhUaO9PiVn2Q9rf6CFOiJm36QJX5LrpgJmh2KiyvKXFfl0zJqVxZnw3cqgRDx8/XcqR/ceJgx199
chtGFDiaoxjx1Hh4wPAGu+cLo2dSyHVTIFj3HzUz6bDqyK3GTgUBSnmNJSOj7FoxiyLguUe/RaVY
7MGyolGbLWvL7zf1o7ju/IqhmuBC8kdzWLDV9cXV8+1upHkzXIPYddSLzOvgCcxxSZXqxejwdR0h
3154cH3ilEkpTZmllINimGEWpeMAxgTcRnln84+xQjq7BRsyftItvg0JIOxnaMt0VhejJ0lr+9X9
cDrLKEUs6FPGzF3ahXUwuZRzerU/30/XTcShQR9KCURCMtcAplpf3ZvQyC9a+3NBTBQNc4x3gUr+
Dc9rZzx4fTOAdap9lWDfxgnJqY0lzHx/XdWCsv1mb3709Ju6UfnN03KaMMKDtKB9hSPipe/m1sKf
nCWBNchnIBCzI5XY7JT27cCh4jlJ4xjUQs0m9yRDKNR+rUermaBUNEy/xIzg5vsS1C0XdKQMH1GO
4kHQ3tHEJ9lTitiKJeLmGV1Ec7M+OrNq31CyGyFfRa5e2LNHsGyL0CllPr9fnVxptVpMjNfv9byM
0l+RGDh+sHMcovIQ2Y+RG3oiwxBLjDA18S1V6Zh+8oshfZ2UxjYPQoRLE5HJmD7QQXpObSNEoJqk
Xwmt3LROb4IxhA5jS6I9BTHiR7qhlNQ8JF5HEQCgrkRfn/8eXEKTqnis2ZYdViIC88tqhXaXYgH1
5IpiaGGWIHzVfVGVYqUAjvm/l9f/p1LAcBygBSKqrhIiX7GMd8deqaoWmrBhLTYZtQZ3UwSvzHI1
aUIewMOWZVdvY4pxh24gkokUPXmTnHZQSBRZ3vEk/9U7nHrOOJwgbm+kl1Zbu2l8GNUZysfCsXM2
KtHW7zGSl88Su845amY2JPnWpCBxQweJ/f9bBWmHJBYY04QjInUHPb9fCC/9LJnMOOA/+tF4CUu6
Pn21IA3syu5W1tc5ZTgiGXBg92S4/sTIWkdMj/eGNfgG4RWZyNOD4jAA+kUetXwisKWBTCtHT5gY
xvYnY58KYWw2/H7B5YbuCztvKIql4gKUjsNKiX1cZqqjkcblPZK0zZwcwDq+ygeRK8s/oIY8Tn8H
mFhVPfyRWuU3RfvfZyXKAOLsHOIli/rqXD1lUyC4UYl7aWjQX2Hg5s/W52RFlJabfwf7pc5+hUY5
JCHg9g0PcNT5MoTtCbyHZS0ZhckPbXoaE5/UWdpfKVsb9Nk8AILx0HF3t/1FItOvcGFeG3MpdQol
ALBCesEEBzJCm51qZXCx8RhiRbaSUZEJzHoQaVehKcFy/w8SISo93ATsJsw/w4oa/ScnEN3roykr
JAZBwQeaTSZZbq8c7hRNXHtWD18WXVvPQcahwrB3Pjsa/AAsa9a1qeD+H5SHJ6zms5fYGRNIKjNW
88yOdFSaYFUcfnhakO5Gy/0yvunOJ8/XhW0EAt9z5kUgBh/1u3joADy6CJeTaDjdRrsm5gjswNqa
gv3OzuWHy+GRjAgA+EL4InXFfJV1qujhAjn6V9DMsgdaR+XbzPcCt0L/mLvJyvNyrOTJOIb58vkc
wCoJPA/zlP+Rcrwhtl00lY6difu3VzpIVDgUrm1VPHgsc4VQKnqP8X/zoetMYQjz/izFv+WvSGyL
DFcgc7shiNZ1ta7C4U7Ek8WH6fMlGZLSctorZXJk7oF9adNbVI53oOn5hbiol9U81h2u18pW/Vv5
rebCqfxU3HNGIKFKVKcM/hPFXu8eEuQkgVp4lHIWiqtFW9Z3wNMI/CA/s1TztP3FG2PFWsoQtLMT
LRB/RnMdRuhRc4hG7whv7SL40DzxBCfkxkGiOq3tZFKJ8ni9pLjAjnam485VNBRpB0h7iNnLowjA
IufxoG/8XqNctqO2PsqJLYe84Ka0bW0OYzcLIrgYpmHbFoZvcFUUjDpZcbsUzSlUTS1J0fdmTBJW
pU8TGUVf7B9SCwoePLNgCHMo/aYyVD0G48zkWyrPFi8GaoMPxXA4dGD2Z0cDAekA3oF77Dl66r6x
NYlFgCut1PSkZMXKW5lXvH1vHNh+7FlT9WbNkoBhcRqAIcYjcRyfFJe2R+2+a6sf1Ahr6MIvRe6v
QAObD1wZfpkfO8+Z6f4tFvRKMIVjrjDeLUF/P0Dg1oCyjffVJ0Ffq4Xu6uhJEwNjnwYIa0z9inay
hxAI09UCQJ40Inwg9IpvXkV+vGn9XztnvLQsLc9K8iaMwX5tdpD0K/MLgE/uRHDjhl27oVTFFzAR
kUGeBuQxCnerfKrPv5wS906Vj+xfPmd1c5G+Uti5DOz2qTkt2k7Oys8oV7w+tluOQSPippS8FKEw
NZqVOqjKTgOacpiaJyu1MZB/wg2GvwnKYxGjpV/Fnv55kONr7f1UK/915OraG+z3wSlOuJPVKr+F
hh6LciHHpSqRz9ZYvK7RZXUDTRYmaVrOlgZM41/SKqRhrk5C1EBURKDqBFojKT/aDqt/YP/4iXKp
96dDrrc+x8I/PaAAciQgOEix9QekAMa4DeTaoRMWbqVckvBWc5nLRI3cvh0ba7sQVSP3PDyvFRit
VcgVR/AMUw976Pj3uaAkhMTradWLsF/dZH5ZgOLnvW6389+h1SHtNTRmj72yclz9FB1SKm9ttEXh
4CcXH4T8G9N8nKFoAigOMJy2JQgOh8DvU8cUVkWWs/ZLSJVsb5bxMJkoYz0je2oYmjiXaxo+TmVr
PErv8xD9On5tXmue5tQoAtjU5VH4roR1lsJx0iNyfhlcsDevpUrmbLe8lI1lqlA6VzeKSTPgWbaq
ivWUJgJPdnBab2SkT+omAUVvgx7gHth2bjoBBmLQj4g2HBlMUdti9GoZt4Unte/nR4S4If9VfcbK
TSlr3Ihq2PmCBd85FHko9Kw4PVLf2fUfkTHImub8HTkM6hZv70KX0h4Anpq2i12mdfPUKmG2SIe9
DEgyJgkUa0N5i0Lmqg30qC0LVGiM6ABRwxHZ5QBKHgvQ1dDDZGRcWBuCBKpR2K5j55Q7iu/xYeRQ
JJebMd6fkoZYikosbqra8HXskTqGdm5IZfoyAkAwya1RQlbzdAlkTrr1Gehaf3waWWppQdg/yMT8
O33CUAKNCgmmgUh4t23GjIWJSC/PLUO4CF8YvA2RUteRH+s/rpoKgSRthWwM9C13zXIvkg0+G6bs
G/4E5j2O9HWHdsGHpzShr/yE0bX9p1f+iLFDnrydqYQAkTnmBSvXT+WNFo7PVFjJNjmIxr52jS5H
4oxrTtUx1Li/I3/+5MAV2Yfm3ZfAjkkdUlWf1TM+APKz+TuVVXJpSFGlscegA5h/kL9MbWm1ajzm
79px3cfSNBT+5RtDeEFODBVB8nRUpaZS6L8WqGVuY9C44Cu0wHGzNOof2atwVX7zrjIAykPzWoue
Bh2KxX6LDMlztojqmRPWzdU4+gGHe3ttx8bhvCj95sNI9m1XMZgyoMvZJSYc1iwIyLPvDXynV2l4
wut1KHxL1p3rtkOmXyOz2tUk6R2/uOzNHrLfZcQPfzJTHc9095KezrOcsWHZh/Fkk91kcCvgENVH
tz1lovU22BN1iqM7KSk59+9amj/nTxRJ7lVZ2iH9mBujY+zR0FtFJRycT4CEghx6r69TCAIRKcIj
BHfDVksxyLYuuhDJeH1+jp/rQe6HQO9EJJm4Yw/AaMTQM4sKmgdGQplSAp2rBpVT6c+arxWGLAMO
8ADnijxYU/Oz3MvfpDdyzhxsTqOPuc3VsxL+6+071qEZRgGKkbaMkAxMbnPxZ24TKaHNl5J5Yf/1
fYfIl7FvmCSAjFgHf7fB1FvyehmDgaYs+avufP4Y2rkkMgsSp6B0/0dXVVgOvtBIfP0ajbBSc/bA
x9OdnRsSPBt46rzNy2zqqMxlZ1NFiPDXo8+tshBP5LcngRUa07XQg/mFlCMaX+gSAMlFwuYENZCN
os5+N+J9ZHKLlr9WVygrrdqbYFYLBkCy3M0+spz0OLLKxpKdKZCER+Cird3eMrmy4VHoIZq8PGXV
wzj4cg23/9dJywdYorQUoN87PuqIPi0IoVUYrdJXueM5Dyws8/V3bbpbts92+S5bZGcZ6Qjzb+pk
hWlrc9aJsJy7vjoZuMdEcH4W+HwbnAQZL18d29XaKtlla5ev9HYzDKjkpuN8ISOO23Vjob6IU0SC
qaglLI6VosEwgdByWE3QwFevLa1mwcL8M4LIkEn5dO7cO0Owo8COVSUV1tuaXJa0kDeb53o3pxC6
F/CdJqPjFvyNJX9BmXl70XgA4NOHB/w745knhIsyCdWWyzgk1hb4krRdbnG/HqAy8bG3O5gfMlAF
yzI6S6rxXfxvXZeyLEzol6mikM47aT97O+tjOorAvmEh7KD7mRQBuSS1aY9X+y+kqIbwTHpIwQYj
b/g928gI1F0XlOa9iUeqB7/ZbIQdz88/vrc/oESFZNbtMuQUCTj95f6n9mHrb6+kfd2u/tvgt7XT
hO7MmLbERqfIZC5oGPQU/fUyKcOFQAQJVVyg+HC8io/cSq6nYwCNCOsanhrlQOwISSMD+o3XwW6c
gLE3WvfHHPfaXyH/kvrIRvQygmpjM8fZz7O8f4RAwoxqEm1XW2PR56xjdiHKqFHOEEpnaGIhLu1X
b4x7CjIVHhYoa9d8rcLZfYN6aUc8xDSlsix9q4qZ5Yf4a8mLwcPW6oZTT7b8LA44PPLGk/K53ljL
SyzMSGdQoI9cPsETRi4LRJx83PpU5Igtj+ppVXC5ptbvSRxUOQlEecG1gPxoczW9qIuRGrjaEhlX
MYEDr8mIN669rvc2x4FAthgafcU+dbY2qPSROmH41usqgn9qj+V6H0fNR+7gunvLri7pF8TM2xjm
PGFacLDo+L4gnKD3Q2vLUBXE6wU1+fsOgyJEf2fFi5rlVWSfUBvkSW78sTMcI6dBCblN1hv8eQSu
ruJFYeYPop/rHn9yA1dty61mNNpeIbwJ8R7HHt4D+Ok6IgiLbuYUdRHG+uhiX1www/3gmxb42xTP
UuRBNuq9KM24CnyLM09B5CHFz2XzX0JISYp1+Afxm4mmQrKuHIbLKAIjsf/kOpxhEZZEPopRH6R6
4xgiYBgTfmtkP1mVbefo3f14zsSerLUu83ZkdgZEOcSyxE2K6wiCmdoxFomniS3USo4pYnu5BCyt
NF/TdGwFwg0j4AoSzVy7eQLdE8FCm5flChpMiRgqZ1sO9PIRVlRelSMcyOOFp/ZrB3V/+Hg/6s53
qpix0EX3xW2YWtAihRE9YJd1VKkf5B87EvHE9v24Za6PAVubfZt2WHoC3rqiPxa7TpA57vOROhVK
xleLhNLHFr6EUa9/wBPriJtP4sGh4hjUAVMUybZMIUcgkz9/Thv54SZxtu9ecqqwuASVRf8Ltwom
BF1m2LMv7HtEf0KY/tGGA2h5voHjey/MAUWi2535qMai9ZSBWJEIKMt9Nz84Vbr+9ReVf0DexblY
KFPflP8cLituhtyT0qnVP+LzPYuJ51Iya+vH/dlcvsM7zU9Hh0hbn5sfcgADVcwZxKehwnIu19B1
PVC+QSWBIhK57LH6q0BSg0J4oSgGGlRV3D8Kca1vGV2gvWhrSV9Qiu2XSHeGVWQOfedmFmowHbrJ
4ZmcriRWjTJhBoIOZpgfeOPllKO/cjGzWWdHz/2LEGUMZO/8B2fNbVksu7pFJpQaBpYWvLCAdQ/7
8l76c5tBwuayBAdlMHj/8aM8KdN0zjy2f9VmXtbYsmFSfCHvcQQ0PiH8r9B5C/qOHYe7fS0stUjj
30PldvrNXRSv4qHA6bZEoP8wxKtwPLCgPkKEeJbCfXkKHwgxE5GO5yFVwi4mblby3Ff0QYL7xQve
/q+3mfrge/j/WCHBaIBfcrzWBl12juviWGIrr4GmQImERqGAKs8x/9doQpmES5Q4sZfgFQI5VnK0
foxlAMAl2G4oXEiiBlCnqIZGyw4ptt/7aFRO0NacKXmBlq0PLBnQSQG97x8sT1GjJ+JEZhYC1j4u
IJoMU8K3U9v9xwGFT3gx9gsXLmL9cx6dVFizoo5DIRn5fsypJgMRLLifVjvOaFMwkLvo+AW18HNx
y3vw4axI0OhEAcyPMPJeMUzU9tv/Ey7kNdlc77BXCrqQdz2sCrCF5Kwm07m7rvu9NDbycnGIAXSp
ir40LdzlMh52YgPVu7hrzUAFBwbZaoC8mxMF9AHCadR3DibCv3rue4YSInMNI5+g/SDTMa/pgbLm
+f2dkCn4JPT3xvDH8mjsd7eyv9r55w3lrVLnjEyNROAr8TS95kGQ+OqF0Kvp2XVH4Gpz4ChnyLhr
b0MJhsmBR3dbloyV0gdZwzVcTG2NCGFfSZyvVPiSD+G/Rki/P+bj+Cz5/wggb1GrttdcYoEbSkmK
uxJxYM3llKdwt2G6mCIE0Kizw2WqaoaIAsZO9VnMJXdJBd69q0b/aB5znyd11Fa3EzQtZH/ByAZx
o9jMj7FRYr/gjwIlRU0zEg8C/bN0PYGPlubAdRy2UBHnMDX2bylmqMnR6S47lok6vtka7nWxiJdF
1ywYCOv1UzbYhmB1naLly6jgKHaOfbiZMO3CNsJCby6VwYAr2apdsv/UQJyZceEKAs1zOweUepqm
dd/PgUZeSLa8e+NhYoS27qBXK+HToLYiqAdziEBwaz4U/no3EgCNYpdT2zGCUWiqnGUf1XGno77z
AJ2i9ceWr+cAaWJSUDVcdyEVLOPOJY2HewR3mxgl3RRWVTkNcgBK37ZMtSnFNZirHyRU6NGvHNDH
BG7nJjXXbqehJW8NpXfn/Hi7u+rAQNIK465WTrDvqyYyCFtrp184GFQGfsI/Q8kPoZljq/dSi4G6
+FpzX9ldvp0fZ0mH3wmdSQdetC0mwh9vYvsw525vAnfMlJ8QLMaTGwcuOQR0j0Nx9TLLyDGT05rH
ayXyNTWMDuE3fAoifXZCeYewklAlH7gdCsX5MwNrHh6ld7OcQS1iJCiFivXi7/wfe76xF5I1FtiM
Uy4UV5IDxqUAG8AUqtiQwZ1IqXYPwWKOYHnBw/fwVg++h4pzH+uTmtRDLoKZmguhQ5VUmeMhmmJ3
q5y6cDkcO0S5EgERBXkfePuHNWwfdTR7JVN5N2Dh3Es71BdBUYTPA03hZhVadlZElBbkTie7LHqA
qOQYKA327PKAz+Su8AVy2G+URbG7vurceniejl9KZlfBXINuWK9QwzVPP2Mjjw3AhjPIRwQm56rV
PixRhJAaIOwZ3glu+gLUkEMuVKS4yhV+Fl4rY7Jgdh4VplSFtovGEYhwJxUR41g3Dz+K4A7VvK1f
aIMQViEMFf6/33nHi0jshIJhPbK1YhBNyOPGMPO7XDzs+46bmhS5JwTH5KEkYl8/hMl4OkDo4DRW
0jEQxlF3Elw14+6lnf9WtM6ChQZ9cbs42XJdC3xr1PoDGJsz3NEL7C6V+TGNVJLBShFT7xUqc3dW
7HRsTb7h7MRN92ipYu/9Ywtihv8Hkso1Tpxi+01qQTaMNtqwh7qTOEINaxjLIfBi6HNEESyLCZW/
fKyeQ4m8+FU7E0m2Bj3HkDToxPgbV1nAkygzRAjAZc7hajAYg0QpiAX0MmLybZOCyajWCZqG0gjF
MwuyjyJJ7CkfxUQQ5r6+iswoKp7enXmBpcXF3jmEVCBxuwALFcko006M8qh4ugmZcNKM5Rbb2MgF
VliQusj8cxnqrcd387PwuSajiWyK8YRHq8vfHUQ67clNxkhGLeZuR3Rcogz1pGg7d9EvETnUUerG
37LDgWa99ozVjvpEfgX1gFe+K/o8ACRHqEY1CKPFZ4qYixNcG9AkT5Ki3R5S2hVtIOckctFt5WUw
kcSSIuAoHAiPHQ1kI3RetAwKQyfKv55LerOMUf8v5un0UieMKQcbaoKBlT30v4thkwnhbTlk35/X
BwD8hM8tr9xt0lYkFN1LanRDgDFFBg1DRnoW5swlr5zQf8x0S/hOPnAoKSRN6ImD4E62IOdzznMU
jLj8CGVJqLtITFT8DLw5MMzNz9DQZjRzC4ilDKbfbr7MnWLOg37xGhWOoZQ78JbRKW4nf2LZtxjs
mOXukA+wZXWZbYhVSnE7+xX/qCYTLnYZtUOsGLLiOgIJIuo63dZHbqoLh084w4MKqEqKWFs6OShn
fyCWDweHWdJn9HmTPFidC/RTrWglQCjeR/UOGUgY23MGrMaT0Zff6MU2DIOmB2jqjMaRMOG74aPy
reSP2sArKeKh0OWVP8r2ti5CpRZdRXd35gqdj8KMEJAf/y+7881GSZXd0cnmmmQ7hA93bok74W0I
bZF6s+L1+cpsRFdT1wS8dsEbW2/vzNYC37AS3k+Joj2FfwzIeYnIXJRcCOXt7AW2QdOFRWFMXK3g
35lmddLZ8QNSJJ9Vp+Ab23k+yRLLgyJdCgPUMlkQUoCrSDf4Lv/MyqmUoCufMoy7S//3VYHjcoOL
GvnJc6r8PI+4dhT3hVAGyNvsL3F6J+hWLcX8LFIUNv/6KWLALpQpDtUU7q4aAtRIbZplWzQC6P8S
y7ByDX8rKxjukXxmW3sLNMCTzctN3Z74p1+9HkSclbM6e26osknxaCHXp7R2xSE5DKSYKunafy8q
28iCpADK6d3JWn3hPoKQ3ol2/07uGugviVsMoY29N4bTdvQAw6bK3L92vkzTV9lCiAFcOzk1XWUw
i06Zr5/pAgwNf6wsZNqYjIOmVxTRkmkoMgZ450CNPKAQlU7xTiXBp7dsBI+mBnB2LWRGuzggTqS6
43UxaEtlX/rzDg3ZBuPDd8WXu/6tq4+2bR6iGaw52afYgwQaN3+udDZmGr+QJbaNWjnBS8xBpSxx
/lTR7K3k01mWhSljgfC04jnhp5vHmBgQkl3aEUUgyJzMfVtLF6BmE/wM1pmpeES/0rYUluN7eQR1
CKDxGg8xz25iMHoxYRnstvnmBj6jQg4c5I3gHo1RKZhkjGgb7tsc4P54uHqy7QbhIZ4zBpG/HwYN
8w8jI3gd73FHlI3+gB4YR8aKcY0GTWDte2jKWmCwNHbVV6H18cgyXmpoFNHO2iV98MtM+mEQyG4k
mvLWv3A5EUDsSKsnDmInykfMP/kKy6xsjog3NCkcbAXnxCu6+GcuET6LLZDmqqG7M5VfKwY7Bsx6
YzMFsxZuY8pXNSta373uECmymVhmmvuzAaEZRymtIcY15wG5nP4n5pg1tBb6nDxQy7V/YxT0Ed5C
axlogn96D/WEePOHgeJQs1xGHyTG62cOa3cSdVszXQNbFs+9/sxRnmpgEYMtirq3n6izSRK0BD0M
wGalvLlqXdCwTTojX4I0yzqv04Lm52MHtPyjiOMCvazZBL9j4BQS9vq7Z9sXWyUSTI/z2Y9cmd4B
VXAT7sT3NwWpArb3iKoNcqcEiViYlboYhIJDOuSkK82Ugq2BbEDFSzgJ3ArVNJ3vzFGA6aU17Tj6
tv8upfFh3rmM2RgfKGvG5MDpBBCSh7ii9PIaJsfSjPgjupgX1MPAwuhowZ3VbcUW51MWqobgu5qT
6KjE8SP2N5bfH8k3WWlDVoBoV7sPCF//CN7k/MF35lt52AegzMLRORw23GTKtWsgBimT6TZmqGnK
Sp1clGfyoUQGhOAj7bU4Y5Z5+MADqPYk1NuUgKJK2bQhq8lD918pX9CWC+f30yB8O73VSVpNXbzy
mmtRE+CFCtlES5v19o4dDszCJxPxKZD/7emyl/Fzl/+8qga0LNoVU7H3J6DIPSu80856eSVBdHku
lhamfIksnbvYyJn0XY1IPjl49D8H2tCXmXX/PCtRk/78wOl3zWqCFCaPZgrKl2e8MUsclV6dgUdH
fFi2ws5QMx+ClrUzPOivOky4aSiGkEy/8ZUT9b5YD2cszsuOd7Xl5FDJeZj9etmcwFnICcT63Q5K
aESGH14sMBPPstwNxZKCWLoKVb63rEs/G1oZtQVBi6TddCefYImApLLZpfY2nf2oUcBMGF288j5t
Xjee+41VtdJGUu5Q86AQxQ9ndENX70ousnb2irJdZnxH13NHVNVb9E+5V/BmE0/0VA9CI6hL0aKJ
KsVJDqaxLcT9QIK6Frn9Jv8dIuj1N32sIIq4yx4I9vQEvT1sF5FqrGMQzxJh6qfji6Rd6s7vManH
G8S4QBUc2b/o0bmT+Im19nc3h8LsSqkZYjH0esIWDAn+b/VH7ecJx3GFhl8hw9WUTnbLT/1gVgnH
MQOLw0vtJx3knCYHpOtck5kfGOX0CJ0ucB/hMPchxdhdDP1XnLyZ8DD7hEzjXsjMrcXw9rXkiJu/
N7rZnes8dipK2L41tyZHyh8fUkKARGK/zPHJvqDd+XKZsv5PAeTgSU3gTv/VVvSOWXwdVHPAiLHi
ITlcWALbUah3/pDeoxLk2E55p5fEP8WzfG7k9TqYoh8SDiLLpB4vvtpIeGkqjQiCfultJlLyiiH1
gxXrH8wOVUCIIUFJHp6x79Q08xZ674x3AGCxxPSPQaQIrl7aQCR4Gzy4BUllO0LTXjH0KnuOqsvr
nX5+RhgMOyfkR8LNSi4fXHejccTen7xBoUwVgyw54ggpikG2uJCgO8/GxK2Hoy1/O8NkmKYhgdSS
SWJBI2G8mOg0xYI3t3OaIioe9hk9kmF/Lx2B/WvZ9V8GAMec/0O9V3HNnn8WEmHlcXfqwmulHwm/
kljTMI8LiyvJkj5meiMJPCykKTd79tHjnn7se7MqQ3QlZOj322s3e1kVxFm6mXyibOi47BQv7FVm
rSjyHYPXHDd2ehaaJRqIOT6kE3D2tNuhciP7Ae5pIC1fWNmyXLLhHKwmpGIned/ApMXPg+U4Mglk
lD1OE8pAAOFDVvVZhgdDkPNagyDrp26ANelA4i3O4nZmCbBCvMDsVPPTXwKpMCUQ/Y1BJYrUNimr
bbMaxQfmGy9R+R8nBSrNyE+uVXXZus7ew2mMI7ddbNdvtsGWZi6lwe4rhpfpCKHc4rHmikAaPzp4
j8XSksNPotVIAzf5bkhniyMESZGUU3VzGOYeaCfR++nZFFZdTjH6jTkr5s94jydlFqTtMkH7QFlh
Ymtn6ML7LxGBRukC7gpgOQzFDmh5EiWr0RVoa6TaXxg0r5yqYMdh21NDFvnMfjOGRylNSYZSEP+R
Yw6TD211DAe9O2qIC2K803K2SYZ8/7VbtDLk/mENUYtv996j+hSRzjqM6t32deXE6dU4u8R96QXW
PuaM+dxEnjLI2r3VummfxdrTN4EmVQ7gBOU99B0WXuc5MNPTBq6ndYmFx5bie7zCbnYPqV9vk9/A
kbrRAy/TzPluEZrnKMeQ8TeRImKcnZrBljz4QsoNDPk+xWxUJTjUsU31DRM0rOngMAR1fB35x/Sj
R2CRPYpJSFhlyR9O3D0rS7iB7G/3O78TDZ7lC0f0SRs8gKaKTRBGQoPexD1XDC6lArelt1EyTnAF
hMJeFcxoLYRFjIy+1tfvYR59TxQX+GYCV17WG+hHTKTKLdPO3rKW3Bi6HAB53xnx04NhHcOMkFyd
5HJDyDTzl4Eh0CoiwxraJSC+GpYRzROgEjKnbaW8refk8ETHH6Au3/VDDxAHFLdGjWPbu9cpVGoZ
XVSlY9sDK99otXSaIN7veaWpSl2o0qDk1l3f3MKt5rwvNDhZL0YF1mLJCQTnpVnHmxI7AthN4SI3
QxvtGZ0xDK+f15SlAuFgCwEVNqVkDiUVuBWtnxyVTSId9tfSDYRAHLONsPs4F+PM3mNECyBb2xef
QAS0lo+wGmwA9it6mZZSkGMvxzWSQ+Pus/o+v2RFeLKRdmvjUeS22BkCGbCNKU0OlZIbkkhALtvC
ECJK9uF6Z9wjJ6Ahpsn//A7xWBKyJBhDLH6P3ps90fwbnTJ7MZu9CZ6I5QVYzxqXRDl6YWnQzC+M
lNIr7mIZzKsxmtTN6WFbKLEsSOp2GlLyVLnp+DfnBDaBuo9Fyp3zrzieoFRCr6dWkMQ+/C1dk8HL
KsMZa0mw2pEa8zIsq3/0KIC36ErBE5sVG2gEBSRLLNkEO8i9SWnkbzXCb+8uiONedRkQiLLBLxsP
6eJJAc6ErHMDFpucqGfPUsVOaYw4E+hMadavLd9n9ZE8Xq3HgFm2xzf/XFG3x5MaZmDzU0ZJQ5KC
4Kpex86U7vn4i9VJ4ZggcL7Fs6jHoz0LgKkKV7Y1VDHtzBr88CC5GH5eoqU4nvtwxr4WxtIl5vEf
cYiWiJhLHGjMikVP3h9Es1bC3kWfybpFLyZNoPWIMaiVI/ItjoI064d1vme0GZLza7zDjOPE8ubZ
zcdEAcVIq9NsqfwDR8gzKMar7RPspKhSQn4PD8q6NF6gWFs3sXYREV2i4jvwFfv9ll9kVzCTtgq8
IvHpUlhU8v0pVVJedj4rlbC0mZtegrnQxWGW9viboso1B/YVlbTt0M0Etb5StOLaVf3wC9Nqm8ae
4sELGPY242AzAgAL1FkvzUnsxBl4f7Qrvclssl+9at5pwaZY0RXnhz2DoWsS2WAKnqLSRvJQiO5a
HcWzT0+HqgtSG1LrNefq2SvLCco3AyufcTWiAAvXfQ7bwvVgfxIkEOj8XbPBfOcEdN69OPJveB8f
Q8tDA1J7kNd4bWYP25b2qhjF9hyPutaXH/64/qdgdOx7Itwm/ONtMBxTKlHFaqymDp21IdMMqefz
wyRZ8H6pJRC/npbb+FTV2EJ92xF1gWChTFLCcUXSfd8TvGwSk0odG6dSK1HLM/b1sp3uMocb+q0L
6QzSl57kjK78Q0xRI9I71jtGbQDYvK7T72U/TUAtqkcwnlnqDoif5ILPyLHm6GE5mDOK15k9kVjc
1tlfAyu3N4AKDualXGdNkPGcq6ouNBtdyrBxHXATZoEBRYzYcyYcut0wh98CFC7Bsj5CuiAFi7ZO
8C5pzPSKZKiGmYKEhjABtGkgU5ugwHosi5Ryr92z2g9+BzeJuhIkNcFAbWKUAGF/yoUjx9sxSJ2E
b8XtYQqoC0GhXHEgeMUqEMz2mmjP4wHpGn/3QaZSaHJfV4Jlx4Ib3aPAeIgzTdrUifI3f+wY0lj8
je9rwNKAhpgrTwOy2fKdV+0NiV1aGXMR6/NqgonhU58MPxKVb01UPna7PORiT2jm3iPCXlRWl0Dn
NaslAUnwhhqsBxe+oFtBkP/XBLD0YR6XM5BQDQac8j6S5USYzwq4TqIu9WkH+je+jQfoEQLBLd1R
BxcCNMVXJits0oPtCJG3aRTrhp/H4SXD1ekSPLq/ApD8OvcALkC3zLb2pf89kvVZ6ScqrUWFv//Q
xgrbyEor1kXm9lOYTqL/CcG4XbcrqkprUbuxshyaIG+rWEtfkhnMNbEuWFJkG1dApQaXP3MyF1sj
fKgWHEhu+Q+nxQoJkNstqT/RCsd+b6iSnQwupElfZWPzJyxoQ80xfm3DZhxbRHBi2lJd0niq/tB+
uTVdi4uKjXXSV5hrcYFOebbGKbE/ZSYAlqDZqXS5bQbj8JJH3DXVGESI4xbTH1jCWI6WszuWvR5Q
objppl6lBcVaPpcZu8QYs3bLmID1MEs2VeZ7/UiZ5VC8yZL90fEe273GURCxA62RGM+yOdyaXrJX
3tA2H+ukB9NGJ8H3vicywyI4v0Zt2IcWP/E+eLBXY9Lsu7o5FV8zqB2KL9tclnKYKcSwIczCZNos
zcvIqNOnZn+0StFpUedMMC3UYpeIZFMkjeWDeuk0uNk9OgDnpNsVKg5PQcCgXin1lid5aSK/173M
ZW3tWPDh+zux953XOwXD6nlW+MeW5d3xLqjm+TBwBvFqO1sdYGTDqJKrdy001oqUSJI0RJEi0Ync
2/bWLbjRiWtNfO4ndCwUhHOeSb1DBB/irNGVMoWE79NxB66tNkdM3rZR3/0Ipq6IcMJu8KQav5+4
7jtbDK3K8X3xhUANCMbvk6O3a1KoDO1JPoNw6c30fzHjBZU7rqH3fwSx8Q96MVaLTqCHFOvXqlHl
sCHw/SYSkiNndOFnWk0Wn5mEkMJAXKgH27y6QQl/xiUi8BYR2h4DI74sJEgcMOnudAxs9jrxTAXM
+vO1CoJK9oQfNidSNRBTXfWuygy984pr3zoG742DF+qXQTW2+mjkJwCX+phbsxOzbP//hkMPXkQW
urADTwpPfhhUQNxXrN9NVdyjMTfyQaFsymIcmyG5s/1vG2Px13YZyqjUWZTsSxGWOTh5mMwEXUmF
AtU5bNCTJW9Upjya7H4pzOn+hfqZk14Dx0H24egMBAV2OxMsm2mZymO3q717BSl0inBPCTr12aW+
I1OP+Rq1egL5RD5e5RnY0Mwwm1XSTbPhMR8UBDj5OWzJwHaAXNA1azXVTfa2RMChEgjD31Vp0OdE
GD9BOdhrCi/HVl8VBitvu1CWPAphS3uGy3VW1tfoorVpvBvXY4kuENpiAQ4hkHXKF0eFgJhEAqs0
4oObx/iAZipr+Pq0CTZrRRkugxiP4k04IUfCgkbE/2FVQJTSYyB/Zh6tYufGSRlbmWDtjbLUX1Kn
JbOmXSUdnzpb2hwb+3oSvMtwHOZuyFp2pTL+FnFnKmR7emgve2EPRVK4TA3/YXuGq+Lf/m6p5m6Y
+eniYAD7Rf5lBE6/mHr9V7mvbb4gd4A7fCcVUPita13TPE3KDcc2btfZcsLW2JFzSGW93UFWK65p
CdKb7ZPGP4vErXamd0SVukzCIQaQ1FBaUWlT5P/a6rm6KFlCFcwq4psVADh8+CjvOWBD1xpk1/aC
GBfuUhc5XL0GDyvFdlORMG2eKe/kO5EfUmkwuj8uGVWcojMfWkmpL2fuQfj3vOU3KOShGxj133Pw
Ru+9tWTG08NwbVwBODQ2W5eHTTUmk7UeMhKWLijt3ycvmJHpYe1Lx6GPXhkOcWETO+vguJRgLVBH
DFJPGev7g9z51/hELfTwTUEtW0vxcr6Pfz8TJF+Sm0IrqsMsV/l7nKHREkxBo6CX4oHY66A1W+fR
JUNWXtdMIz40tzmVbeAcizn+ruY4510G1uoAbH3jjd8+7ehyV+0mnzl+WS9fiQxiSS9IrfxfyamK
ehUd0om/MGF4fJk3DuFAmZMnTNYt4H3SxWQumwmE8i7oeMrYfXBtgM/IeujiwduoH3Um5BFYyw+9
v9ANjm4jwJqGWPmkDePdyCknXIloLZ3hfVGm3FxQBa921mI3v6kHG5boFLxl8XKsJ1SX8t/RX3q6
GcjbfYVBj3UYSKuHOA3DFYVUYl6yrIOmE7x192ysTGvh/3oQSWiAgPfiyp++QPbvsxIRlCAyAEr2
yBMmKSnzKfLq46EW8EAqO1Kg6d4WJJ0Bn++AdYQQ4Ghv1airsxio2PjrGZAfVZH4Y+x3YCMDfcny
Tj3kV/QS5HsSIF05XdvtKuo17yMWxB7BoiWiWFWpjOiKVcInMzSamlSmoGFMa9+yAnYL7rOEWAv4
dP0Jwpg/kOJdZvovn6u2iwVpWsHTFhQ4x4ZnK1MrJKB1FszJ+H0KWRf+JhdpzyZGSJb6YnNHSl6T
KrayV8Ln9TSarZjkjHTrv5i8HOWWA4rUo5QtszY6yLtjeTddbMc4drDn7/fs2vb/85VGjdwLPWI1
Jhyw3PBCI4pndCvK9iUNXxxWCuz+TN4l46vGj+F3wLH4lcekEPy79sVhDm6H/1v2xSRtPClKEZgj
7VcGYoj11GJ7lRV8nGfaK2gvL/39IirpZDqOy7DZUcg50TUbVTDmxwpOE3bfyL/NYn1TNakmBpm9
1XFESLfb4V2ihPA+m/qaxVVKQHd4gU84YbpMtzpRUQXgfaY5/0cMqPByZbF6xFE5dT4Ynd9d2ASq
W6RFgZ8rzoyUlLt92Ly0zLr2MmSvp8Z48a77ayUfFpMXuJs9eGMidqEZSj3eOoT6na53wQGTmSDH
FLWJXsPC8EnKZgPlFWZV0alUWax/tUDii0kwLyaeOwVBmT7KMsdZSnC86x6abcyImo60W2wqe3Rf
gK4GlcPHyPkAH33+Un+KneOLDCxe7JzCgRhpY2YTrjcq48rOBvkrhRAxwFxCgM1604qP9UE8vtLY
DVsN1O/5xAaui6Yt8IA90rY6IV1A1wjGkNmHIXFIlOkWYG9X4uhesBENVn9qxXV195BmN//oOTBb
jGZh0HMEJXxazQOUTR7FkhCmRo9Q+vD9qioH511p1Q+3fLJ4yEhgORJsFDsn5CmwydXYHyz4+VOx
J53v8Wb1xO9dNl6Ql+mDCDvGa8g+RG6wkCpgkUdcVOy6Og762CwQSmd6FNwfuInUJGNKND9pbpkC
onWuxA6mgRWfSAgWgY3ISIl2y3/iG9rMi9iHuhcDIdofPlQJIv9Fj2AUgSctXmOqqttBU2sAVvfl
fE5e5y30cEjsEOBWtfeZlnR6+e35A7kN8mKZHcWdL58OHEHvnFX1ZdAsfSdZ8IzoSP7fBlyhTNhO
p0IuIzg/AzMedl/QYoCKZrrWF7RyotqAfq1xv5ODkNRDDF73bHOFuZ1VEq0LylNcFHC5okKxMq7C
5DU0rH/c+KX8GxIyVbiWx8yDsl18u1hKoymXKfo4VllJRlekukF3FdB4JqX8zGBKFYS4d6SsyrUO
yUo8wF9y8yx84XFRf+Q0zZnmnXaRJFeX1seic+oTtC2ctAiNKnxHvhCnwQzAR6L9KUe/gYZH5rp3
FOSCLjxJ+NSWd1TA0kkKoEsGiV7q1WB7uSQadv83MkaXZzxosmPbEZI36h4Esg9VmN4swRB36C4t
XoGf50r7+kl8vnYREBjOhFsXRODxMyTrHiYnMm84bI9/5Mne02WJJK5nnXYptzsqAtlRYmQCyLsW
YkXQIEiFN0QmSMMgLT9tZoORggaqjX9b5Dj/0KfiveT/yhPkR6EIhN+JH2P1RbEIOSy7RLLCJuJ5
VuSyMus0W3w1RMHuE4A+HvaWoh620r72K1/XsoTD9zUwyoKK2ir4cmle8ZfvxX+l6s2qVckfMdKM
yJlSIbQ2USkKOqcH2AdUtpgZT0VlrS9RhC0eZU10DURq8MBVbaHWYt88fakAWslqg1XdBf42FdJ1
ucro6fPY+r73v+0rtRfnxkJYx/9m6mmXOivWiM1tEbYDAY2ek31v/IT4+we3q/uPTt5kJxcwFGGQ
emIGWegphIGZVV3KxO2v/e4l1t3MDqiZKLCphS1KcgRUhqtd1d8rVGcHsK+Y0M5D/83mtEyT0/pm
WfdvYTehUVxSG6lmjrjeyJiPutzoIP9ATGo6xp5kAoVMrZOSQurmeO5XbZcPv4/TXgDKeyHKNtqC
/PeMAFjbfovLVkoPkmU2rSjR2w+josM/K3NT3fqF8k79LWTrXtdhxjervIvq1bv6aW96k3Hs/VK6
zQQPrPs9FWJ8bezmX5DfSmj6D5sqaDnSMuej9zKr3ur8+Q90fTbbM1uVkMtbEOwfBZOqWs7g6mDr
sDcgdxwHVlnqzis94DTDG45faOWxH88jYr8D11GyhA3ICXVvRnrh3QDXx6cNVbCYbqQtDNWnxUSj
Ll0dJ5wOe6Od69WCDIEdVYK0xK++0HmnIcU/2gZKQjoecWqGg25vkNo6e3UPuu7Hgv6XPUzFHbTV
guTi+8uuFvdcTplIS9EvEs9+Jsun/7XAjhQNhgyMd0dG7D6kxuSezWKM6z8rr20lmlg0JVcGYwsf
9Y4OjOQHcCZSxi9TSg1DirEktWZO+/A7FEQ79K+k/qt628FyEfDNbbAdqp4VUXzIlRSxrlAkTNrg
p2Oa0Aoy4GIkCG13Hdk6WlLs4cFBb83L0h0g1s1JRuAhVzK8gRZ39AMiXT81mpZOkpuTDDeQscpr
8XwcNmLQ5DPrQ0EfLbPUSR+CpGEZaSPszqtm3wOnH3Y9ocRB09gFJDbTU3CH0PS/a2cgqTyMncno
RBxjx8f4tdFYyHpwzObsdBgvkaoKe+CjSeU1S6lEZPMdvBaI0X6DcYdSewZEbKDVWqHLHS8/W6Lc
93ehRWGlIMWdDH0qMrR+L8ysGSG1PfKc7MVKTQIsCWkx3UH9MKDcyLIf3v6b2iUzyCKym0ePr8dj
ZQHHio/D4N/L58q2/aeTv2yW+mu2U744TggbTwCGzWa96oTrg70tM0L74KngfJ6smoMIeagpm4Ah
TfZfw5MbVKKg88qQl1XVLk/HQ0ZxHkMDXDFK8YeLYjU28LqsBYKgyUni9fTV1R6+Fobnis1t8uos
gJK/xO65k1UOIcwuRLqnDC18WfVvK95+gQD95t8vcGLqeMw/OUe+XM/krR4hKQzhrunFb46iSzRT
0FwMBgHyYdlFqiSG3CjXDpJVo12pEbHChWjuwZwpsOvxYxNqE7zayNIqdunxTa34wgo+jQW/CpXk
Uo5vn0/8NoM6ch3w0+1S8TqYRSTtocv1+8bnpG66kFtj1U8iGY2kceE+fV0iA4U8WWBmrMz5jfRJ
7BvNiuhvMjKkMDktqcfHGc/sA6eZ4ySh0BaDt0VKl8PqPNcx1mJ55SD+0fAnCXOLYtMxjhivK5ba
Q34dPLKGBdeUJ30IaGWQ+TjCaAypdiTnwUAMCjEQ/OSzXJHWnZkcuzFj3s+TdoFe+/xk46ezjdJW
NXKnDE/AN2tfXoJFHMTy8cNmkp7WP8/nJ9UQdqBVJx7KoqHVwpeADL7gQgmhjdtlJTVjk0qFC6A3
P/dIUxc0w+OsfhhN6rb30HWq0i2dQO678RuSf8wy+zKpFo5pYXX4lRReypnXdCvlYEFXtO7Abfrn
tooIOKkxg/WEQRa4MsYyQ3wU6hpNE1EXIms4cceMRsGXtnaTRjM7vOE36jd/Mk167AgvAH6Proua
g7s6tnk4yYSkxXnQ50UxD0UwAF0k7mBpqK0Wgy0WgYvfOHo5egNGDuVyO51qVRzI29yEicl4IuBn
vXpY5sENZ8NHuwaPH+EVvCRE8w6oQn8SwUznAI1SgUb0JVto8AcAgqQ6ba1IOAfKsORLAjeLZpsJ
YQ5p+30RsObyLsx5uocubsJSpNMcEtOKgDu4WN8eUcCoiiSNuXE5ZBwfVT5MEGaSAXN9Lbs33UAb
odT18TSF+hcPp+Vldl2cUlMK4CRNs1olB0ayFmjZInsA1+nZ+CHnBxEeFSR+2JOjIlPR+Mv6T9lx
5DygIHPLHLfMrbUsFrEg3Lp7JT7m79SzaY+/7icGNnnfqm4JP+50MvNt+wF+E512NWXvfGQm1K9r
rwVa7SIHGDevoXrc9gpcxq95RAWHMYTyEWa/4keJbN+1CLQQ92OXL/s3fQd6BRjfVRZCCVGALYvE
sQ1RUYzVdepUKTBdqXNnyJ3FXBsQ9hYZtsaPgTNU4f4Y0XWl3W69ZkGaYE+U2XU3ziBxRG35E/Uz
iNnzegCX7PNciZlCVfLe5JMiNbFwUEfM2wKymSy+afn+AtJrNzYyN0l5OQfp1idGt7R9gvexvV1K
hlLkTP6HkdUFb896GAafSSh4DrkmAzS3ieH6kXBKAwjr19fVhLrN2QZo6vy5Dx4QAw0FeUBA9QJT
BIlLWUt4l6AtuOG0hkE8S38gEEW/UtisFb4I0nwM6f4Y828XP+4pFCSKU4NCQeTcQlQgG3AlOR/0
H4wB2iEXwaHkPuXQIWzBrE8Ukx7Og3vQJC/7TUHE+SEEOZ3/KayUfInH/zskVvfBz/DuDDtJtWUq
1M8+AlzhwUy3DUQYqwP9qi6px6sQ7hN6uTgELxqjJ/ff30rqYDjeHZAfE5FxBKwv0vMawLNzHF7U
+5saV/3VGBN9pAzyIVTQokuZJt7Fm7INvlzGaNPTXXnBDJdLhJnW5alicDprMAmySVUXJP8qRLNt
oFxWrHsbSmkm5FPQ4KXfpPorMmoWHciHCP/DSslb/wYXxhoKx0ajGocZP3pid6SLuylSoM2AVQZc
zgZNTQ811jo2ebKg9aZ7zPwsuBqDzFM/dmVogArgj1WqJgzJClhWw0Nvw9hJu925TgQm6x6iAVpT
yhQlwwFIWeDjLEwa+EEruysCABsNIcAUwo0knkWOLTSmMCoh1RfWxO9fgC/Bs3+ZRJDFKuw9+Yh/
HwJJfe1aVPTrJCwYVw1U3FFmi+8jBAqIyyDYtkT/yMjEiJX29bh5t6Ff1g+Er5C0BEu9JsLRhImC
YXf9n0PpIrywsvxQUBIRWA8UxUOGXS09/hRAvPQQE5sIQeXIIZuKL2W4XmnVtpVnigLvw28Pd+jI
ZQcwi7bgQKYXL47/gUEFs3bi7m2HsXratZDlJ0MgJR1YUsI/KzqTG2KPDKf6JYs5jzyFR1qEfx82
5VnbU1Gtfeo3uATAyvNYtB2O1YuipWXM+HdrTe9e6oDV+yTh1LQJf9d9vaURtr+StVZ5BzilRpwO
52V/z4VrknviMXbCG+niAR+efcul3alO16D3ftu2605Ds6ioy0PYfTWonL4G0GLXhXUYDL2q4/so
ctdeFCVvO+hcL3JXvCtaGKMcOf6RAoA0NIh43vD1QPAr5PAWeZoUAsRe4tTlkab7kv2TlPx4liR9
8bytvxJPgArCWXLc7ElmCDDvpscTcPeJ1SAOvgaQn0n1w/iDc/SuyA1WKVGetwqz/1Bqa2i2eeVb
FgsRmkAqfBAMa8jZ/n/iXCm/eu4hIG+0yxsZFCwvJYJt+p5+IrEWg4qnZRSZMTaxbmhpFZo2U1Qd
LjWQNugNGafc9QU7l3vdQCwyLegkQ8p+CEeJXywhppQRscVhrDFpNbflJ/Jr9ZvEJwK00D987+0D
y97jSyt3RclEzKQWbJfGgmhMgiKmGY67/wXjKSOnOS3/R9NyaxVR/VjAHOUt3RPiHECvrjVm9DEq
tVJ0ONggXC6Yr69tPMSvqJFR9ceOsam0a0WhX04sfBlz9md6mBg7DGrezo1cD3qdjdZnUP0xne0s
8GAKQfOrFpLIZcAtNE903ffjFENn3XBCqz3UfVfn+cBVA54xZtVj83SqQK5NbEbthI28Ic7ORXT6
7Nt2hQ9kqkMlEM1T3aFtdrFS8XWz5pP4YiVkOH9KdKad4VGgR6qp6ChOU9THlmsumi3b2Q/dPO8i
bq5yh5LB6OjqAGC+pNKy5FL+eCCePevjSGhEtaqnBp5w52rkar7XxMXMa7iA8iiTTwPttV3EH12N
IaYPCRWdrd2H5WgoyFVb/71BGOMP9GeuEtdG5gbMirUmAyZ8tWZ7Q0lYAkH830D/32WQryd4HWsf
nqLs62jj1hk2Y7a7XKzvvr5oCEPzyCeYlEhbDagCVCgvAfwDYjr+vAj42J7zKcjPYVfI0U6u2WQr
71IFNxismXcCJrswCSjEGszUHhOtN9asFUGdHEUK2hhvwV1xwst/NTqDAFzpJtUb2zuR4DT+LsQE
fRD+HwRSclyk8flF6ncNvb/gcFPT8oBD05zCQ28Asmm8DSshSreCucVrBnahwes/owJOKKCEup5y
pfS9tkJe8kVDkF6BzDGQzzNIlxoeCrS7c9M8Gxhu2EjIUdMELxEgN90ul3FbPjlBH+op+eWq2lg4
/vHlfT70r9lKv5wPlr8XwPO6OW9gNqCXI1lFoT9XafPDlrX3xmOjmPkvPf1MlZRHJxdIdgpzb+/E
wzmrZW1Olrj9akVdhGC5l6P06XkIm64/VHZvytJ9khvvEW0mZIaLChku62OvxLgW8RenCMKrqB/A
XPzEVQv5gtk7d+wqXu9WiAiHdsqnd1rHf1bT+sZhrJXkdTXVTZsSLwVYLsLK5VDhnnsAVF98lqrb
Iquecdaq02/PJvsPDwnSaTPM+VPWvjut6sixhgs0w//SJDrPD5ev3VsWpxABnehGJKFzydexcm0Y
S7TKEPTWA2Zu9aDu3sPk5bUNfHDD8gysAd7p3bJOA6qnk2dn1U56xnJUA7hhinVhUWKYCosWDszs
C/KEQ6tgaOnFpaNcN6dq50kaAFvgg4N7oGRxWDeddMvWgJdbY8ZvFSeNsiThhEmqg221crCbAI0J
qJ8VE2GiFNWNyO97fHGcIq4k+tk3o8ZCdWltcZ0LbGhJBsMZ2NKzC53IjCKhgi3p88aV9DWkWMzq
wdsX/Edm0i7VEZ/23PRur7n5V7H7kE6K6m5MOTclwD7cBrP/5nlIwyYGLzHIhwjddpB41M3KB8T2
VIeaQygAef36PBuyoUIQ8o1/TWMCbr98DAA8VPWXAAqWnOsF7+9WimPe4Ghi63ExqrWf5OvZUoFj
66RScxpgagai//Gfh46V8DPePE40yvYrC7K4XyqYdEaQm2TN3ZcjSQR3iYiCQRkcSMy3jY1ltQ7l
bO5IWElF5PYL9gzf1drFD2d48Kzy0jQV28LcgfAtpu6X3QkW0lhnhyfnah1SL3bBKaO7PwHvYHWG
E6arXkuq/ZyBkkiOlYd+GRcfp0ysMOWGjTGgEztzG9g9fV2R61MUAiKplEOuWBkrqHjQ+o99iR+O
fS8XqSjPwrkso4ozZw0UvETWqlK9uXUooo/UlBIL+P7TynxCE8tLwp+Ff5HSWJoxkeA2hnirjmDH
IkcOHIWX3sLAmIOXRfSfAJrYofOawB7b5t1FrD/rZ5pB9w2IG5/C2g4Wl3dFUXEhG+9P5sq/kHam
Ubl6x+4anJYz+Gz3CntvkKPFLgioYE0u7kuA9B0m7tfOn2+zXBmnhkvmuDJSXIx2i/bck0v2oiVi
yK4QR9r9GJxFBL+MXKTsHtej/1edGxkcPvspUHAc3NAz41X1TLH036+faF5RkcZPE2WHd7ue2dIS
oghUy7Ltxp2PGAFGOPj1O5g1x7vb88X157cLUsk/I/AuUgmrjURSSjTLdVJs3LDq9tBSmVTnIm0l
zixM6+H3p0N4gWyNAoCH0KRhhtB7mSLSvEt86wJPCX0T8mgQBf43IxrgOLf7O9XcA6qWtVYA9YMh
m1bnEb+NCpgQn5U4d8Op8ACGHfyii/1TkRSpf3q05/QTEnaByocnuUEwz+VGDJzpCTHju3EwFp6w
s1dC65LRTSC9TvL2QslSARxgeB2d0tK7CkI5ZM2THQYMingK83opDHYQn4adQFz163mGtELcS3Tr
DhpJ+pWRu1eStBYVlYYwg1oqh/g7hit+MxybnfW6pxe6mrnt8A6OwB1ijZtFcSDmUh7ckNFfnHr4
XwHmScWhRczCFjp42mshAKJcJKo6u8tkrDnum1SmTYbt3mXU9zWiiQGNc/M8ieOiFkbwlwlq0Bv3
RfeE6ELW/uY/B5erZhMWH+QJBxNzUeqlvtR8Tz5qWZl7yvWDtYmaXu58aYVMB9xLa53cVYPdogjZ
nlMTbfgV2x1LZk+CubEPq7jA8sd1XzSk8uikkwT5eBA4BBJ+0dRjItZsy+VK3gg+vDi3gm+XP/8Y
mohc0i2dmbHJjWMs8vonfH7RegBW5fek56HRgwyVYB0f9hbuus2vAx8s4NGHiOaq68ewqRGKTjql
tKmCDj7mOULcwqPiO9tVOUu6xgOVXvrDwRqAAa/eY0vqAMRkGR8NPxR5c0sQMDgqf/evNDz8vgOh
MAY8nkWhz8RgkbS6vxdzlJ6Itq9HQFyznIhN1/fbt9iiUG18T82VSaDAkIJjjP9p3W9i6m21oW1i
5JAzbB7xuN2cjHzjx6ZOXrB40z0tX0FEJnOs63i06egyo4Fsk6itahDolyk/auVVnpQsjZKa62ej
CZN5FCxHvnA+4diK/1ycRrpBpXEuPWwYRRFzCG3KejsfcjkMdry/M6/bQIaVJa19oGBSsl6AJmfC
NVXps5raEl5aZi+aIacODbqL68fBLc/jaLT8SpvRqDuu3AuyEsN3PJbcSsON0nA+rKO2uIi8A3BY
f1SvBQwYa+wm5BplSklgWpBaxm4CUee8vI9WHabEy4SL8+FxrUEeKE14Q+1+EepXgBwve8O+LLjJ
vLNK92RPnvnbBSNK6Nz04wHfFrSn5tDx/CbTLCwshXzr+7g7APqyi49PJ3yZVdNZ4Mo/EDhVX7A/
Rht9rh5fsjxXgnTZWcb9Z3cEhpAbFanX/zpIaE0Ys8rwhrALCKxukYJ6SSkWDVIxDcQUr18FX2MA
9eBuiveFPZ+nU0e8BGne8Xl5tq6rvFUt5gcv2EHfWXqIgl8ODBOrWOXNdBqs3r0itC6EMAVOE+JB
oNwEMSqCmesmpYdn+5+WD8hV1WmlbVkHzv/zoc2EUXarnCnbzmac0jxTY+es+YX8DkRDTyxcMxJG
T2/yxdX5vD5In2SyK11IJc2sLMKA+vuAVUKTNEmGqCY/Y0btzS0mby8sDvrZCCY9KJeZquMgoBDq
aH+stPHqzTU2/YkkKUsspF4lTO86TLTaJ4dTh/KvpTcr6C8qY0xAQLHPny72BP1F1ksWILBYo3iN
iz1SgZ4dVFQYpNRBYSD/XbLqNdKAmAlkMIT54et/cgK2NMssE7m2hYDXOjS3VIJzyVdvuwZ8ZvX9
Rfg1jFocDK2/D6rNRKfrEKURboEl2PtEERcS9m3hHJ7KzxPdyEPYb45q3psoqLrkVcForbTAWMX4
h/+128QwdCQuWf8ySHtqqV6NY9a6pR8+cnPBVxO9mWoklR9jcp/+Ijf1EDjaiqRO+76EZjdJ1zBx
oOpX2FfeUgy8vtWWfrjiLiZm8AXoZwdjToGz3vNSTZsdKP+/4BiG1pU5X+Jjv3SLPMbaxBg8vI85
rqdYN856F9DsMakP4BYVAP6uYBo8yhCKJc+cPXElLwvlobYAis6QT3P4kLYWzL9l/pZnxUgnetK/
hiH6XuZYkG2OYoF3ls+gdUUr1lbsVbxx4kuNpT4NnQ00qgYVzOyr8P8Awvqjh70CTW4drcUY7sD6
6fXqGJLWvjzWaTJJ+wmqoSywBtKt3gPpl/EylLxeIdFpYjZNM/XhEf40RM3JWsGBrHldAjZkMCsv
lAJd1nAUUqZAS4PI4aGQ/WS1ZfMsJ3k+wxaZ8mDFeoXtyHsTyeO6RpCBbsGn37STGWLH8VKWQ88J
yt/qS4jZDLtJXvi9q15QgNca6RFLHEw76FzgfR1vxdOy5ExkcHAnaBwBCkggPWmpxzhtOAFwU3ew
7X++xcsRp0/svSr6NZGEH6j0wIHeCm+3Sj7ovAqUzco89P0rL5k2tmRS8kBumualZcYDshgGDCmA
pGojK9YTfsvfKlV/bp3/T3p0mXbmLd6wqAZ4T/z7GWlFF8a8CE7/uvA/mMKmqDrzya7xkeZlCxf2
AIYqQSqe+CJnoaJGdWlCicoVtVXOjIGPR97vVjPJikgN0MUS7SDd+46Iv/gMzX0FkhinI/8Y9Doh
zLFfnrmerw9gGbCxHp6Zt0D553XdkCiTLoZHuGGFv2y1wDqwAoDfhIO5KKbJmRQ0ECECMuo51VCP
+c//2+AbKYCtGxChrQmr8Nf9ZwuBgkiEHlsNQaKaz344mGDB5jb2REdV6jFUknn8/Ftjh15/+5SN
yIGedurg0gpM2lcWuH/Pm+7sTRLk8NXQsHzyKOIZdvVBZ5gk1+zDPJyVjPH5D7+Ll4QkSMxUcMlY
+vgEJ8yWlI0St6SP0LSNW7+x6jHYY0o7a5SYf/SwAjDJaATJEwyKf5nuykAtsWP35Z0jt1h1ljT2
+/ctFUw4J9iIk4UOkOE17K5QXhq2hesS9pyIXp8EefOM9iEKnQHXfG6Egyz+qpKQaGAFHb9DuNr+
iIYauWizx9mDJomdBTraB1VTJhRt/Z5jFn2pNt9sl6h+Vul487EyScl4VjmCyjXQxNlhWg8MmHaE
EZnphxJ5A0NSm/kRJTGHcgrNFVNZ50J8/3VEKJdYcFLV36RqTqRwWV1eyy77P9qoNa4bJblWk26R
K8qHeoWqcSM28Uabc5YS49CtPvuxneeHV/sf78457SnvYg1CGUDtnFbUzt0CI9rF1G1ClW4qIg1Q
RurFf68iqOvvtvDK53cGWGIMznfk+OEXXqQAV/h0Ir/smM2keoiuLgEsOjE9m6JnNhdjEB8mXW0f
qd9VwTD8OnRH8ST5mNOjBVRqjclwsttfv/hPRO4p63FqnnAVfp4IJmZ1hQpClwQYr2QUibjHIgE6
PY/TSgr0ZSFvx2b4LQIeaMFVOgnFeEyoCPn0755LhIPiFmhcaU3yQ3Js3zZkUEz6HG/MXjXKcl12
PZzpffXoI5hv9UR7uKbMRiGeierq0JtBN+cDxSsn5JyyOulMBH2eiu2Yy89EzcVRsnEC4sBhQFeb
+9ygEJzajxToXLOUlbAnvFWU7CGvROWP3qQxDGf5HA1Y5FRARiLokP4+XCpGN2HRZnvWgcw+fUVM
xDeUE8QVeBbkdP5YpTXLN0O4dmhQIOCf+UTdZ1iDkgg/s4w5Mdt0sqaAFfAhrAaCly4pIYEFUlkk
7copCsgfXVNKi7gMr4T1q1Ig4kUEjR925/2JHrNXARK7XkZAc7hLjFXadtHEDnZXHunSI4cg6VLH
N3ot50mhiCculVSe4sQNfIF/C9AQDnMa2Q1Xx5/bWdZCoIrx5gOCgF5DnBKwmx3bYC+AA81hWPvt
/wmkqblswuS3CdUWWuNpuMIV10zUIqjmVElUGBXkHXBQDKUGW1CStBdC28SyxAZqW3TiF9kWBrlO
z8pKusA4mA4k6V2pnLJcJ0A7NrnvcjKhUuqm8p1qC6ypDtWQ9jhHoq6ImYgVdYXpdTzZz/Jg48LF
yqHk+DnLjVYGp6Kp4blWgxHYF451onccr1nH4L8qmsYwZznBOFd/wWRBvR1vpiIT8mACbTWVSjLp
8GkGmLl2tvAb/M9xLm5+sheEokJgTrHZnxa4MQrSoN+Bnc1EqcJzhoNEvRQXLtTxGE6wTxLU+aBJ
J29tT9wtNYWwCKVBZxPndBn+GThpU43lCX9V6eUsHLKejSxvwo/hrGgNcahwyrqxQ3Py7VquLJP4
15KMz4yc3WEItSm1j6mWa4Jblftddto2RmxM1gnkXBCgW17iyT3MIskkU4exBfrVpee5gf99eoxc
PzB9ikPdy2rvN7wG6RNBkdSYQEqvnif/GPDtQl4VUYn7Hu4wQcJO2PpdMPwUPrHA5QGu40qND9Rm
s/124PGaEK6dV/lFzifwmUiSGR5BjP8EEpltJaH7Czy44+k3d3k8hXxjW/jhyPIGTcpv/t2Eas88
YEEhSNS1yWzNvUxjfQfW/XFXHV8K4wf/L8Bs7cXLzYiYCTyr5NDm2/JEJN1MbRNRxZpiCFsgACQ1
8C1Ce6ql/VY3gtts2LqQ9m68Qo8VO4r+AzdXem5a8vi+EBJYL1DIQOP5hthqF0zt11SqLqqsHxJo
nbvAY+l9ir2zxKp9H6cE3nFarNk74kc5NNItmVKPlXyMHWaDYxQk1dTE0dXilLZUixObQB1iphXu
KXf3QYDFSsmQq5qR0r4Dgt/UM2EzqvR5sHvSsUaB1DhMp7BhBxpbAmFLtE26IAXHI5Y/fxF5u42C
WBH1xVXUO2mkijtEIXRgSfsSba1xTHYyXGFl9xqxC+cDTyEAI4+wVtwsRqJ4eJXora2doH9b1jo7
5WqmvgIcm26P6axAAj8X9lsZYPbBaweEZi41U6vnNrHS6TNbUX1qzGI3qeNSAa5k64l4yELArm1u
qF/fyFJkNjgXytqr4U507ODdF5z5tDV5l3WfO4dar5qJ9Y9Nq1b4lG8U4eL6JFpUT+ah7fk3pG32
Kft+6Ss9Vhc9/iGb2SOM7Xt49yDGF4TqNhrCO5FzAT8AVVNRSte1BYJZCMhZw5waqCVtexbbQe2+
gxNknDBprTH8KnlYQIF8/soW9lSufR5EHUIRsI8hkQh/dLI2vDnh5cRfg8UvxFQ9YHozTCB8wc5H
8CtszZTOndKes1QEEihB7KPaovti7tk9y+9saA8MXi+ch6S0bpni3zKoT8tFckYyFgIrURPW82RW
B5fVY4mCSz+bsnZ/P/5MG2pc24TJCyOgABFJYfbA9LCvIiC6IlKgczSiiKhVGmkYwle4bhcO9TSj
CfPTl15cONB7qjGS5lRCYLXSbb1Q3YhdNdywJckzHUQqXys4LhNmPylrvqa8eS61ErA3/AHF5uFs
oGQIZI7wBGU7KOhWNJ4vf8RLO2tRvFsoBqY6b7pRh51kcZ9tWdzq9mITnmuJSzNVdc42D/ddWtMK
Nswo9CKESZ2G65JpZD1sxIb1qbV3cbTAP9y5tDP1FV50kcygPQ8k904VnoN01FCSEAScN3rQCs+X
Vfmx3IgEzIGFWVAo2vuXhB9LoKxvKnZwaUO7I58IV6Pu233gB7GVA5hrQjkovGMu3ETEHWI/pQ1x
r8jf/cljU6af2KTtvXq42SnaBiro4HlfArb4etD3QI2TfCjyMaa37ilLpDcjdnIZoLuXzm9UoiKz
C+nGdnJeGYd2+HWdCfWhd35cwkrCkSV1K/s5+QPeZDyi8fdqNieQp+OWBx9JddlSA9saLWalxv/1
glCAMHEntm5b7+b3JADU6mlS9eOnO5QNtOklBMd1jCBS+XOEVaeWTZDtv1/5muAXwnhAsivEaeeJ
2Jh3vH0QgH5b7zBbOfa5VXsU6GN0D62z2GDTIw9NvHEpAtngLq4pjbIfflcYNElDxSiirzGHncGd
O7L7NUBSlzCSnaH0xAWLVESPDMNf2Vghn6l2UZws3LNeZcc8qKhvrz4S2+OGWGkb57zKIgJ4VqeJ
v1qtvp7nodThl0t0v1CpAXbbJVPyyCIu7tCdd7PO9DzCyzSXtqU+T4puHw3xbRN4eIAiDIeuWfy4
5BQDPJeMxMvTTfG6tH7gaj10CRy8LBcewMwrEeNyT1w8C2BCQP4AjjBg9MTvBsFlGydaLVa7Rt49
wfjPGbzSG22mH2cHY/Wd6yamvmNrKPWQQAWZbSqOoy6cabPp//uOY4CRmW95jLAFGKuMRKOyAqHB
yeyDvle3stPdYyKI+E++U1Q72+Elvl8k4G24T7MStRhAe0UI5nGRcOEjITInEc/jJZXti+JAVJq+
jRtlmBloZRGaDYb3F0OjwzqvcbpsVPL9rYiMqkLJnYjai/yB7tBirJM1/aedb7qsymnnxIlpnqdC
twd2Tqsqp80b6XBbNMlEr8kD2F/taJNIkuds2z8tVbp8mKlVCJTp4n99aWL5GSx1hXjuTKz6N/es
lWK1KPKDOe5F5DL++kBfcYdQ25E1ilv1DoOIGUL57+afOO7qR1T4o87LYQkrszuppF90fw2wKslA
johQ0LxKoOM7Oj6Z9n9VBDvGa01XcWW7qhj8vSa+eJwpDSY/F01vlPktygROgyepugsNjmUIJ9rc
Y3mdA44j5t7lEVJ3+d1mtu5JmAaD9LF/+Ig6RHzMX3v2SvkbGHLlZ0QwNldIqdI4Q7byX8Q2DW01
sWLY5H2zwTddyrx/X6s5StYbCbu+qj0xW/gWZuklKRZM6AOU68OIybm18dW09KpEAZ6ybZqcZ/9+
fMlQ0PO1GVOscKkQzO8A3OJ9TSCyT3mm8rtrneEoYpwoxLONAkmxS4DzOf2gWNvrfBxT/wGRAfSF
033NtP51yBlZHdCLjw9rzlyWArPKVhKJFuDTOf5c1vdq/TzDbk8QEAzmf1t8rZIMYPbhiRZyYNyG
AX/aElfWqwnjaAorPVwXt+JO5Ay6C7jXpj2IpvV7ZUcOGZeUhyAxU5XKycMhnioy6bHYp20cmK/p
8JSzLduQQwQyGgT79xC+FgBOXII9ULXwasqf1YlTxrA8GBHWE8I1rIRNqcf8vXQZtoTG5gLLmgtx
yPyJNokUng+3PSmc8XLCFX5UL9CwrLUvfqp1mOW1rFBfsaRAeoRQDXKsBiCuHde2fScvwDWuCIH+
l52j9GVY/Ha2Atc9xE4UWvs5nSMbidy0x5fRe9TZIhR8KVH1sSy84J0rNvEFlTRaUSQJaNcAWOP/
LCDbwTlQqpXXfuD71yl4qMC1KLPhJDarS79jxa9xFfXiKA+ba9i/9yn6n8TwSdUfV7UadKokfysc
S0DZhddnXl58B8TWNY+gMwVLBr11iehyUYf4tDQ4W9J0RDQpzYetxYkeVSbbJEBK0iqNTgBgW/K5
mkB0/AgnOFipkFZI7g5b53uVk2Q/DM/xCDP2CqNoBnov3yLsK/jJjunuThN+uvnE4YTEuP4SdU7X
ySkRv6oApxI0cbrqmtMdXex+7rJGYIv6d691kZ9h9VfO7eNw7Vl5s8TE94YmDsoXaqbKZ4sk+RI3
gP+nDkiBYTTP+IWs7XDyPt1TA3pAtvVDYA0UVIX1XNllOrGi7u9i6t+nq90tz0Og1O7Do9FvX1ds
bvtM6KVWJK9orRC6z0OuUrtTaQAPY6qZ/rEkAvCHILal1b1PgKki8m7sdYUN0zkQjUuz0D48Ey1o
ungPTb8/23pPV7WfQtyzcR5xELjdHsSVvuNEhSAjHCSbkRzPnjLHsOJvF4AQ5feLIy85l8DGGt7X
7g1zPj7OTPZzk006YkvJXbLnuXGlxjNK8hZWF22tia8tzNiCpWf6ueilYxbTHk5bRpO1pAtw54TJ
k6YUH5cj0fRTPTyMgko9/AaqibvxW0dwGz2e7ID95u64i2Lq8EU+e95Y87IOANk+OW1u5GyRLx1C
6fosF0yKHr+34hKgmXgWoMXz12v2q1oL2NmWEmbf7/egO993qLuIPI8a/eM6UwrEOI+u3ejiiSll
zqAXCgcSco/6HfWeVo21J+dT4pxeXrKUUrjLOrFx6b4uHqbWb4oFVhbBW9YdvZkqYfWKjKZxEB9q
6P3g1PTF24lyHy9zMkF/IcBzzHcAcvUPwbYYiBuDAKUsAPPp/Xe2LNr5OGDLvztAehO+s0UdP/LY
2ht15qDWwkEex1VmMINHcqCjE/uK+tJVe4FZFlK5sHcGB7dlhPKaLi2zob5BiSyVimJlG0M6ppqL
X7bkVewWPZlJiFFVtixzGpP6Fd1AR0hag4h4Co0Ua4UDT42OKkbbeF1ySv5348FAmDs1OFIG/41I
lWOhqqhc2NGh7XMMF56KcLDT+UphBBn5rCATAP/mZ8m6pOFAqtkHN0CCqMy6ODKy5A7LeymMIgP1
8PBLPaXHKQHK0DA9PjuP+4f6155FuhwfL0FuIsGIMjne57vQy2Yu5OpJyc0lW90CN8jdBWDC/HPK
mXCWZ3fBftyLC/qo1X+Vg1/2FqXcha62W3GR+SG2YY0G7M+LmU4WqEoO9eyzib9H9C2m4R5pxku4
Oyuslj5BnuxhgW70LcbHUO9To/ZM4yN7yIFRNH9v33/NHaaALBQqiYd0tVvSCn723ShU2gopQ3VF
QA6nYoXQoQBerelR7zGmh8qFQSRCSSwTw/3xY9lMQJxAUm0C/qaTpOSyJrD5tdngFKSpJuEtXdGz
UHUfa2BjIyF4JADTvGHoNH42HFMjXQAWymqCd3efb6myTCi+1fPd0yW+YRq4lO6eFVr/lpX6lw+z
2aujABwNh5x4ZGdtmF2Wg8/pWX/d59q+qUjYnHky+M4OiNZlqzM88ykGoDUY1hXXXvMghC/fcUDh
2eHfr3zMOfk6+PrfgpzE2hfS0RwLP765idEk+Pifsf5xbGoF4nXrTTKLB2/fApFyI4rAQhY9gRYA
Ja2alQBIExYXNSPeGs7lcfA8HdOPB1aca+JBnUeeM6Hh9JlfjeLbjRVweKYhpvKg1OYL1XJrEKZ/
JataDtEYhTqCBXWgZtogBcUe2AdlpTdnzf9QjVpLtWQXveHoWbygHZ5rbh7P8WqpGktkCZNMlJyg
432ryiLHKQtliLm/g/0PqZbjrRvwuCIwT/UZrElJsJuAfA5jUmqcJxvza+Bddm2zuRgaBYn1k0Ii
IEkfH8KJajSSaQM9NH9RE48iAdIBuJ4Costc7lqIXuzJNEc4+OXlUSFrSb5j2WyPTyDcnoa2PQqb
nn/azPXEXZ92yINqWLQIk+kvUANyUzMMcy2iM7VA8mrvIRjQZVNd/NDFQdWA24I2J1XyHS1OV0vh
UoFvE9zTl5w/D93RaTL4AWI7efijnab2LgLuNpbwFsNPMWlbhZ5xPOMw4KtZd0Jzpo3AwWr3v7VO
dapwNEYqutkXvy7TvkxCdiGGfy9U11WY8bppwOnjWdbhpMOpO28tI3x+9MmMwxg4480D+K9nrzPn
Kt4enFGoQ4/ez8TXRva8PhZeTlD6TKlkvUkB/d9J0ZHqoCjasc+qPOquFh9yKy5RvyTwa532Kq8e
fmE9XIMVAlK5FX6al0U0a4vJrN6rjbJcT7lohpdKe8JOhB0jKQIoQcwWy0zF9BcDwdZj5LdvtBRH
6h/gfxyNaD9CY6OHN6SaKHheQXapOYSz+WGv8/zwT/9M141RS2yN9NLH4Y72LvUU7B24OPEgOeXg
Mr5I2KqUA/sS+oZ9CwQ0t1pWlvmc206fJ3BZfBz0siX+dlGLfv0Irkl4ATJQNlzY30I/BS2qpd3T
A8LWiG+tALTSKVwCtwCNk/93aC+PzS/as7aEXej6tYFZmPHgXn5uKP9te+2+o7I9psxYvTopDr+K
1udiq22PAc2AkYObdeBiNxpyraVRJoAMmuWZIFlMarNxwRC8x73CcOYgoKAflaVymsfZj9Nrioqu
/5D+ZZKjg88hd+dQ5Cdy+YmduEVJpr6esPNKvHyki5rFFu8YJ4xiL/rJO4TXiH5IgqIkUnMG6+XZ
Y7hsQX49/gRDTNZPl0wOj7LQXTAAzAig25Nka/UFrPo5jZE2IaXVLfzMSAKyqVAlEt96C28qvgz9
kWElpppZ7OZwXNp5GmRh6+ouo3I+dzGg6Wc4x1njws5AFb4847BdHGjoDuHAlGPCEn9PedbLyDmG
iEaW9KGGxeSG1sZUx62acl4aFpituCMmbXxxOqt1DVctf/tmSGsgcabCABF+0r0wefbGmBjKqdY0
urTz+1eAWjWSCYklw/UJwsA5NPPThd5I06SaSzcIdDvtHD9FepXBQOf6GNOPj4UFm0yvvWVz5bdl
mwZIfroUy+Wd9GvniWTM0Poxu5HGlvDHAnNa80cocVKUClEE8erVONIh5Yjd/q+8PCuT2aqN1ftc
m1QDgY+ZdWZq4BZfmMe7twM6p6mao7E2L2lCSAsjnxV3X1t2bzyfbRl98h/vMOtMrppHZPkwMu1X
w0ovAeLylCBhzT55z7f98UqbPIobgT/Z6kvshbCAgBjVjUR8/yTu+oDf8E68PW8emzZMpetQ2v/V
3mfFLtHf8bO7mL4JCc5quKUQr1pKU0Lt4ovINLtEtA6RhuKlutyAgGMciNoRzZWp8yNWWcklakNh
Jm7bq0kcxOncxn7CYO1LrJ2NRTQhK8GZ/9a4U115JFDwWTOEB8+IcaOLvYXWXNnPE41vCCnAdNUL
l2zO6aTDNpfY3JnkXgX45A8uDjYpqQ0E3ITvZLYUWFtO/uLeFDWYQeXbXdWULK3xBfh5OW85+J2t
ikzDpBIJDEA2WdvRYY+H5zvMXEN41ulHDIEGoLJL0cphhTosMU84aiNPUXqGPOvENrO02wIE817y
mI+c1fLQ1Fw4z6y9Nqc1k6xoF9xgeeBf3GRIT5jP/BKpHviDhmK8b1dC+beTwPBd7FpbfzLdQTGu
2Vxg/Ywu8b5rSPjt55NSA14I/cWhlqTzNKyfzr+mbTE9UZx2Tuc9bfNBvMY702A/y7344zY2/s6C
Q1e4QmtLTX2mmzIahAcU4qZQCEZa4Qhv2P3/CKBMnpIIOu1/Xap/+yrtb2VCgZFwxoyq428LXgGa
mjohL5f0IxEwbHWrI/y2zS/csjWvl9jVGol6bLIECCyhwJObhX5dLmC+8jdpbdy5t5qEyJSUjkGT
4hVnsfknyvUL3aqHtR9L165FdN9GvlRJq5dSKfOYc+U92oQLhiSkR/KHAnlwf/OJOSI3e2+46kWY
it8OTvAbJo1ft/UZMQlA0NlO0FjhzBe3ktrJXZHpKUIRwBxoJMBrY3TK9EgpE9/LOVpM6JgS7RHa
s3hywVsPjeAwfHKv6P2C88IlstlzUC9M9Qx8sdT9r2nu2fAA2mEzRibtIaalge9ZDywRcX4n11nb
wWNz6AOJ8T8YduB2HlRgtBnvOa0PLBzJJFiT1PVXnxBccmOH3O3LawPKuSz5AsdgN3YlUBnKKQvs
5UAqfpupRbL4RdCnf2JedWU65XNwKJ1kB0NnpjjxwK84smx01CdJoeiRjGrXn7/hEmHWETEexnDD
KR+/peYo0tw4vRR9WYQebN3WS+WyBQ7uhbH7RnQuJa1/b5QTwJMiEp6YVmVV6ierg+eT4Tpsb3ep
Sj8oYWJOfqa0KU8EFhmaV6Si6iUSRbD8kJ6wb9e/JJu4Fu6wQ/GVGKaL8XC42e9l8XXgl3AIs9c9
/AYVAfeypojJyGkyUwiO8gPsQ1d91SnewgnuP20OPomIONlpFUVXW066Ta55yjKv5o5/yUEPNNWK
8rq0Dr78wa0xpNtTm87PgTiXlLxH5dAMn0QQsfspoZe2oSc6YIGMu4WT6UeCYaIZgmc+vydhV+pd
yB/qfbhNNERrgr1nxxthQELmlkfJ29uV/Jtt+fzipktREEIxSQ/8XftEpPbe/9VJRcq0WVPkp5N1
fM7LikKzGnfIK7puSE2Bzk4lM8628v4YOH6m8qduGS9jK3E85UdkZMwkI888USOLO4apzS1Jxg2J
fMoNJt9/Nk+hHjClc9saOfTK+xuMgIwGS4Om71272THd4xX1+LiH8AmYLWMC24Hha7E4ZCgBsAwT
MIFl9qYvHCT09/zn7+kehlQNY/ibLnClwVibDcqsw8Nkye9+ExhK7wSCiCsQo/64RgnODUDGnG5p
MQL2YmG01dzlTvGIbQ49yi+9zytYAkOG9uLIvQQqQQhWGbyi3IexKTdnb8cPl0mRG06fYWn1SDt9
XUVU6PzlUV1ONzCIT4O4VUoojMVDIjCdoR99oTMLiigZM3kAYh3leDr3t8sShJojgrlnc2AwInEl
wQh5yibCN09vmlbYLjpsxa/lIQYssIvKGkYhhJGw2uUZASUQ4jvjSeRsesMrRbvM0zeUTWBg7UvH
+d3EcXInVVSbW55I+1FsySTlbRpRqoAlf9njuan3xSFIcRLYWO7zVJWAa5EsQlYkFLbhz26rnhQd
fPyJT/0RbiYg8LFxekdUyus5SosFjqGkvZ2AV9AXPS9heDcPiswby+IkLglK1vcq9/6pyR6NDr0G
+dXZgoGM7oFqyQNeVL1hSUR78ld72ikaRDZU36R7KzoThFl6bvwPJNYMmr7KpXICLcSFk+cfZgQ8
pyRFLIj/IP95TPrhklgNIrDd99UBRBcIg8jhBL3RJk6Ro4iaotviSkF/Jgv5FZxhXCvpgr6jLHhm
ujEVeuMBrki/w7Gz03Zm51DHXeiyfK6T1GbLYyYUX6axLOgZgUK/RVrow+XhUoXynFzNMgej2Kx3
BNPll0vAKyJJc/gDBknxw9pdprc3w9/q+Va2jpQK09Iw1i4i23UN2KNgq89VGJMkAi7vEy/CqFK1
CdRSMtdYZrT/ZRTsYcyHSs/ShabXw1dB9M3JtSUH/jaYq/schP1vyjNgwPjre+5t6FMBYEMgPgrE
d7e7WGxNjohT3XHaGcO8V807z44nvzVJ3RdzCm7Hu8F8OWM8aAGVFA+3ARFuX2iPcWTxnIbiLLU8
KzqUybntTE3n9k6tNhngNicuqPqvpQECksWBPmc4dGZPMvCp7L+o8HVd2mdRkKRgcC2B7CRyWYOO
PqfCRs95vvHLemaCJ10yXz6HX9KSoqD6AEbNZb5XFCGAp10NV90CTDUnbCc23GH2HRWdGhq1DfUS
oQCNJPvHpXeL50S9QnMe1WqpwV/DHYO8lURmMI+qRkOX2m63Wwq75749tMI2JwMT5hiyFmoVL+pA
0BjOJpd0nMl8udN6mahaYterTNX/6DnVxgvnk3AMr/XmfNwhQYhrBLiedmsIgCWOIXONagUBoYgv
ZeKpOErZX6kTmM/7UBCJYgXRdV7oOvV/10BCawWToKzEp7YCkB4m6vlUnwGwI2LnYJKE3gyXtTyE
TR9aVNu5IWPN1en4yBBS1kKPy6LA/by7kO11uN6ta5KeAiVsS9+KoCMEr2bD9Hafm38C1RGWzsNr
+gZGXG42yOEJfJ1d8GQIAo2RxqzjJD+gI6EIA+EI7tzDltrR8jO9YilXnVjkd8uIzEVWlk3wrZ5f
aIixl/N0uoabEj9YTQDrgwrIRyMplR6dmsDEug29agzGsUa6FNkYpbCdbUa1oFcMNd73nKybHlip
qxe9goOlDMpF75bqHALyV4Ko/ub3m9oOJGIAjfwEhEsOiQXfbGtxoRt49ZD2peaA/KDUJ1T1rx/2
ZuIxMmg9i8PI0ruEYXy3H53jJHmhOnT8nvJ27yyrOZcSHfROyYxi7j88W0IoDL47YmiOIKgF60Wv
VHEI4Vb5pmIeVPw2eeOqETFjAzA6Xki3tUZMXdetq4OCcn2IEqhakp2tde9bfQoIya7FqO5tQX+x
OoZQ/G/RQguLQCPKdOajU9Na0XsCx4gnU7Vs9kpbl9OKxbcb44mTOH9GHRF8ZJ/dsy0VIn1Mdibu
Uzz6wSGWOhUnNIlhM3tP/7y+KAOjaTwsWs7zH5SffCrLWVDxS4xqqJxdLjA9zfJSByGNfiDXROCG
LawxXTD43b99dHV0L0OnjDECV7t3ycLPalgU4CaMSDxB6Ep1hBKkEWjftFKpAmQ8l9ldpKdN/tSd
Cq5PWCNPgkFSlk5T5zxWSF/EbfB1GCv3QhCaDDzozDAI8l3gA70DmB1XG1ERyVSByL5mYJy9zAjW
VyUWOerLNC8SWIfQ60opoOx4/NCJza0B5jDHYU5XzTQfE7axQfeUp8r45OF+1O0BpdOuHIEaO7C9
/lNenn+ddSmpr84vOpnFE9V3hXqzOmINFbP/JG1f6+0U843WtS1RsbIjcwrKVNJC94SlokjsXqSD
Am9tmy3N7UK0ECpa/B2hGqtoEdMrxaGKsOSp6ZEeFz0guhgawlsgjS0IbrldQ581Hr1v5nTMmtd+
T6KgIny4npFzKXYkz6RvqqyR4d2STp8e6qJKkGYI76L0XZeQeQ6Z8zFJNRMY7o25/NcXHAtJa0tM
bQ/xQONWI13QcuRc5WT5WMyHcBWU3CXKWQ3EUmUYp1MvG/2eyhSJrLokoKzQxgK6XITIHxC90eSo
LDgWdtXFF6A6W3zVF8vta8Vf1+SSN0HLu5asH1hl4/WN1/EHDUdQCJRngqe6cxjG+BiO/br/tAfB
i1H0P3JTaCMMVXyxpHsMEoBW9U+xrGU+ZF7qjHjUEK+9/oLq8TR86OlUmQq0pXZVxUrYLy3/+KQZ
VT5M38B7mefG8kjpwqRu8w3CapVY/IdpBLrhu+CqyK8mwU2fxqbWy0O7rCuOHPXzaUPum1+iqbp6
suHnB34/mY50smhXEdD2J6eDOViC+tSQaCZ2eFyRWmBkoBzmIWioBPjGpIJkjRq++7BenJ131dNd
6YKz65JRl7ls5FCKxtLAF9ueZIkTdz9Kh63O5JAlC9KDfjJfFKwkpwCQz40yBsLt0jziJ1B3kWKd
akb9AcdbYiXHP4rN8yoPmbcHExm7BEvc9PM1UDM9i/TrX8iNd9PHW/VRGGHCemNYB+ZS3VhugvVz
r+qOy/qLFnfHPRzgOQyEzqgXVHtrJtgTGgJE8tPPkm9XYSPJeFJyfKl/z/+Ek5YXWBofUOI618d+
ly6iwCFNEvYAONr45JUlEj2sfhX2noGm4g8E7BBTPP5lm9Myy0rGooU9y2SoXECJnDwHMjIJAURW
B+o78MjpzvTb8QZAun6bJLWbOHs/rwrBxfyLaf4x6c0K4JguOOdLAyczWAo6COux6UqvDJTC6e43
5oZBjXZGQiuD722Ah2H1u9EQz+bw40QMFV1gI4lKzK1yH/PhjHPJyBTXb0jeTjAQqoHUN0VZHi6l
fErHPK9UhydlyJPH16pz5xFmwdimTo8ZJZJN0aVHBnOlfjcv4K8d7sVgevTRW0sTDbNXsZpYZioQ
T3PDjl2Zsdb27E0/aryka48MRZ57BXUn3pn0Hd3qlQBK3RtrlSci4ZiCFLxiLi1ab8rSCCvNiPEj
2Z1BJl/HPEpl2h9SLDdnlV6mb4SZXC+E6p+7pt3GGoyYp5z6JIhAYDJOy4sfDfzxutiFaCSEzRCK
2ooBYb6A0HBwj+faRgugYE1FuGxDh6+pQ9PfaokO7T5Qyy4gdjM1mlOWUuUK8Fx+lGyO+0x4Xa1F
4t3y0l/oAG5NcPU/JLj3xoRNFtNd2u+54WNDkUkWCzN24RwcTVwk804tG9PxZ03lOTrojrrSk/AK
Y/0JS1OGEW6+o9Vk6ZmhNhwfe32iXJoT5qQnah3OoX87KNHuPkp6k+K+Fnm8ctaZYMFXcItfA96D
8pnp49AjDvRK1gyP3+IWIPyEQMFqDWYRn1nVU7SKIQKxbqt5PKAMzIcxoAIhCWffqATCEDsLn3Mu
PZWekTxPVxsBkdtayeSlGV4T+GHu/GnjKIkD9oPsr13Mcb/O8aTOe+dQzvEXJJz3E4DD7h3sLNqW
zS3jfvlEF2cwh67lwA2CstOE09xh0tqadrQI8zWcwD+Ox/i9U5G+jr7FbNG3ZIEN4rmBNSiDjCuX
Zk6UtnOBTFxnz3fmTUjy/ajj0hAnMqqVQIMsBsuMPLIBuUHk6OMM4N6fn7LyBaexT+JwURO4wehh
ZiZTwN9xjAebM2X+hXdqWiCeAdcIFE1av7c9Sv/Vsz6ODuc9a+/YS2+tBY9f5u//m0Igb0mLeEat
RnXn6G9WKYgT2th3jgFxn+u4azBkb7+vGqQzWuU56qsBrg5jX0nIusV3xPY4skm7Qah+dXy5eO2J
LWrAP0letP1bss56Xs5doQd2cIKsBtxeEvsuCSyJvdjhmu11elndZiI+yIfda6pvOg7Yx9pC8K7J
P1y81YYUthtCNAJ3sr0Wr/3kfTyuu5mxOR6xOPUaQHeKxmCioqJrZ5hMN2Rmszdc7uiFvz60IssI
Jv4KOz70tOGjbXj6i5R5c0Uu2XtGUdpSrfoXswK5PEBVXSnrXeHgoF4D2ae80IKK7p3sEvuUkk/U
H+lS6/JaY53L5TSfUTWFUpDy4cP/jbA7JwBtOMRic3v9/CpjhI838z4/YxvdHytMt5azYu/hfTfE
Fy4yu+K/MlN7VsAYayZGR/7QpqGrugiaMKGzNrCHATqS5yKxA9JNHX+zrH/xmAIikrR+dYW2lvEB
NY+foiV3dqQ32D/XAKg6uQlvdK0wgSWIwtCOXjU8fcXPMkcvpORMgGLiWtBnUnozI23f/+zhEKcS
cit1N0XRjgOPLw8DggJmC0Jeb/C5n2/QO6DnayQwQ7KE2lfHM0n6Q190qlKp7fI/CPECv32TsRj0
3yjgOgWl7UHsYqYrEEeTbZtD+G5+aS6eANURNk5ENOtZh96E3Fs4yDuU6P30n1cvCvRH3fC2g/yX
gTz5hN386NVEDvH1nJ7/DBrOODwNDmGSwyMiPlXknXgfZRa13xNTGhScT/MquocpCmuWM1CfZHqi
NODaJUHK/oStG9xYJLahEjPu0ayO4xUQ2oq3tJy+9wDKsNFP12BC8AsoN3EKSQKt6KWZNNyW1pBe
OL9rgSG1Oe90KOyHFuGgTL6T8QfgdTQGeOzl0LvQv9XLJLNkKhtejlIM/ZV96fXqHi88fGBx+hLs
e0T9ChRpBNeaNjFDlJuOw8j3UL5OdydaaX/JMAuQD8g4DZ4MOMAs015v05qlskNBStTGaZWMzTej
rZPJ3oP7Q99pEKkyMXhu6UMH6rLcU9zlB2KpE/l+Oti34752lzKY1w+T1A5O3Y6ZjUqhR8+nVVLE
CxXk1/OXzczHw5YdwQHYF+FPDr/QuTY8TOlu7p9Ex29JsIdniZFMNe19AHU7z9XqwSmoBpheKU4v
OVuGDvH9jGgzfWYO/Mse5Y2M6uBrBbvQ+Sww2tx2lP2kO2VSpFRRd+6vACU0bC7PavXJd2of91yU
ijES7ABc4DLAH9n27iai+siMrsZHlUHF5xRvFb7PRp+u5PhfBoBR+yoRHANPmqJVvcx9GRnkfOFS
4jFhc0lQD4F8ry+H1yNteaWKt6McdwuC+ik68AgmMayLSxM4kV14wRwMPcCRHNwux898mzbtuaJ5
iJSbI8UnF+JuDrrmoEb9UBIb9fBf0JeouMFNPTUlrd11RA1w19Z3TAj9BhVFJgUv21juCZ2VLVo5
qjvt2FDnehaaQOImlZec2BfDnosc8Tnli/3nNkXxOP+pEThIHogyR3C+1KshRP6omIP1JqOPc58b
N2a+7F/phI9WlK37IstZe/UBni+jV+2WZTVcy9Y3D+dsgsfDWuaYeG7X6q07hrmARTSPlAjtH3xK
lpoTZ59dP+pAblzLrn6jC96mll6GZ+k5mUkCvPZILcG+tKMHSzE9fZOavxjQ0cQ0DvBboaqWDHP1
Sg+trh40k8ALYsqkO2xtpNUVxvzGsy1WJVIuAnl06b+A3ofBmjnkrBX7CiE+UJrIPQb+BrYA2UGI
DFDR/xRri1vKDAPFjs1G3Fg93WwIgMX9yulnh4hghllQkcZaBm+T4sfuxuSjmv02ck8RT2KXTWyN
xyI5TlCTD5JKDleIRG80COTD2Lm+ziypySyUneC52w8JWIh9zlLcQaSrhMJwf1MREiGzV1SV8YJ+
iMK+3QZ+VIN3j33ArDV2SkC9Xcc9P9fKcjpDlZg98PFc2s6dCesBaBHGc6PTa7Us/fBqYGrEzWsS
RfLLiG3JKhx2sblFCaGShyQuntoDaZ9Ir3MeLvJHTYD5Cbq4hkWLStzvpFeKMPwBToDxem7GdBNb
xHy+c+4LG0KX7+XdyRGceCjX7+G0iO+ixCRrqYUgixlSOdsXeWr9Rd/nnyxjUK5YBSSkRI/thaUL
1PkibbThG7uy834+Ja3wNDkqsurPRRnRlanamLidtr0iPSPZAre/yt0nEwSTRl8ce44nvX7Vkz48
YJrMWDYoXx1rVW03E6rsWD/mUx/p5QpFWEn96JvPZph+RtkZ5+5FWb2xNxUJ/3VrXuLPv21ECmXn
cwtNmMQ1NL9VPoQzozUKPMwrrHfjBignBMLACo3GHIMCc1tcNEcfUNozPM/SXaGAx4fF8KrRBkL1
wU32gCCCVdpiRm71Zw2XhCokTeWYfEfZwKtWVR5q5OvXo8cdNbFxzaL3N05c4iOohg6alOIjfiag
lIWXczY5DdPyp/ILEP2I/bqGm0DeT3vAKJnEBKygSZCVwKalMPitJC49heUUqGb+eckk9sjzgCJ9
LT5DgMOjaSEPwq4Tjsnqi898HiOJ+oNpFqCkfws2akG6ZRmNsKmDjfYHEFfd4x8yv7iCKjb/cXYV
ouZnUHQci7Ko/b9rjtYj6P+yNCdigAzaHWYWOethusJvEIa8tWFmP+7p8YNgV1tGl60M+YMQbz3O
5DnkaYznjoGB2egz5KwTa8KdUeKouaK3GNJBAZLkMTrcoYZf21B3q1I2cb33J0uMqLacBa+vrcHy
C3fqdzgvaPBJpGnIHyGpIb6FBX9MKTzmcFjavNkPrDz8/mz9SZBi4etmlr2xFi1FQEGEGPSD/PVt
vRfRWJrxrSYfyUeW3z74n+qESfVVdGtMH3aFX64ENZxy9O2GsErhw8ocIdr+czs2QtPRQMl+Kr/p
0BcY146x9qexgEp39MUUEK+TkunSEfnirrfKzoagipFhBlhlP8arZCG8pNtK+JO9psmkSTW7/UJM
HYJeCHU2g2M9RJHJH+PcRdjwVA91EzKaIFAU5fOWPQepkpKGtshAsqybdQz6lCBVq6Z91pKTnht/
gsuRuY4TQlBoUyBwdGCJJxWqBCTMQPjuN4LRLUbvHk/YbZjoVG5zAobxpO7t+m/1BZib61T65EB3
E7yfI/V5fwC2dEI5yb9bwI42f5QlJymtvfkIOIvdT1SWTaJoYszK6Tjsz/1vUQNC4+zBlIjhF3g5
KNkbwszf4sGv7yiv7xiFmDg1H+w2OvNazzcvLb2LzsCJzL36TOS22OCf8jerzXpaxmkXQpT146e7
f1Ri/ocKxJtHrErsNg+0O+zduKpwFpP2DW5yxk6KsWtzV2BBX7P6fR2FSexxSZwRZvXxQRwtYBhx
38+m8EVnIlAPlbWBlW/Fq4Bhudn0GNiWbyCa8X1l1bGjQzGzw6cUatkJCuikqq0mfiQNw55pndtH
NStEWLHP5oqM/ERS4WeeQyiqyqZ5Y65ICPuPkEXevt5WrHbeHy4BSAmlC9HbSy4M36Zvrn8p/2Fg
r29YVMzpR3a4/jPvLiTGDuLZrCxjne9L/c0isOItp2qUmuFQeUx94ipSvQqzyb9ATStwQ5t7VfrM
C8o6UdnFC90LS+P8gtrXi7m4ApQfZE2SN6Lbgx397AOIQc6Lu7brs6KIqGvqUG7jyeHraXjBuLG9
oQTQEuXxy0dKMGO9AiBj2yBWNQcDcDI4MiAygVyKXpmNL/oGwGOWCOu6WRba0ji+Nw5cJ18ir/tr
kExKuEp4CWq4RHod9iPW6aEuV0zLI7XXWA1LKwYzaegtA67BhbQseDaBop/R7X0+B1tdLFYQ6Qjz
MkTZq+m81V2SGTbTcOtPNNI8JxMX/nd0y8ezbxLJHjSymUpbXu5g91lC/ZQa4OV6koe4H58qKPWP
RDhdvFvFwVNtPN6whJoC7Xd771muCNzBj6zMsX5P/4XibCkIRA/wMEGyFbwVNesmR1GmyBsISsa/
lY79wWCSomP9k+BjvRp+fxbz8RRc9ihV1xp03BOcM1mjLh2rwcJqtiLQVBkqhG3qOOOhmEPwY8bp
R4WRQ2uxP0ZqxsrK7f0VJ3hWFOURAHC14i759vYZAY3/RdxjQtzD/vIXBCopGcNriqK6sMZ6/2Ku
H7NjbHfJBpwF3IcIjDvFesKZAxR8zP9/s4A6G1FXcL7+MnpRFPt/gIGJy+B4FuwjSCSFenzc+cHn
nbU9K5mVPwgNM88A1G1Fahjx5Urshx0OPnvYozSq1IiU/oWmAfgKt0Hi2q+G4CDI0vzhLFqbplnK
900Ejf8aej+NMTeOBUUAO6Fwq002DzF3hdz0B+jTWfZFO00XFeCRHTF36g+qLYousVAhpGESkWgj
tBzM7VKo74TckZOHuvDls5R4VuoRJc054FekMMumyPNlT/1Mp1wxQVbQzjwOEwdjhC8jSLtrSdi3
4fj/P0UhBHjXeVeamhgXTxYjmdeGTcH6wFZvC4xtZrIQTySlMPK15kyopzzxbx1BoAT6No9eren7
+5KCuEKzQLmITm3KU7krJwp2FcZT9cHtPALJAxfT8ZJdrtDenIOdaf/alioHuGp0PJYz3XPf+zqR
X4VpQtasdedSDYmZwCXxjMx3Dc17kl2V7AgcLLUu6h5MWk80bE6YKswMioqOI1exTWkW+FXFuxk/
hRCoanb6JW/3l1IA+YyyYkIoRieTf7VK84CCy0kSZ89cI1Y7pK5CathGePqXDUPOVynRLF2sqAyC
cynMYew7Cq2ZuTg7j8Rt54nt4ZDQOKI8iCYqroCkNuTNlrMZbfL0u2t8oqZRxajz/f3QnLi73nzF
Wg5p8jnh+/FpvD31vBqUzg0lXqjRJDQK1W/EWPTCwcHLALphdOzbSefeoPVHCECJz08BAI3BjYYG
9l0SBCyHsiQnFCoQ+/q7bCryotg5zCdisWrY9z+UEAHwMASZVPSvWHptG4yYmrP6yp5bLOWn7dHx
JsVIopo+Etbor1Ie9hHmzn9jC48fOhpekI9FfcN3LGs0kkUe9WM4nMUDQ/WIBFqKLbZAtZUMEwZC
EyncccxR/PHdXEujQpt3mc/2OT67KeCZKTOlH0qMmgi7Cg+r+xQMiOHy87yV0l3k4UIWsaiqroao
BkTj5V79M25gxRey4v8ae+8fOz1oSux/igyxmROo67hMrygoCX0pDHTBdt4fQgniA+kfQ0XUPGEr
YGalnWOIIKRg1vlpXZfph+PLmBIBepMJgSzIFAeUWCinWEuOwwo7yZ9bxZtLqw6v4Fr17bnbmBlc
BUPNqRv8HcMTlzjR0CdBqdRbXDvgrDKphiAWuFp7u9Mn878jB+79zt0Z/2dWyP1jswlriMxCCIdr
zaCXKmNmbwo29YREjoUWvR+jfjEowJMvtAirXh5LpI6vlaTnCNlx5NIFDzqUAusl+UQa0ybjl6Ow
qD+neCqJJ1yMIVoLP5fMvHHt7Zl/40w7/9lwJtqYYeRIL/mZX8atXPuOiTI1AmQBDxE3Y5dGNwYO
rOjboVC3gXgIEb6tT8CBtvKZnyS3RzjGmUte1N0tUkkEnEtSihSMLlfznU0xbjPfLh3Ki/VUTG02
JzFEzlUc12wPS08C34hYgJK7LdggcTw13kbLUX6lS/2Zdflr13vE7PE708KmQ0Gy9PmqZIb1CV99
K9g4IyeG3TiS3LAzacWllS1/YZ7y67VYIx1iTfV/rkUKB0LfaFN8EF0rehKh1WAiMDk/uD7HzaGQ
8GxV6PT0D1zF8ckmIlgPEF4gqaoKFqzN3WXHGH0XjZxiIu0VxqIHJgakFy1HjjZv8eVDR254zYy2
GVeKS7gdiVLbh7F2e0cYlHuuOjDmztXuOROKHvMde5YEuyQxwpWTyfOAF13idBrZPNPL1tOeTnyQ
JYQM9JnJqVfZHsBOUnd7fgfm4pt43HHIX6+x6RXiBYZsdBuVFfmxLBJRj0TCZ5op716QlV2hKoW7
XBxVSOGxzySSsGM0A6NHm/xGI7L7vbuGJ9IO9dvzo6ZSeBdMPwFzqpbhPpa2pssDKZbGW9LrwDvw
IqGm1u2B5TYtqnzmvjURDhGGltHNJDjKHe8I0GxXMV6kivHucnpHSHSRnKPrsMJLPwT10aKUw5sF
7u0gxUX7Hjkgp1JDeIqXwRoXfJ9rcqcEZ/EjJlWjOJUiKaByMdt0jnMDts4RjAYM7OQEnN+U0JaK
2QJbbe82Mrt+C7q7aGylBp8SEcYoZck1OYc9EtbJUZRWq44wUUa87GY0t/28YoZzTwf9dnQN6dc2
fpQEHX/SGv9bjHJgU4os1/YkLc8fFdqTwmd7OrWvWRix+sW6tlAD+/RRGS7GwkSNceYtUq2mP2qE
9/ze1pPm3IUOjiVyNvPIDjTbF3aGyF80PU4eR6x5JLlZvHApCdJF+lPFI/cQiZksljLTDA8MYjVd
pBOZBV9pfX6ALCC889Jbf28pKciMq36wEgqLVWODVeGxXx0wK/z2WqcYUzrZvGy4toxEK8rcxvFf
JhI8KjksUdhtlKxv0US3tacNdtEFg0wODDCSQ4GmxzyKLNpP67NaLPLIJcegz66Y/+wtREWGfWxj
xIEgBqa9DP2ZI3sR8hBo6eKkQPc8j3vX7I7G5eEGKVkweB80EAxBwoQI7c+H33Janc239zvYHZCr
dbyd4GoKuRl5BEA0Hu59y27Y8n/AYCmG6kHnv67r84S6id2LbBy0FuYtvkyynNa3/2XSog7LdCLH
YKVbfM/s/sgiLqFyM7/aZC5VcQRWDWH5aWr/aeD8J+dmIKqgi4YwMxPoLo026J6HJNzISEZixOjv
mIGg6/Y5Ihtpg2LvCMlrZUIINmZNpDpjSjHKscvptJpNqmMQEMwq4muAoOiRwUQCWlSZyiZ9UJ6L
epgtqYIXk08GuztoA6jl9VO5bGNUsWUpgPxt+xeWSmW+eIcpgHZru/4RmNzTsRpZzh7HoKwixVPd
ekvl7G/VhQsNEyC7/W24j1AkzizONpvZLlNySMQViQSiYTrND/8jfaLX9rQFwlenqKGN+TpHQ2Ag
9I9VEeTXppa6X3XfrHAqvb81CJ8Lbs1A9gNGJn1qqEFIBKrXCiYMeo/2ZPn/njV9ECDx0YmHR1sD
wLNlClGojb0H25OKZ9ISRnW7DX5+V3+a51VHnxeYdD5U/yN1BfzwPEmXhw4v6RmXexAAtQYPhRef
dJ7H3aFNpBjIzo4rvwk6ysxhy7cPpIl+1QffAb+HguscAWzJdSzO8ZR1V+/DaPzYkXoOBqLWDiT1
Kt5/sMvNZXkM5WgMtGknoZao7Ig4lne8hCUSSkE2oci6q+lYBVTo464r4I27EtHa+ZLtFnpkQZeU
PQcY4cfEsqCeF3dNKFMAACpO6ZEZOphd8qMgaZ3++atAJz4ItIqwTRoeXdv6A+TWGIlBqBIpk3mX
tkAbNug1KYgBfPcd9ufOrKGn2CtPsE1AS6cQ0+yVGrb0tAPTt7u7vrATzHT8obPkRVdQVJMBIpeb
7yE/1I3+V8LKz/X7rYoA3zP1snBnJh/CJGkFzE4jg1iaZx6jMfwzrqTru610bZyXy5Ks+P2DqdH2
XU+0Mrpg92n7RUTfXx5DqpyRjorynNPIl/V0OzoYdEVskqBdENBXWGgmmubmUhzZp6iplhuHfZuY
ezISv2/HaHbXSboW4bTk6cCMIJOF0O2W6rAwecem++tMbakLlb1SDfM6tGhjl82795voZBJ2yahx
PFrQ/uAYvFHiFrjebwApSWpNHCeEzLlAYfqGhdSK6x4QoSksEQBmrh0uOw4wqvT34r6EArXzDRwD
56/e8EDn1lmrGVr1wK4eIw4DyijBiX2hphUO2Qc+1kdK243pJNFBrFOVq2Zk6QxX+jbkJFVTTh7o
ddpGwcpHeXA/NGhs35UM8iee/n4dL2pGzwQn4l9BFLnff+0Qxt+KqiFo2sxf8i0B5IF5VEbGVMe9
uiKnF81A9ajX6Zuxsocief3BSAAMpHbcSFlFJlYCSxaixLLGUHnIXhK0zW/HWBef9FpA4LWCa3Sy
qfcvkwdcsymAVrpNI1OzSHdBlRlJrmyvLMwhfDFKSMT6qXYQaDKy6LarirlUXH3EgDgxwTZjOY9/
mlOzp+OjCEZfgMbqRRma6sMFVZr68NcmHySUecqY7kqY2JKJECV4hI7S20AOu+vEjLJNjhDUC6ts
5mo0c1HLC2j7F49Wp27roSoMocySiGCAq4gjh3UtqHgGx+hn4fGF4bSjR56GRAFdNZHeT+EE6lu8
AZJr1Z270EWrOVsNUZR4VzgBs2FsmMIrubIyxW0lFoWsZugEWN5pmTdQzeteCx46OWwjI48NhQ/B
t/emXkvaHTQtYI++QYKtlvQ6tK5eUqB+ISS7rwN9F6Ssb1cIadhI1DwKaMZhNVmzClRPkMSHNWpC
cWn58xNNQbvPdo82aJ7GH5heSux9MMnXS/xpBAwEYqaQoLDCeaVVUs9sz2QmZf6cGVve71rmpEZt
1KVFhIQJJeVMSgF25RYVBYRhwu22YadAccigftH1JpVqlzLq8TirHGnWMYD1Q1TFkh0hYnZeIyya
01rZH8zUfaTu6AXwQOZ/cnhVzrnmFzNyw3Y+Ud2cJXsU+xK4uzYaU6w9K1mLn/v9fowstbjhy47t
7/jQLDzxiKdqRKhYJ2NGJjB4Ws8BfImrVJPbBvqkC29Ry4S1Xg76dhHKjKzHrq05Vp7zctPhjD3X
1Qgg/Zkcq0WOLIFPutzWuMH7PIhlgvgE1S6JAQaC3unJV+0HsckA8KGtQwkguf88yX+VkYgFVfUl
mlCn8Lmi3Kt9hEcdBopJfcJwGMuZkk9bAlXL4OH+2Uxp0vG2gHh1A/dQuwpiwdgh8L9WEKFHlbuN
WTWxqw+GL0vVH5wCNeoKQNRZ/rKTMe+9N2yoJNyytEgbV+OjgvE+pDnVzoTcAoAnYgMNvqSKCNhc
9pOEPnHBxWXCvIJVomiU8WMYZcCRiW5du3/8uYP1RvE1i0pZq8O74thYh5FpKyGnda/DnaPVO1pY
D0Q6wT9XjtV5qWO7LUVRqmBqs1MGaej+013YhBnnxaGPpUMTjhKGQUnpIAMoTdch3qHIkakCV7iv
CJS1uVpuk9X/Rp+3hNL3dXmi6D/UR+OVP+CRDwsyZWB8cTmm4dSxR3Ki9aOWBT9UxJvYGb+J6zpW
245NToVS/xImwMfE+p1NT3otAFYDRLPGazmu6odo0j+3i6gInke6NLn+0U6oA4+D5Oc6VtIo8N55
RQbnLuKbGAmpD41fEboiHEY2WHsjyswaDbmsZxNIjz/Z4yni5Yz7ftV4KRHF5q+2K44E1v1TA9fj
I6w9lTEj3A/Ni9VUWc6hmws+ahQZjEssEobS7Xhc8iRo7EeJ8kmTIgBemYuBfsYaMrN/R7hIbLF0
wMj6cJ3QwGNNA4HZ4ZQW05FsyCx7/LmhYbxBHi4cP40gCtiNhvTeylgCALsSLUpMce1XBhpBMU2M
QvpOVQXIsYmc7qH7eedRu9h7qoCTwhD1GEBHsGBa3LSJ1JsqC0tpe0P8KDHDYMbwLrduGiKybiTE
uVACI6aEq0/8BPsz+cQivl+cirln6AN1IvW0Vm8g96G/428la6P1eVZwHnPM41kS6h8/r9tococd
i7tKAVWkNmxhGkP2rjm58pLK9Xu/XxhL2RGuvRCTulc4sp5E8pY2cyeApEhqPp9PtHO5I6+NlTKi
jsh+AHl6J9FyWtPhtmIPANdrwmSW3FvHN90B/ZyfDzkR708Oy+T2ixtML002p+G++444IRzsBorr
JO3JoyROL0Sx26KH+aTcn2+XE2JxD8BVk/kn4YpZXWJEk0NQKC/Azk5zRId2BBP09mjVhLEImPJc
CwHomaPGAQpgSs92DBlLI6cI+sGyMrmtLbIFcAxKq5YZJj6qg0azAhlJih7Az0HCpAkM9RCM6K6e
4U1Ilvupi11beT+zWoNcUbmdAjtcT1FQssvCwmHFFlTPL1oo4b7lAoL6WPdt9wwyTGp7m7McW+Tp
Fi9nvvz8v0/TIUBSwAd8TAbGF1r2Jjmhl+ygZIc6GvEPqgdGONEhjkZvEJA0lom8xp2xgGfKahnt
0dUrGxulfyzNyrBQVkwa7m69VEaOe7p8Z2RShQAw+Z5TvxP9PADL8P4mxK086sltwVVZqhGBxHJt
W7pof0k57tLRTrZ/8vTIZi/XSPeWCLMehl6UIYy8ralihXRe6JKptV3W6W18GmrcuGkkLU2Vuh14
WNKvJCMwHv9f9aji/aoZcMIEEg+LPzeK37jsC5VpssrUbvzxdgjDbhyLcUrUaKnzkTAc3SFokTVQ
sRl8XwdT4ARC0icWoDcqGHtHaGfJ9T+plYWHnLfWy6Hg1JDnUADa7NbPjVp9uQUeyD8ieA9qWBP6
U+M38t2UPrm1G8JgjyNFrB/TSXmYEA0CgBWfYon26Dyw0lhV7N300Nohn8PWMAeemK1/IHN0UZo8
WChnctwSvbTa++ZsC4UIMgtTRKbL3eE78qfNnMkePtBUYKqrzOQ6zZDIM0sa1w/JQH43E2QHXxuc
BO6j6RZkaGkZjmVeP+2CrL8EBztAL6iZPZ034d1eskScwNPVG8Z8X1WQmf+nlk+ES1LdTzxFvoiS
XDGCN5rze3vXxmF0I5BkrqnsEkC44ViuxLzoZV4eBceB5Y6qSEoIdZmMhqxmNqW0DnM6k+JN++CN
1JIeBBAl47Jc7GRYi6F1Oa4wcRBEebEzV8Zg2zpJ9gc7Wo8aWmUGkQt7NyyTwK/SiweTc9i1RBni
xhu+uZVIXFn0ePGApT9AhF1cWXRKLdDAUMAvXYjlSQZn1chc5KcM0ppaveGFzhPyTeMewN4ZxHgS
rBBQWV1ugCBMisROo8K8YscrfkmiwOU3mJ+0yTO+/ymz8DyW7bC1rvsNwJphDf0y0ZRUK+AL00Ji
fdnmx8DBxijSvUyQo79fF+/9tfXmROTFbNs4hqT5IK8gqXRL5YvfZNZhxZY8IojjOTOs5CYu1RxO
JWWvFy1AeDS89FMn8HOBS9Z2XfPoVLf5XTBGS25MpJ30k0uyqLCjBlwRV8ewyKxLPlyBYP1abyDj
6cB2WfGStpAqCN7xnvSzhiX7Y2oKErSB2LOiEPkj90wOdzH6NYMjH94WQTrznC447IMTXlqOR9cH
4M047YCrORg5h9ZqfV9F+fo7xgm2zc8vzV2aeC9qoTXekAuEW7/rKybbjMecziXf7+n/4ZyhcM4J
nz56Ix1mOZRF9etwoCmARNkwI1t1U4eqRGQEs5vRy2DO/236mPJ0AWrL5DbK/ypgnxaRjfyIY5cr
1NKiHeOwgwR4ve3XSraKfmMi3IwcNnkx/0Ohh1UqST5dhG9okZ5uENdvqrX0Z95FJ75xHCyXqVvE
gTe+Dd0zDmSMdCe0RdqRuLaDJQImRxv1A6fhAHL611OIyYT6pJeddrvX3WMapHCrC2cragaQ9F6x
wQ2aRX6O3wLXvtDxcqm+lzwVyWdtVo94IFRb0zgOUiWGAB2lPcT9lf0t6Nsp0R9V9O9CTptsQly7
PAblQe7lczgnpnfYDo0QYUh8CTRp8kYcmmOKkCwCm1o8f8p+eoc1tvEbVQglxLqNup7rc8zry9AP
IK23UqzqvMMttjRExqiL2bRlXvSe4S+3NNHAgSJSlbPSfxResx7zs69zo9mG/OKtXIS+4n+wXLMD
DXdnaGhZtW6i9B2PIzg9DGHSi+pSWMu5V0tTpcLF/sW8Y4Pq02XzotZd+LJWwYlcW/PEXW4uPZFn
8KUY0AJsv3kscZ/figUmPO3QRRFhd3VVwPLoVOxsrIlNwmD+NTZnHmsnL2DQRMaR4VkpEuLSunuC
YuE0xoiSxtGYHxyVZLyJtGXC+2tWk/QTWx9opxpvUVueM7U66hBvTDHxoXKh5MoueOfO5i/E2Msd
vSbyJKD28htUsJ6qswnqWxW0THx0h63u/iibdlKSl2GDeGEyG9u+yOm/5a2MazOEHvnmNvAt/DlN
dSUEC8ZY5ssuQb5XJmyCKeYYeoK6B1YKK2/PVd2yoB00HxdfZmEW9dgQwiaUCVrl84EbS6vtVxfu
l1xiOJ+HqS8i1BODpqxujGeN0KpkrEerpUs77QhbZsZJIxBkO3HraZnMaNK6cfjTnLQzaIuhVlJA
eH3A7DunZjJCXXQeOPtIiMS6K/KKzv2aiWWmrH8jZtu7TrMimEkxYFvwFwi7cuvfISBoeBDWOStx
XB1bpjL5o/Ybu2GWVayiO8DK4ZLIwWkRl7ZonwYc6eK65ufUmI+AjeYJjxfDYPS6PSzokwHrxkJq
N1JSYv0tTVwGehhd0YBOb4F7fjfrCZZrQe4Z6WTSXU0a31VZ/v4wsmEvV2m636ofJZcbPcv4YJtS
lK9rWv+O9PTfNy2+SIt0McD/Rq5jITiTFGEJo6n78NG53nwRrVc8Kl0f/avAVObBRE8Mkf1237yZ
yCG1183eonbqx2n0A37lTUxfC+PD2SB/XI+u3Jab+zw/FIItjso0+3ke53CeTUMr/o9z67DIvSff
FNIE6QnqmCTMw74uGfCT3+xXIEKuZdYZrvtl9eOrxh6rVrcJfZe1FZty/e5keHp/dH7ZKKQR8SQJ
gFQmoSMlSFRqtNUCFHg4rJt9h1qyLtTW1i/+EtpSVIOv9gOeNXKZnMfsIE+ubiNCPe8Jwm4/K9wu
GzL4/tarjriLiGZNP/9+N/uY6R3fl5H7ew0WYjTJi9Seg/Qrp/zinzBe2VgIICBCI3sjvCJIHWVZ
FrIb60Xvt0VLrAVg3NsdgCekIPzZGRNJqOHfOfpa1az/e8EKCzaSliC9KunaXTrbP4BFBRxdNJWt
9NiK1jBb4MLLaIvWTNRit79/1Tky/HAtLQ9UH2DdNTB7NOJD+Vn1iUdkWhW33GVWlI5QpC98IpLl
3BfcksTO/MDrqxqA3Lew1lCMVbnzSSVLD8TZcppIhlRb8rG6/TZEo1kBP2HbFI0GDhD4gD/W0D07
HasObAzpL9L6v1+UhZujWrkRjNOwUXmO7eOdTYkugMYaPQwxfmFr8fKZdw6s3fOMmyFW7XDk9V2i
guuwe6NSGM+hFnfioeZxAcfwofLEv9aUYjXLoTtrauHvDdXZ51oRukgwkC5cb90phcIAI8/DZIAA
r9smnv0h5adBzZDRAU1WKDZSrgz9q4NipraR12iateu4WL+ERlXbHpDJ8C2XMEw6ZJK0CdjqmMlH
P9eUjyLDmjil0a+fRqVtDI7Im0dJTXl6o9vSe30lh+NgqQ0nftIydzJZW1rvOvaQft14+PXFOM7X
LWrriuJsaoxEj3cChaI/cpX+IaEn5fq2Gl5SYzhkxncyvOjy0ougPeDXpmK+6MbSTsYlJNjqW7BU
wuMa5FP0JpUxWFgbpt9E1w4FxJ7nEP3dQYMcUqPBypZq7Uq/G6dGP6b0icaNwSuXPkf/z6bYSLAA
m+w5yjuFtx/WmCnJDyHtay+E3PcADnxeA85qGdG8EbmZKHc0+snzPSKGFVKa8scC9KiXxKoGyaRu
n1K6Hcdq5zl/0j5j7w6rD5wtoqSoGNPRW7K1wspk4YpxU90sW7bF+tI0A1c4gJJFHNi8TIwv5qm8
8TSY3OFTnlWxwjZETv6EgzMWBbgiZBhyTkibMjoqGL/e/6pNGw1DvDRoi0SvzvO8BrbV7gGgI9BQ
HHATivfPYWV9lXEj6GvoxVX5Br+ss7l5HT0FWOWKz+6gS9K9JQ0LRtR8HMCTQt7S3ntMLDFUtBzD
0ZtAYGhUeedG5VeX5hoh3vQSxDG7mV1Y5Q1GcZkpmPXa5mucxiQD2nEQ7ATkwSz4DHpuKB4CZ0q8
wtyOWfA0bBX4XXuoRGR5C/+w2uPkvrzYAcImkh1EXLExWg4lLcvWU0dGz1nXZdPUfKSnpVno1XH1
iYdfC9u8TbKw2H9in9RIxJlSeA0Cc+2Dmbmg7dLbCHPZ9hKEIsK3xav5FkkTLqTH8sf6WE1Wb18P
RifuqtrVwof9bJWwm3yUHXFxi8tO6yDZ0FlwimlyNz5Q74hj5zsvzJXiom1WGepRCRXSxGI/nCWr
9Nk7rmdl4b49DE37JKsbxbHCYDffz0ltd9r+5vyah40TApQitjhFc3/QgujjzFaaXN+8BuIyztfI
C3v+K72dgefPlYbmUDLtBoBlNGivlbrfMYlqr48UACCHHDQCEt4sLsXHEQOvZTIk1sgZg7hF9EUz
a9HAK0rpuYMDsIYQ93qlLfN0b01R6EKwmIGraBgKEiKEtUk7Oo9+wp7XZ3kOwWOL2IAj4o3Flv41
wuWH8MhxaDzopxht26Ms0VCCsPD+RcB423OvA3MnLVvYY+1dJy/K9A5KH/BUCl2uQfNKtTxHF+S/
36Xx7br4kwcvARNhRZg+oCUVzriSNhN5V90h74RNw0SlutGPoeH63P5G1c46VPb6gzDZEVgnKxUJ
ypS8qUxJ+UzTreEEr7i1aB1mSIOCK/g6l47N+iOKUXtbZI/8yMZj75+3q0ysHMa1dvmIfr1jugtH
2zhDg0w91zZz4DZca5jETvf+vpBEvV5v59JHgHM7tIi8FJOufu58TLd1Z1c1X9wZ0cR4vrQI2f+6
j+CcqdncuvcRkZUVoVJ+kPMVeGAvUpX/bh1kfiyX8ftsYczC02WVUL881OQr7o4heb1fTOmQPH2h
15xknwvjKvQzRiwuqXJG31AcTQX3WXHL/2bBUy8i3gYyt+qy0VIV8jjJMJ7DMsBoo68d1HBAWnZa
VzTOPkAmNnC5PTGYnSDkn3ZTRYqsM+m5G9JLiL64dSKvFXLVpeyMMVS09IdxS1XG7o0+AnGEWf1S
HtvuI0Ljc2Nbf3iUhfrTdQJoz00OM62ebMHOhx3vDofWq8G2tOmfjLYKFnMA6uzRt22QZnVZTlqL
6Cb7xj+zdSRBLL5ERxqAnsHo5XOsD+IKvxFP5D3XW0onTsd1t/dJRg0Ifs3gXctW2VUAvLYV6g2Z
hSQSM/6fsRIGmjmXB7bCpPfbSTOx6EZQhnpTMAkDLXH0XkFwOOdomLzfALafzFNh8JyReF19HBq4
KaKqa5D/9z23P23H9SgbsNMZFYFWxQmJpeptreZ06H2jRPYUzGGC3YyHK6b5Uef7K/xwvIwMACEe
T55P18Dh3UW761zKW04xLK+YUMNAYMVMiFquPxxNxWF1fNkwWCbO7BUJw2ZxZ9v1L0X+gRubCXHv
RGAJBwf3Mn8maleLVqBgNg4HGYUohYUFZXscUU7c8qxwcx75/ttF6oFbe8bmZuLrWQCgGKEOHBK3
zQdm9hqK9x768VmsROJEKT/v1zLBWOYh/58vh58CER7LFOg+1bAOxx/3YSW3nKsfPeEi58T/ECGE
W8a94JLGULWuvTNKersoS/DMgGKEb3hmlrhAHH02zLOLvwp+z0yyJlRLEmIv2STs6vNdfJmORLo8
u7i2BTqoskqlnW729CiQX662sOcupOAHiJhRwWUoOMxCr6JV75bIdwrLPiBkO+SGyuAVOI3jDcKq
G+jdT5PjMgPHoi4Lifx0YGMIhhI5lH4ZEqJVUadn2G08PvefqKfsQuOXGF+MAgY4CEYVV3ikRmmR
EQpFiLUB5VbteKIH5OHjBDWoAiVETjOKQnr0kmxf44Jr6OEms+MoxSWSGMfJnsUfZk35UZbFtsb1
0kP5y54V6BuZxVyyQCuiDPbn+X5f2Dk767NVAfdmHD5jF1gRr3Xc9+HzzcQSVV061JrStIAc2Vfh
pHSFIwv84SPUjtHV+nDlnwEppetSvL9E42s/BywWa2iT6D02U03AYJL5KKZ8xhZDI4Dr/NvXoBKy
QRJrwid4vPrJSJuZ6CLRwa1PBmDTbLB913+tNmKzpsRd8kmh04idSTiRLnaL1YaeANwVeITo8UmM
qnwfyfBExXHSuQrHYFqG6rN/h8TwpF5n1sH790LMXHsoJPWhyYS0Sw00dTyRMc3vjsR/VWkKihS1
nA6luwgzA5mzZ0jjSGhZiuc/nRzGuWZtizumwTMTa8a4ygYtxkPDCwNHHtRJGPTKHRMMBPINncbo
geN9F1KKZPFVituntDNHlCwyd25QQNYAddWYN6PrmSf9HPOuxlpGXbaNYofP4DintDw9MH71HTwp
wZW54trCZnDpNVxhotIqKyToTeVq05oMpnVOkDJfqDutSP08n84aB929Pi8aaYxeJyeNgJvuX0mD
dCAl0L72YUF4K4HGgj8z/p6rxB6+AUX0SOm7GDoGTzEhPL+u7T1AuwT+7t3/fsa2wVU7LUvYOipG
M1+GD4ZC8zmWPXZ9JuHyHl8DpZ/GFHyFNHBtkhsM1eb8q040FFjwRsz9Pfj9JDmNQX0ZF+qvuEIj
s9mRDu+YR40Wi/PsAUQLofMeytFij1ZpkYbv+AvX5DdWuKYkVgMwKi5G8Ffw2LjfUg+KIeDDBHEV
0e7xcw3vGozQbxkTPVhzI2fsJF3sUjtaf6wpqDGQ30upAaesIN8pMe2TWbwP3lZccHaAaOSSqkK2
xkijiEMp/J2yUxO73d8XvB2jouQBRoeAtAXJlRVxwbp3fwmuDfsrwjxCFu4wjOhZrpEyquyRQkEH
XGqQxFrm0+1iGnP5EI9zRDROW2OAEq1UlrOwMWM8yPUPSkQ8QgDakfXbIBlWJEe+QjEhRp/CyjoV
Fl/sB5ibLdeXlgHv4Irea+2+4BXhllPBcNNUZg0WZ8vw53kMz4s0XUF7T4aBPRC2q/IuTKf7Dcin
g98STGwd0rcvS4FwEMA3AujQKDoqGEiieeJUudA7FO6kBly9PQ00zLxLf6LGeZRu/dQWtWXoaS6J
vw+8wLxBYJVWr7vbz8FqstQ9chd+J8DrFI9CYvm4JeYx4jfbdKaEK0/38CwPwHLvQau7WIg6NxX5
fpOEnZ9H4EWZM2xRwgCNKB+4T/UzSZE0Br1VtBn9xjAbmHdbkXaHiDKjztHUZZGcnWo1bal4J2Ue
vZv1WhdvZVbbaOtRdtz3tPd6HHR/edUzjySMUTtRHLOa7tfqJSRaDVB/VxqdC5LpzaQzrdOtOP2i
tVhHIriaaIpKfCS+HmGlmymWRIB6JRhqyRsLsyzqy8PGbertZy3Jue1qASf9uHwYnTMQdO0YzNtl
vaGBnvKZSm79r3Okm1g69w8Nrbv1g4dG863ldpAspYc701kwKHNqfll4dKKMLStJ1TgvahZw4Awq
v5SEr32FB8a8XjYrjmy6xLMgoz/APIqYi74ovUjmj8D1P+0AJJYqhmnSPOxkPH8inP+P7pyUHtIa
epyGymiIrx+v+VxbfXILOO9X9Cnv2kVxfC95qyGSx7kiUSHk0/8ZNFQdZ9mKO2xKcZPIy6gIgns2
DQxsreZhvlbLYXYU9FD9UUxk6xmUUx8vqIqka6WZ0M0ml+VNBnFbuPxsE0JzNRs4q41EdSmF9FOh
sBZo9CtTAYzjPvAQZ5VX7Cl+S2ZiXi0ZcpCHuWX7DjtYbAvTMgMGHt/ybnJPMvcui7NFyaMLl438
inre+khe/wL4mMFw6wRlLJrEZt2fTIzThb5vSNfJF3PJe/uutchFGOuzuCNFY21LGJpgFAuZWCxF
3FCoe9+wo78qSbtdYED5oJEpGF4CHEGz2N7BvcBHq7xRuPuqUri5AII3sccBbEDI8icJDJQWcWd+
WX8TsapgW6W+DhuDNgxVjDInY5afMG5s3nz7DEQW6dS+eNlCr3pt/EPhjQanmtrxUwGme4pgc/Zi
70czXABNakgQq+tlRKlEOX9djnLM57aYjY28Wq4owApuR4nesS2FjtaFvfnKg5qwL+ycFFjSofrv
UYmGSWosdt0DErlfKtLwR+vuvwOBM8AO0xtRo+eRzT1mp40+8Sj7UM7s8fpLPs7uo2eJZ525EZ1j
EZ6tuyYSrKVLa1pZ3JbXUNL5H0gW9LAozf6ncSD1Hp1sAKsUt3Y1SKj2SyUvBWmtX4vzJ4Itbm+P
oV8/1fpOynpPv6TYX2H4V4OybgMBWUYQX2iCc0a9SCEOP+3C776QZFDpi2aA9g+C6RM4U9s6/d/C
wTSqD+nzstASVFk7p82i7lxDbQwIgXs5VX3158UHUlwILKs7/hAdPl273TiL3JRe9ArWZn0gmF57
iNG/IglB9Bobp2XlODbFYS81dyDyG7NV4Wpg0VdRJBaY3M+1jGQ23F1CvdHrgVrHGubREUShhTKK
qy6Ft76N66isVK+JX7+sKhMMvKkJ6OeeW/W8Ke69bftvLJU5+/NtAJzSY8HGgAXz1SA1R5Sx425E
/wO7cPyMy0vVpZAD33Lc8+GEXVEBPOrrIwUyT5EmhknALCFrZ3YGzJVppSXW7G+hHxM8sFiR1lhU
15MWIhUrhhJxMlpMPbx7w06Kz3n5wIjUYrFZr/6ZkYM0Yh1fNPzr4c3crPUf0mT5yHw1W0lmP52K
74H6TMUaD07hH88oAoQNm7rCpi3RwJitNhiIpTeEOKAh4fNd7zF3hJp0sSaUjlu75do2oc6cOGu8
KBUN6YoQMvUmVfV7ZlbGgYAd3Pq2mcFrw7W+pjFtDVZ0hKf7iVlU3THV0P6c4T2fXEKDtXyVu4SE
gkIeM5KhLpEPmkOqQ8r+nDeALnomnOXwPY8YIj+2VVvHrs0hsBhgtHFVJ/uI4nMGIt/iteIJZ/hl
/GPqkVRyqhFPiXcv1fpy960lUB8FSRMUw15+EoJadNJbb//Ztw1P4g70MONysAierxSzcR6ezPt5
AmV1VNpFz20OQ0K70LR+j45HhMJMVkNP9gyvwJbHld517cCsjgi4yOqab5+qaGDs1AGwkNG2Ilrp
LPIyyie37i839YDulqEcQBsFjzi5ZhpbyfZPOdZAMVqGqkgCaQvfjm2XR2dPDyh8Mk69VZeQC4vU
9PDuZ2tz+FOypq4PVPFGFG9fgeVosL40Srf8CaoXOLHDXiLZXh5KiM6pXA/g3fyELmBUZpJfKwdz
/vaLPr1fvhd8Uu0l1iIwKa6flmHNVDp62NzIHrPRH/WBYgTrms/fe5MicBbfX415FozTpiMQ4hLW
ua895X0+tnSC9Cju67j2p6PR2bEZ0tAsg6qFE101di0NsPfqqsLDKwCHTwsFGkjv9/VyLczFfdQT
1qvEG6V8UYZ6Vj7DY3Wi3PMTKSOzkULDGHC/N/G409i2vtqGL4lazWaJ5DtXhW2gNdBlvsJBKm3k
23iEQDQfhMbnXjWfllO1LpJpwWKNJX/E9kv2x/0DjHvbc+PFkgY0JE4H00y5VCrQn9te10esswkv
XDk1lk60bZha57IhbXRDe4qHJHBwpe8ETh/M/NM8Q8DWIQLYL1by56rY/dxzOSrq8nYtSIs69yGW
CFvWtmBO1nEKNTLNExEsRXSMSiOjo+48PQ2G8Dpi19aiop7vDxyvR8WmRxI0VvaF9oOU0BaXTo3d
xLzyV/TI1VbJ5Y7sVZkhQ8BwVFntGwRzVezo2STsQHS1l0v/3QXsQEeEGFdv4rMXa8Ec6pQqKl1t
0jienZj9mfgeukL8/iQ3i7gfGfx+H/u2L1x0O3ZeJvnxMJDy2/yLQ4b7MBIcOrfx92jnTjdNeybW
6uYshZ1eaGbaBYmGvu2/eACg/n7/Gp5VtvQJkBf7KxZPbQW5REU73CIWBlBfelRXYCNMsUGehZkO
cWrtpCiWU5QF5z7F9/HIU/2EzznTQbgC+e/kYk7EoAnS6w4+jcBv0uQYJVZGfBDFVDpYOHmZQ9V/
2RiCDaUH9r46JSbW04GwgRJbPGp1TBKuuo7c5O2MJHoCJ1G1YUc4eMzT+YT+QANR0fyM0CXd899+
Unkrs8rXdnY/X8/PxIw1E6lOJITOy39zGaEDI32Px2iedrnKjYhkcIboC+z9C/PcohVUyn4mwQIs
CkaUgJ5zysMvSAy22AArrOI9ryjpU+zakXNh8fnFEWq1Yy5gIKhoBQ//1vfN4DSZIphyV0t/vDpy
xmcj/K98hcBE+0sOZwLI3bEnOXJ24KfbEsrBClc8YW8FjJvHEaOV90fNcVYGGjz55vnFY9N+E9vN
vtH5llfel3ZCnA8PNDZEQFmFXYwk1XdmmIoDp8O0Lm7hZcm5IaJ0pSXU1LtfCFxfNJ39Hpm0Qv5m
uRq9FxdUUOJD3v6M58tJ651m7FU9tG3yikd8ui0qbhnHRXEANQncNNmYpoo4C7/dN1u2fqpOTu0m
Fjfu3mJWofxZUzrF/5TyNkZqWMu4lgQVxw2y5MDUE/8EiZoxq78dtdbPhLLnVfgbQdr9bX49/vdN
4aOcsjbV97EWMeNQvWGEhyMHAOSdDVAyNYVMLvSl9P+wTFDj3T2eUQjJHnFKV2RLOMnMeY/puZFo
/Q6lMMjJliP3hTJHfipSX8EdDgCc6sYGzeWXcaW1UD+28zbZqP2SWTp+Pjz4Mx2fdKWew7vAA0Rm
2xHcnENGNe3LWwtICYCB6FwWhkkthJ/Ib9ooUCGjNF4uzPUuEvcYhnmCFc/RcbDeLxndIcwxDLDU
5phcV3k7yvx88NkRKxnKkHtngiKLRPKo2n8qFeqqMGMSLK/LsuU/2nzMNTNWaH/iFLknBctphtyt
5zTa5OHRuOGkJP02ejIW79e4YfTRTjY6BQTusTKNOf+fAhPLQ7ub64+vtlNGZs2VZH32e2ZQSzNt
B7s35//r5eAvVEUiDn/US2tTtThYAXZJyqqgPTrRc+jqDom9oo/OBLfMevTrcWZ8adrEXZjTsqk6
MgCjVr/Si/B63UWTVVCu4+m/LOgylhSYcurWmowlUNch3sR1akcrIPZ+WvK8U/W8kJ9QWjD78vNk
Zc9im4uh35dHZDalfzWeYOIxkQSZsOzzC5eOroUSRB1cldLuVWoVfvJ4pnNJivch62N/opVjSAAr
lh4DXjYv9BMuEsbnqLYlStPtNuvYK7zc9EVN7kWXZN4jruANzjUS226y3nxPQR0PNFr7BCqcHgmE
68rUtER+s8Tvwbz9pK5MOlLnhpCPdDNQBqgB1plZWxFU6m7cHK0HCWRa22y1ee3yscoXS58hx6cN
dC9G1oQqCWG2talmTBykl+UQHSoTKVgKNg2SPlIHauiWgXTtrW5eTYPmUDT8RkFnGiI32cjB1Sh1
2ABFGTvH1Fv6Lxwliw47P1epLQmJ/4G36YU8JpZShJrfArfjYWRSzpnb9TkbT0LKdJks2bf/8RwE
9FCBqxJjAGgz8/4JmQi0+t+tNSMxzMeevNVykZfN0bktsRXeX3u74Ts63m8pUs0v7YsqnwgQbVW3
D21NURjOmIQA3SWy5/O6lwfhXnzY7n0tjEmROuqgRT01s1Sc30CrQZzC7tz2xZWhhRK7/fzhR5Ni
vMVMRva95qIfIhEjTTG5HI6BnYffkX+yycrtX8ESUKi7zOLyQrGzo2QrvfkE0VpoJPzE8wVV9JRs
1Dol20bQdv5uwN5nN4t1+Urn6EqwHvm3ZzAIA00XDlMdCHkfxSIqpMxOMFouKSILqmNAXQv77qvE
rpa4CsMOFLI/7QpFfKA3sgkIhlBwwZo4sBhmA8GDMMWTCcnPx7OHZLJAZrPfZ/IChCBZ/+2CBujC
L6RfHBRhLVztdQH72lB4fIwxNAVHZeZEEcXniAIUdPX6X/mF5DcjIGEETng3Jc7nhyL0HYZqaSDF
wvbvIwccN5n5ckULWpXjDyCRwLpzF4b1pdEOzMDbo0V9X8Mlly8hfup8r6zVkQq+xNatFWA0rmSC
0JOBPSJDOZxyY81dlF7mbtJQ1M/XUWt/mEJ8xMBH7IwlgLdkdcJV8EZXdarwK/pNnTUh2FYh0r1k
dFjgty71LjCfUnSl/PKHvennuJUlrn47CAlWbS2pTdcdi92eZRC5IlrjOKfFQLAqbb/y09zMmFjF
XG5TQASFvMxYpWKev8A3h7BQQb34h0jwvEnP/6RaBvjWsyCO8B8XAHR8l7adZrBr2xeSN1PylHAe
pVLYXvXiSiiYwP/2ZW7MsphPWWciTbPAYPWsJ+u526NO+bI0pOcJmRoJalHfcElvWsmUFQ4B+Avq
5+TRdF4pGrajlv/EM+bgFl1uSHkTymGxQrufms9JcPjNVmkTa7KpFkO+jZUfv+f1gMgM92tUpO5E
K4TE8tdJSGwU8SjYSHrpx/IhBhC1CB+5vLUfjLd/cqbmeYUlPwCrUaEAQoDebaxL6iBOLJKoO/r8
VnsFp37zcWoCTAbB8wYklOxGvGm9h3ixzAYBElK5W96VhjjLEufrhpILphLVREwgPWa7vA9R+ow6
Y2h4CmoBXdrXQnogcwenUF+ko+LkGkVKxAah1vT06uqi38zYI5FxoEQunqFXuhdSdK1YSEeVZokW
+bKtaxDKBxGpdHBecB4H5u9atTP10jndZkKgmd07s+3KhBMJ0aMptVIVeG2A52tDWzoGNGu2FMWm
RqnJZlZex1UWphxZZiyBlyZlzKZa/UkWyDvG4hOuKK0Rmr9WfANwmHyBgW9bEeHETDDRfJHpTrvK
eeoh7XP2Rn0+kbfFckOBYH/NDTdW/nS/VIPwjtTJc5+XzTE/wWC/BFJ29lFSF9z9OWTv9BGM52mh
ulN/Hhf8QcRVkO/Qz+yD1v8R8E02H/tau+0cLuNiOAkBgxbzUnx1jAxaS5o0iu6MNekskT6TjJgV
3goUxz0/cm79HGX0pK/0tiFY/oPmzC+lauQtkwKyCeNJC4PlCXW0j+hz5XvOpySRNX9IOMNCnGal
mkwh3iqzXvGTbhFuri9cavtwDk/DMREWD1quXMQ7Fp4kJBMlRKGBgqnBHnHWwoyuh3PzdDM5dvTR
mhuCgb0se2tKvBRb6Rol8XYm2ZQOoF47VESFzUpN1u6pfuZpJFSpuZOor8VxD2u2Npxq+3SjQ6rI
dI/AnH7k8Qcx8RLDk0QCiWr74oBmfnL3mjaXJHD2R+rXxsj0WvQwhykxVT1/W6qPjIdP60lhaZXz
08tvPzpDl9tw4kgjeqldpqtIigxnVuGCfakay99lM7QezMfRVLc7DGFgCNBVvz5QGQAvV+G2/n3t
taSsgHU1qXnL4gbuTt5rY+zN/ZU8ok7nOsf+KE1mD9BPclnLGOOuOIuAL1QJjIF4gpxKd2COlmbp
JX2AfwcRH8xzYOqoRpQISOLboOUPGN3BP4rlbkB+vjjL5Q/NIoyVyV/9GGZreCweJrm7hyxIpfe8
5FOAovpcSmhh6TAADQflJbA4hpgXUFRnCdm1AhtebyWhHnV5Hs3H+AieYkzR9kAzCDZCNJBOgDqG
+BTZW0noiNtrkBjBAP4ypZdaOLz/1+RFS47EPDbGmX+d624+s8Sv6k9TDvZn5ADO3MDefnu4xBXG
UdyPo/7nTfXkfXbPHLeVQiYOVIVsfDBGTlqyhAiNlwVRAO5BuT1fdMY4CM2IEIaYVo7WMfRayrBI
LEhewrYawyZU8JcHk7zVqkC5tICipmT4Vqr4/RAE9noFnO871JumRYEBodXF/n7RPPGKyiXu5DDF
9YOkMREzw//rul321lAW5B+dzMZsq/4zf2haXVMiSbok92gv7vKHIaGcrOCT8rr9+Q99RZs2QSE8
swYIGNQEHQ0w5HDd6m0oC0zapfSxt4+h3NvCXrA5RG9/MCz/BBWvhJZiIiCivXoYY3CUfu+GkdwG
F6dfDFunKdvx8N0uCPv0Jy+U27ZK5iNiD34YfCxZIfuHtxgsuk1T4zAMwayezg2FeozY/O5DJpSU
M4simsRQwoQqXqlLJMfk9KUERHggO9x3p7JuYqXBK9DF71Pfeh0DjLcNXtXD8ozxCVmKtX1vH9Gp
sRGIGXR8SqBGYSldOejwst1sdSZtjfx4uXnAl5o27yHn4m0tOqUnFE+SbjPsEhtmdSXHHUg0SG6+
YwxveQkIQXfxCn+b/KgVYyU+voYFY8ijesz0itKK1dlKqXCVfc3IwQl22x9Umorq1AN8qKyQWlCd
X0m98KGfY+/GoS6ZvprysUX3z3MgAWBgPiB8LcJRT9kt7deXfO6mqT+BpkKN2byiZgCKW1KN3day
dKD1pnJIbdrahXvmp1qUvbX/TQhlbdig5P2VAdJP9rJbX1skAheDt7fdJ38NUxdd42KP+gGZizgB
kynH25TOs+3Ng7FBEnJOJeC+z2yFmUO7HcWPMYtEQNZW5KKwO+9AKKiDf5oN8ISceWv6wR8xYAQL
gjWdkD5S0Es1xR73PMegEYCu2yroAgPuYnlL4sPOqcTVuKqYJPZRQN4OISi1YUZnEmorsCAN2Kg6
XOAIf7CS6Xn5JKk5PdUTcmGb34WjYk/Yxnnki1McyHycTW+rCf3mCmB6wx4KHYNfKgnE2QhPw6lG
30vJk4iG/cqQWiQ+NFy475i9fDSXrA9f+FjrK1w7rrQ6S7HBpDF3gx32KkFrJVpDJK7p/bOokfcI
9PeC+2rqtssFpwSKEM/rdkJvN/9QABTw+st7SxOilB+YQxI3Yq528u+060zWQ8CmN9njsOBtA7HE
M48ByHeaivdxy2kJ2uez0hr4P5RgZg5DtAkwji5nQbDgQA0w137sX+luM0xz9VTb2DvfRUJ0J+yP
tUitEXebfkpgjUu9mHxz2XnAwhrwTfNYteWfpXUGzzfw2HkGHyl1wSKOOrBMDrJSCQxN/zfe3o6+
uJWpgQajIANH6WaJ4eyPSIIBOy9PVMnA8rMyrPXVaLRTg67h2fHp9D0kCJeirRqZVYpE2VfYfYQ+
tzOFCH1G+BKXh8FECUcX3eOIhI/eMPfBW1p1cz9FQoYIby1OUyJszH/zgRQ0hcuXnBtUpTlGFu0L
qS4kAry9GhficnI1H0yM1AtTWkFjXRcHqJb5R0zooIvaB3BnpYhVIVgUOQcmjpTAxKy8MFvSpiil
zHJwZHzouQOqOkiVhQaih9VTpBcHiO4KPkqZFfAG9AocyaclmnG6/7L/IH+2k2GIbdcm6VXNYOeW
EOOfeNjJqnCfMYTMjbmwO1GZq/UncS/p76xINUaQ5LzhKJG1Dj1Ix5486FJPK4rh0tZtmFXLnEUp
Xdh6qhx+izVLqmHsC7Gc6Ffen73pAmYqJq/gi4P9w+w4ldjhYFat0KdkeDx2MzpgvbMopwvVwvyF
zZDOC8qs2XOz7nBG/ejm+KzUFaYnq8UyQNO1rjizx3kAkAtyZVMmY4zzH6H7z0Kue0NuB0w9ndB6
MdsIaSXR56KIrIHt0XHid9r8IcUNaEo5HkuSBTgyNZvl0BUflHgli+a5k2GUjUV1B0/0b7cDZzxd
kxSGOCgf9AOshataPhWGFAzOCjfO5w3OAFzLcKicZFC/POlEGdY/b+RPEFLK21MARvRWGyJun7jU
q3d5+dPseQ2gIMcv7lUZqvq4mqELC7drZk1tfZYw45ErrdeXr2RsNsDQp92tkug0azKjI3qIxjvy
BEmFhC+o4WdnAqkHeoLy/kjqT7B3PnJqWQmaiLOYUvg2elJLJrfOvqrTFHRruu/iq2JiHbyx9PuP
Gc1m/UvXwTA9ZfDuDBDY8PFm/bQPA89feMxaVslZfmj73qPJw9IXSI91718mLEoLxeQjtMuc7rgd
Pof5So+5CMdzcDssK0NU+/DSs747yvoZf65YmZq7PbTAO+/0QzLf6juesyirXVRiPO38ublI2cJU
WwGt2iUHHNcvxk6qgQo3jEK3yggmX62OgB6zJoW+6OxdzRnSafHjFYNhcUvtF8k463bgGo2D3ssV
4i6PxQ51K5R1sX6AMU+HTMjzYJseq6WKo0vdcZtJoNcr3cLbf9xCjBT/JCCcqmhEiE4uW/IfKqhC
6O4m8/vxyknEYOQf6LgONYKrdnEUfHKwb5jr/bnvek5b7XAqcUUyFwiTZ9WTLSt+c1KoKL1GH1np
O37GnSxoeGGWWLEYsaOhjtLZM7Reki9TnpCYHLZW+ZE5ADHlFJBojSi7lma/6zbL87ZmJ02L+Gtn
sz/LMeL7QN+YfgwPKkfEXG2qTDplExV9Uz+6Qpylzk09drlfH/LGh/pz9KjtBLpU2ji0jb9oBbQL
g+xHKXfd2YqmAskXp+DqYSttAQCakiDPoMV8RQGCRg91hMMbk6WPBPBmoDdLZXU5lxNdeEh5HXoj
TcgdUQo8HlC3Jhkpm+7OZ1TQ8H6SfYvDTe/BoJwUhlXrXBiX/YToKRYQ5yUQHENusB4aZfVUWz0w
S37BpfeeVU2RsARbH0CDoMgriSwjsCYWZBWtdgI9i29/8/ZGFmhpdor1ezTOpHFfhVLVl7b63FJm
pX5Inc2ihlaCtQNtnfUvMZh9JfUSVlOTwY43hbSx4zy3LDmqW3bY9kg+kSnhuSXeZEXQy3gCWSq3
y4BDq+0mCKXAVqOjejXn4pHM3sRE52boxwu1vGCeDEUwkotE+5mQtBBbHuSH+sXSh+9U4UEillOX
uoeSzeE59Rid8+LNKuHdbID0WcqVcXrfpUpQA6RnkRIwrL7h3tfX8l2O2VqPN6P0LM1NcfHfJCg8
mKH1k0X3hY4OCw8izMiG5I8ROtzEmXGonSZAcKjl4Emuj/C5TEek7KvQVHPMRXg1yOJYHku7Y5Ek
Z/UDDZCzuqkR7WBPXffJygXZamlefoqHKhndWxLF6qDzXzwqw0+mcCjZkQmN0BJN4e8coqBOdc4s
zN3gdG9hUDET2yctBt7gAbfyUr6LCVOdxH6Lfnd3FuTlbDsd8v76xQsjEFe2hT2pgV9xnxjRBa2E
Kh00IkU1zCsLctZOVHy9bT0220SeM4c6gy21z5gL/DYoh9oKoyyM8s8tH3fJ5u90chl4+sBRaRH+
IplJInJw6Mkamn23baX9gghZfx75aVcz3ocUQD9j4j6YlA4LoMqLPYabultHvN9lb5BH7qtBlXE9
C/We/3/FbmU+9r17kOBK5QK4ERBZsUzlDvBCRgHBoY4GHnKSDk4j1pwkAiQ9I2JY2IXjmhLOwtf6
VqKTgm9CTk32hV72pE3BzoZw8ZR0DpmKLncYfBwDe4De9XB4SJ7GLcuoOG36rgHBqp6ZBwjOHR5r
p8rvGfmKiUyI4LBtnj2nNvXQwSz/Fsabjo0IrPGjx+jXN7n8q+mCymagNmSDlQKUnl3IjPY4jNKw
sOswrLOqf/UuJ91S4t8bW2jDSic0EmpmoG1DBmQ9byk6WJmC9TYNl7IsZb7VCEvB4zUIZSz2zAnN
rjWPCMKfK+N7eR/jnZKRP8VvfPjQuF0MLWqdkkeJM8WRT5KvA0Zfs3y6k0EsHmyhMJ6sPRGEdk0q
ne3lwqy+A1RYFIjeUCZRlfjMpZdivytxU+a3+EmKYwaRrf8QVElpC548R/+blBHp2VjIIWeuvals
18VXQ3g2Tn6XEV6KDX112ZYxDuCN9W41zYxIR3oR4iSSOr3TqzAOxCbDRnMz/YNTYGPz/PrDtOdz
F+cywzOS1QRV+HldcAC+ftmkWUJcfFucjjCHN7RilxiF320dy28s46SF8rKXsX2/gUC/sk13qPx8
BprEWQqjGlXCf7EZXUzTmpvfNkiE8UfP82BO+IOiZIN8qGMGHCZIRwrESzxivQ4K7p/9JBzV2yxt
Hk4XYYC/C+4ZOIPYLGKaX3/tdWKFCmnDMOUS3k6BLvkqjKCKSvZ6aQXrAKsGbzgQ+RtdcouY6cxH
8beeoth5kgQop7imse3Xf4/cnSkSAN1MRoBA15DDXL53ZYsorbWCBSBHV0TyxkFn4kUniQpmtjnL
3vURba7ID+NJ7mPDlh96o7ONa6lHxhWn96hJVJH7qi9oXYyyRrfL3AEId4jQu8ogO0X7zDlFfEB3
fNWc+ysHOY2ddBVkp9I37zMK6aFyb2WSUt4GN0YiO+jHqv90aJGXvTeg/cSe3gsY9vZu902fLEYZ
X+XvILG1jLOlCOoyT1qbipg4745qPRFc96MzPZ3gT5uj/PO/Ge76SomShcEVWZ+F9dw15IFAVkv0
lUf0dD5fdeqTjpEK6TINhY7PjqRI1rP/y+LXBLsFpGkWuc6rlHz0Xp5PrTSq5e9Wx3DRR+UNe3cF
vz0i9f4MnpJPjw9T/4mmEUvHR/7sGKfFjYbeXGHyO6hKF2utNf9GcnAF9b4J70idXdP7MyJh5GJY
WkitGaF8wuBnQGMKi+LoYV3eNWbOJv/7IeVcARar+CRVXzMqwhAf7XuVepbIxWE9Z8JXtffH2KYI
nCGNYRxd7i4ymw3rdaoDCNRVoF92X8uRjzVaL/Uf+915NNyjrUtjh9GrROUMrAZm7DcJqPQ5cPGP
zq+3RlCYoSwF4asIo8ol/MFCyYbRqxLqsh/83TVLHc0UIHSOSB6qzwDcnO1IKQcyP2av8xT/kTHa
fg14c7gehO3NpRfCCO8nH2zIS7W5oB4KTaHMHJByg1SwtgJYITIGMzZF87gkNH+Q+n69ZUG824G1
ufqp7bQTo+jT6YLRxUYAmWkY34ZIGlrMjQMBvzN0lNxWjmbk6gpXpsJrcrRwLcDSAwujuXpUCPoY
dwJwaCagu+V9NLcjXyrkS090AO5JraRrG5bu1fSMCbn+Y4lkgSaGA2bCvW1GNbA6lU+XKQS9b8pK
yIvhtECaYUJX/SoTtU2H3jWpjiUuvQZZN7cvTixbSBM+kY3U78K89xTze3ySN1UvR5aj4rrCja9z
s1Slh6XGHtqn2VaSQkLG+zxkhS2Xh3tBBgiF2X02v1WCxxN10jtbmw/roxCsQMqUDMiB/0HnY2sN
NwCL5AaD8Q0KybU36QKUp6fhrnvhCjntwm0iHQ15evrm1lMS0xrwO4iCfCw3i+/Y3guRdbsWHsJI
qTIIGHD6N+PT1Dw2gaS1cqj5JSONYmVA93rma92HYBXD+/OjywaVWmC/WjqeQT8iaN10E2dOz3Am
pHca/HBgwTuIR7Fd5usUADbjgHnk3NkxcZpSzBcnMOisc8+/RoFTtW2EVsG4D9YWPRguFN0JrHvh
K5F63XaTiOLm7U+dFyoXewUAgFjbFoqEdu1XlORCRcCTrXZnNren7IF9NaZdlfADnqeg8p6cUDbd
OwtLdaDwaRqpqHo6rcIq5frY1NPOTGERBxVBYPwxHla+oSQJBmD87m+yj0dLecQjQwCdi6uny/tV
itypRz9R2Ohl+1w19Bcw/uMggb3bn1KuDn0FkeXvLIjifpdQLNCIho/9JKR1uEGjXadbNozgVwlj
lnJUNn7Mv23DrPuGaEm99Bw9BWZBEB4UOyL/MxpA/XhAhfBzSX45Pk04SAtM0g8EZx8H+3lzgeEM
xyut8AbgNcaCIv5o9rcw7rmXlbzwG8VpLhaHKmuGxEcIPKq2yZHBdF67kwPQhXHJtW9uWith8oRD
IeohY+copvrRXYfhuAZ/HTQMYSJYiZkQepyaAKymfXc8J/y6cO50g0i3Cki90B3uh6+ANfBSewQt
pEj3nuF9M32r5bMDbTnSDw++9Mx01qh3uaSwBHO9xMuVJf/QnsAKfBRaVBHW7CXz5Jb41uOkTLLN
3NxyBj79zY9mKSnELKJGqoeHVmAWvs5HKiVPA53eNHF+NcpDEZvG3l4t8yzlXwPEWJU0tZTa4FZD
oRTpn2MEkt451AYZg33YQxdwdbCCK1Ib06HppBznU0L0l0fKaEreAZoE4NMFx/piAi3qPQjIYWtr
eJoBjfig5/BT/3Sd1yilhcrqn86WYO2eGmy5bxUMTEljsMIhMXA9HLjUK4dpyKE1b4O4mdzCBiDG
2HsTElTbqlmr/sVXMPiylAWRTocwnmjxNTaNVGh4yAoZHCBIYb5mtwM31ePFU3ecjbeGGSsQ8QVF
gS5Arr1rFYZYjMhzSXnA7a7S1rN/C0ww/tOK3HDnN8oKSwOlBNHoSNsq/JDcTPhAbUF0LgUlnq7K
Ujjk3zU6P05EkL/akL6WlbVBRHYDD8qFO+v3Ab/ucSajA3lJ+uxeYv/pC5fVVns+axLUjLi4emLU
CnmTX2yUaga3qBMMmFIVeiF3YWI41QcgQsysd7Laa0octK/ADUmRMYSOzhPI4aGYWsn+jz/BYihb
fht7kCedAHTLxbi4UuJmvK1A2SLx/4YLpz3oxfjZQyfZynj2ULJBbG1DN598Ovm2t5+9ah35Ba53
CXkKNjTwBtM2AenKX0QFkqT0RiTS9DvTTOO9yD/n3LD8w74Q95dcL9y6Ck2pnWxnpQjbwanaIfMm
p/gBIYfK6/bri7jAPP9IqMw2PdUV4+j8iGTRxjIi43rEYlo8QfHN777pOvi+Q0ewmcChBPHCKI/R
u35Iq92XzMLd92szvJE11N74YU85etPNO6/sOFpgx0zlxmsgHZr5kVAPypKNGFwbocvcugHu1rQI
V1P1k5yy6ms1bq+t0H0li/cAkDQ5g27l+tnd/O/QgDqbDRNeS4kNR5UmE+gJxfbCJ3hqFMS4l1cw
X1FD2gKoAOgDjYUvw/MhmqLPkc/3ODbl1C5CODb+NA7IUBFY5hHZP0TuRdium1DYcfLmiFlBUP1I
7PTHf+iorc2Njuk8kSM1nn3BbWsZLt2uliN67ZcSErKoMp0SpriEct1A5hE8vu6gAw+Q2hUBgkNy
A6uWmW7RRPHPtMYC8HkCf1eARqvIql50SQXSPxLf1SZ/M22m6hEs/rFBMWGOUD9AYAMOfdOpMx9w
JFKyrS5s2Ql6RJET1sUWFbccDuEzH7Bou9yT769KhWh7k5jie+Av9DVDaWH2cpJcN2+jQL40zJ0u
eIIB3DI86lZqXpbZ90vFE3qB/pwSV7s2k/X6aVpRsuD6AHdrAxb7Tlsspna5SC1VM8aTFMRmlL0U
o1ieKee+Tpk8+VHoF109VfxDdo9l3JI+2r6YZ9F/eObgkRGChAzNxxDAIh0JDttm7HoW26xU//U2
IL4qU5ql++0l7s6FRGHWo36BExYZIEg5dJoy0MdftSI4SixHzixlhPemfKqJz7VcI8AjZNAvImFL
WJAS+s18Dg7xkB+ncCh8zx0+otmHvVv6pn8k12bD8nJwNkCZwzFuDaoSxtictVKE4dvS48m2zXXf
8Z2YEzgbn1Ijoc69ebYdfq98GODPDwSr5U6P5H5nAPrqePvKNWtugjL241QwALtlJhKm5njvkXJ5
7/Sv4Oz5Yhn2/QPtIXovxsCKATxAlZx3yVohi3fFiR9lHYqfSRU22+2sJOnodxy0AuGBAPcczoRb
sjD7waA/9+b8QOmJYAr2Vyv8NXaLrckYAH4gcv9rh/UdKn5z41K8rsid1Wyzzkk22X7uhzbPRYKT
oaraCTjdFKGNRYZrDlX/cuzjFadjedJm6GXDyg1IvZZPbU3MW9FY4MUXrnex+HeqB7EhNYbbQKn5
7ABIA8weCFL/KfL90utTdb6bOswcGBXUvTCWATwJ4oUb29aDmyJdYcJeAbtaCpwUD9C9uG+JNcMe
XG2yth0wIZxmJ4AVm6FgTZ/7OnLhb7H+DC3P/cFWwZ1p3Oz5NE1SqacS+5OqLiDrks84kzkfziHb
YwzEdt2JV4yu72MW+ZQqQVgkwoHaYlTELy1vBBqk2Ef9Op0jpkYHP1lye8jelytdJGuOhDU5mTEn
HoS6VYyH2gGJl0pI7QF3sisZ/KcamISyFsj5Z7xibhfus6L7eVgkX7A2jY3ym6nYYgRUkPjRFuAF
p+i4GQlvgHBgSyRRQo8alm5JFvp+vb60QN8LkvVbK3wx1ZFo5CxpYxfsXttIlNXhduBz5g8Vy1TK
FiBcSwg2nFkyz1vGPc3ds8ibzHiTpZ93ZHTyeWASSyf6t/TVwrMYwGwIQNeNFKMHZeJRf2upetw8
wZCRxDIOVOu725ZtU8Qj43uNRRSCwGrdL3yM7SqNgzUI7ZnZ+1Li6aNzCHGeDggpMcLlDKQWgYg0
WQScI+zCk1NsWfPRjoP2CGCglQmQQ2/htkj7TnHdElv/FwkfDs/AOdB/Im35WQvTK/sjWtsMgtbn
PvemEoNpYg50x2qgDtQomkjqAiSARVa/EKsUHSOXEkJSTXo27DorU6cHrrFCZLKe3MiwkamJBaiM
ZHEIyB7ft9KACJIISH7oaLcBjGpOyj4MU2498j940SW6lVBZ0sppuUN3bTRVJNeJVkqTT2bQZ1Ko
z5cKuAzI5HW7hYtWIFJ6yhzVdmcX9h+sajMqmbgiDldoTZ40qL51QfilINWZlqJW58mtT8rrfu/J
WoWQkUl243GemClavizZ1y0aeceuWI4MRtG7OcNvTamMKHjr8ocPP0pS123qtJj4aJ3fkTDKnNKa
eXEtdU/HI63RYGBm1EOkVQy+3HR0xJxBZ/uV/ieeu2O117mwO4PpUHN05rx2KcOPGjgGYhKo8wRq
0+Ga3oBQ7lj2wlGcq2Sj2U3CWo1UJCOnmtfg0tDiA54NlGjIu/hWWtjrLw9sl3DPZfnEjQE6uT60
7nRSxavQc9aioE+qdbOpGvqM+ntvS+/jHFgY0mPynqMqvkouPF0ZHs+RS1ooBpO9aS3OQnkxdisP
Wb+n6raKx+DFtDLa3AphXvuWreiHrzRO0ur5KWCW3GjSxKzw7T6JrLrgLogE4QbeAZ5tE3/62OVW
fcBq4+U7q6VFIae/USxmI+n7ewH1N9KlGO+76+63om9oHlm0PiPzJNEikCt/ni7sy9w8jI4oduJX
rJGRLCaTfedD7Z7CqrxDE83HaVoJ39V69N3neoPCrQEA0PwGocjfLl+VGeoPRSJ9O6myLDdb5rpB
uc8yTdpAV27ymYgWMKSAGbPbbElGEkok/3h7YJj+JxbyOBvXze/1tkLAA9DPaZPHp+AHD2fhEZ8C
Lp/tEJHjpz7y6DZEyL8AtUsIhWQ9lhen3MxVSWxaeXYoOb76naYnUnpkGdGwB3GNo40FtSyEP2PQ
aJTOlbfV7qFS/nkqJ3Ibh1f7hAJwL2Ah32N8SyxNd4cCR3zZXgQryQciAOYjmscMcsHJNtq3XSum
D1nThn9u6hr15cM71mAQXkRbuM/03GANURtAUJcvzqaVJMg3laRXag6VEmtrLOAwBmYlgKcnjfg4
C6sEcXC0gkRD5dFbjgQrCZ6SieVldfAk5+lYAn3USYYM3aL9kMCNY6xw3avQlWdmlKFI9zLKo2gz
NAyx+hiwWrQTUmISLBvnWAvnI6ZowKNvWeLVUXn9WK0Hba9Rd71OGxvl85ug+0WQt65QgdHkDTx2
B1EKVHaXbvuGLD0BM7+MMuLYZvWD1eXb/N8lTwQQuD1wURRuj/mbeId4/QJkT2er+YvHGFbWi0sy
GcnR9gwVA7aS0I18jZm6dZbXRkPxpjEq9BZDicM97JIe5Aep69bl0jcVZ9Q/NajRru7TQIOfRODQ
3sXz+/O9K3R7dJkwfQd3N26/cGrTG+TtczmOuu/W5RPCXTStqk8eLYbwCBhpWVQW6RioiYWp6QnY
j4U+36hyHHFFiADz97CL3QKOdsH4CQLoxnUuMPRdW5VAO90U6NOLq9u5qPwsAHXFs0jWGeIuPTvg
MBZnrhoJwlqj9tfz3WsLQm2Yb4gbyDZIm3f/UxlhurQT7iwhY9LQfw/Ozb8fVL/kHSwInNXJTkc5
GsSn/niOF3ho6HLnX5/d9Ucl+CXlQP3NW75Sgtu1/KErpZi/NPfBgyscsui8u1WTRQzA/Bdm6sdu
xYlhnZXvR/KlrYkj4WlWO2ORB9BY6YxH3H17seGUmts72UwHh8/ary6XmQTuluK44IOCsuxuORyl
fCdhzshOgA0php+S6uzR5CpUpIOEX532a3io3KZxMbXHAaReJwDNplC7dEygvu2MBB+uMQXH18uJ
TwEs7K2rV+uFxgb2fSAvLIJ1EBceUZGEp6YkdDxKUOFx2U81IeM5qdQZNa+cyeK2K/8H1CsOQ+qy
5O83lzK8UR81PRxtnygHFYdbVzgUkQnnuzVFkBzsa4RDPueT7gEA61/BHZ7P8ozS5MA66nomB2JC
i0RodmoZPNOgftZhWpKJt8oWJrTFSzKc9qPTFY3vx3RafshU3j8+z+4zMZ8EXbV5AFqOJoP0XFj1
ionf/BHGvybx2Ykq3bh028ytBrROYI++4FEMo+Ntde780ph4EmUameIrF65sM16FE8Aj6bV1E+hO
+Z1bnO6FZZbCJ2gQf2vGHG5NCCz5Kbfuy/4Jcp/rjKP+9P90IFmaa9+lmH9EJRw/m7HgtQP1Aivu
ck2OelAoPk7x+DRhVMB2o2629rFlktlpCIBAtA6Jn8zcMoOsx6RTQzliUnPpk7nySuWZjiJ5qjwb
9ZpKKVEc7SaidyHLHHiN+TXW1wgau/qFv/RY6Z4gARoTCjw7Suh3HEpS8v16wYYTTukw4FR31eQ0
0G7FVmUbuS15tR/tM4BmRLx0Mvdq25JWtFYcuawHNnLp21tZONLjz6QBiYeeub1AB6EYY9Nr2Jya
qRRbr82Vmr6lfRiOqrJXDEL+kKYfYnZTUlDk9RQME8K802fjjCIMGwoDZ4osAItPgZGITophdsqf
wn52HHX4qtYlSK2nmmbv2eqztZyeACX8UnPEzfzhUj2FthqqrsAGJ5nDa8Hcw50aFUxkgzMzsK+0
aguatxhoAsl2di5vA/HO8pyuBy7qPP35MM/DiH6ALrMS3L0hQB/qKqtVmiWJ2myzTHPZD77EtxX5
pDwPEbhiBSo4t9BxxwEemURBJZzlbBneWKoMA4R6CqaIMklPgPijIHeKl7T3ZeQJnSvakXyQDYO+
bV/n7hUs04fjYQTy+AEWEHHFHlSGV8PJcTXgvdvWJJgjXI6/ZJVLJg0G/3m1Hg5TXVOLjcsFqvhK
+gGK3vf8Lg5OVCfAIKi7ncDe9du8K31wLhND/NO22dYDHgl8BHxFgMYQNWPKJ1rI2jXB/60ZXoOe
nyV1GMNGosuXS0yaY9XYvBUYCOrPYnJDxurQdRolZcGx6w7j1/YJU7QKy9pb7cULb1sAIDceNg/y
4MiOdODPZtDeJ4BAFlx2txReBipinKkWTLvI2tq301Pzzp2ff8Bq5i900yVbVWDRSxrg7MFtxwe0
v9of3fhcqoNFmb9+eKqPhS2Y4jAGSEtWWltf5mJrVKWcu63A3DasiSzi0LJ90BetEMnevLgyG8eC
u+gIi9kuCGXv27JzypEjZ52Dpo7QtjFQomH+sK0HDIONVhCMhh5hjvPhOUoaEc0xeFjdXsGhqGOn
hfB9LrNqGk76yjhQl3d2c0j4KFGqQ4F/41z1JxwkyqcCyhkiMKsaOfT505TXCaPmx2t6ZiWjs4tk
8VZ3tyXwi+E/imLhpanzdnHlfLjQOWv/ih+vsxATTQ7hkjdYv0hSs4o8FYKVHoPRD25Uq5dscooK
nwAUq8bf/dM8ENuNGy5fH8bECJemgU63O4a5PzVn4M0XyM82y+KRL4vwCeKQu9BA1Xye7UJrHeTz
mQ8NwDDOU6mObVWK7E1R2fVSGBtR8ktbRFrIqaOBExe7joY2UrzSeCL8dt48p0eBoX/7dl9NBNHQ
TZGQ68181+7ICv0LYgMEsLomlAlvYhoq1rnf1MVmyi+mBhPFyHaAZQDf4I8+Ua0pjZaqZVmjnlU8
UPDBSXrr6F2xo1+Crd+lTrb95d6cVKURmJbG5M5m7aG5rBpf2HugN16HBwPdBDjjOh499bdjHRCe
kurNwaZCE5MILid7GCePEWDDCxgeNQsisKqzro7lqfC7JEshgtyAqZ8Fmkbp+CCgO8JwmzxPa9Pj
d+YvlpOPRLs0kmF9XldP7DwGEy05dFTzbNuw4dneAbT8pohAxyqLavP+Fwkj2rjkKvj0I1E982+2
3/52XFoNctkjz1qpzx/B+jLSww5RKspHyl6vKohGjp1xHM/kpcaLIaDR2TTbOapRNSbTtYdPJaNq
9NBp2UOXRfbqTtrrW78nNLVgjYr0JHPAZtmR0DWFiOwND35fu8ViJo3pIb8wLm+KzNHdeToJpLcr
+uzdezKfTLz/Src0rvJ3H5LORH0dWp+erHJjA7tYHzTVGwBkD9K7GfOzAlGavxUD4VTv8U7QWZ94
fAv5OHDv6/1rjxqKE9v5ekF2TnXL4TuMv8Y1aysWrAqzZwY2vz6b0shrd9TDf6rQcsy6tgQce6Y6
IJLviLsV82ajNyV7UxEKrQ+JJbLvT+wUV3nMIXqzaS/10oLFlDbXdfpc+kCLxTk5BxNs7OZ13j9y
qi9g/4V+Ztq9ja3wl2zU6Pct1eX66mq53V4CIBespKh3umXM6vDjax9zPfS8e/+ghrTaUqDnsTFp
DR2w/jF1ZmlgUrZEgjyhS5Nhf4AKXZ6Xqort5HkePYkizj67QbZVoOuyGk217ITyxfYnrBavHpHk
kDxcnerme/v/4OXGWmD0F077wtlS7n2aV9/Gq2TkoJRHMrfnIYAN1eVJifbDG31pcppQfhIUDUFA
F3NBXn8u0zj9Q0Pf69Ce5DG1fbffd6xIiDJeYLm/3E4AJFjTbnnmN4GfvS9SiyqCstCB49AocM0S
vumQ9eL6JjqLqYGOYh2XuH4GQ7gJF8wO7Y/SZyNtvpk2BiGT4vFSikX3gE21mNsclFGixSKbAorW
5niuBXh5TRV4X9gl2+pFdBn8rq5yc0sr5u09W9hC1s0ofyW5v9VOlXRHiHoleVaWljDvV7jaj9On
/17NZerW+1SxDTgM12j5YTGP+/rrMxuaiQ5KtTN4QHOtvnRmLQKoLkG3UwtfK6pnBPZRYEAwjkJN
QpLirSLEbk0K7SV3a5EauuyoODyfzLOTqKtV7JhEldsGVSkY6OooKxI4o8GKxGeX38v2jDODzuU+
PuxlNNt9ie+j0ykQkWtg+7dkVSb/kpCirysskqjpeNmKNIIhh96PGnIFQLirhiLDnzTuXafmCJee
0WsszGSpR9gDOj+gINkCY7XyangX/+VwpwYuHi7bdZ1Hq0td/B/fDSowctXJ/jpLHqqJd7r7mPiY
CJRsxDPqFzToiRbWci05xq5ZUqLDmlolGX208bKjtEB4X8xWsUbCUKn2R9RfMx/GFZ+CcfVPbl+A
kMMxskI6PFZqh95wFjqU5MJHCvwM+RiAx3Yo8+c8vS9IwEsIXsEaqdY9S0Yuaj2hWMhjHH6czCH+
FI1e4gU33Fv2w/eE3pZCZWw+1lKneAQqClLwNEXNEzL1RMZBvzOkLyV3huDdAdufVweDgnZfdxbe
n6EuSHwZ8Jydo5kHAIfYbd6JkY8adzcM+GkNq+6qal0TNIrRzy9HR1PFZMplq/782+YTchEpD+zQ
9JtgMNPvlIkLqZm6tdlIP5fWPaLMQJOmR/X0JUiNlKs0n6RUL1q0U7hyGbceAKRwv8e7V8JZ1s1M
4BozXCqHLC+FKb6bZHIskVtmEncQe/3Yr6e7QKP/zldkp+PzmnoShZkOen/i36cR/HA0p5DMsPN1
AcqOaf5euvrxXUnI9j4VFZR6QFWeBqK0Zu2Iy+U907imOxDUyGF8+8a7ukcUeSNLCKwLq9l2o6wS
GExzxezSgfm8FWJY/Xme77H0D2HBKf9g8orS7SQL0nw3qSYku6eW9bg1jpl4eL9LL91i8o09SVFi
4uqkStX3pZ4TY1LT9Y03/pfld9yht6vNy+b2k2teorBzHvoeeJ1+b15pkvQSUYf3rbxg6PIbWKwG
SEs9L6cHZij01cFTw71xExwSZL/oLCVQXR7p5FRMYFqnYp/Q7rK44hnapo1IjNZ5446HW4zZz0AU
SSwPkRcNks8FPSjBLX28Yqw/B3wHP4CAEnZnMGBCM5CHqaYoWLX4GpZ+GdrZ2iaUNmclFgrtPH59
gz1xwcwtT/BXPv769E9YXHFRYlu0GkOLpJVIyLYn7H8Fy0At7LVCf3B5h8bg9tpiWwbAXIi1gkFH
kz1YuWx8eb7E3mKFdZPz8t9MsUmC3UHjCHbD+9BnRZKSvqFBFNgbQMEPu600mucCf0MhxMavDfKO
/Ym3+4B5sTzFwKAzdpBhTSSOOFAPBuq6xMNRxkcEWZ3fpV+qxWdnBiShexoTUwzwGBulkq14Jjiv
tEPE2dPUUjgkug9BgTIguunGuFvRySvAwzgZY9Wx2Ke+Yuj0X0DLaogctwKROgB97EGJ5Y+byrcR
3MQE7jp3OI5vFfPVCDu2qPVZhEiBCj5HMsOzqNA+y8pjjx2JQOjpvL+2i34wC3HkB9f77Dg+vFin
ZqnY5L9ZVIPwYF62Q1/Mer8FVT1ez3eOpjFNzNEp6Z1bpqvESLtoVv9v8hW3mGMtS8WNXVcY4UXV
LMsbayPAXAiXSebv6FWstgA1bVAED7V0kH/VPGY+kBt+zT3FVyszcepbCHI/6KxGOlhbuHRIud2f
822EsDt/75zvfNId4XP9kscFv0SC33WeebmGRwgB/tHBP6bHKDRT43YFLWaIeyIJ39O2SafwtvCb
itJY/7Ds6/kedImC/TQTdPMv9IZk71lasYb9A3YTs6O26Eifpb3DEow2Uc+dacAu4I+Bi5NsQM3C
hA/Sf1g9ueLd1pk1qymw6SR8C0GQLdlBsYDXbzO7S8mvJV+hkKNjXUgf2m/TKWfcWvUondodVfLB
oWuA8R1NghmGXE0zL3ZdQn2tMTmWfpr2q+6nPngBQnSI1Dv5X8Wzotr1TWav5jUMEzsRbLmk2z9P
vFRDu75LXY9lfM5DoW3eTRlcyg9Gku3knhquyZRiFoLzn5Zrsq4kw9u4d2QJIerYZjgB3tdM8Eq2
EP1yJT+jqsuPzAj8H5RM0LS5lUVL8fX9hUICo0vJsYM63ob/AA+bBvZV1iXD7EhUW0ZxKgSog/Y/
yNlaBYB682DpPnzO5IysCpmLUWaUgqlvdli6f30+B9f74OhOKDFMoftuWK3m1qXx1jhfvuw5+aGg
7vmYRyviNoWzdjvKxAUnvW8yG5dbH3zng8fuLP9pltFmVmLIKdxkVHIF4S3y7hxBuWgnR17nl1mz
S1GCblJRhdRIsfbyLRTjFVHSLJhlIeGUOEJrKMb/phu1dHzX9yqfA76McpjVgWo0g67oP1j6bTpd
fRRYMLHOY30XUuwV3LMd+Eqp+IuxrUY0o3VqyPpsblAb9tlf8hAswba1riqubuQAudQnOXo1rVGN
HrQK1Xes9mvyz8yY0XnUgtkMojbHX507r1LqiF49el2sem8Zh4sXCOb0+c51ZT6xDfClzdNP67/7
IJ/5VMUuzhfg9uzNeOhx+6Sppowa6G2EpAx9GhZw6hE9cDAOdGDVWhFxmYuh95OQ+MqlH2K15Ggn
Db51iH9xlkjdmU/TdodIw3vQXjCFUZK2XG3mVlqls4zBW9fW2fkmdDrlLssAdXDekeluJlOE+kOa
bhxlX+IrbhoZBcn1MmHKoOAxP4zLeUddP90MbLb+j556VcjYpbcP1/TbjVtpv9WnArMnJM9HVVgg
Tr/gXc1wo2PSpGIvPSbz14OL8ZtPxdlMz09DIQKAzNqTWNaMhBHRqhRsrdm+YcHkOa29lPFMA3Xs
0sD1CrpOif/+QvAq3JEP2pZOQsElxSVu893PXeNmuhwHhRLnPnUJE7xSgxZk417q2YkU5OYn6PxF
RweFoaf7l/x/oBJCi7OiwVmtF9+6zZ850jO5I5l2uI4n9My8UQkWY0+zom+PzPmMpVSMfcnIdJbE
pxcYGeLPjT2EDewIwOXq2NXjlNT9qGK6WfL1f3eR17ZDtchgfQWr+bFaazZmb6iTyTn/QN1mTGe+
GdMqEtX4M6pE4jQH5vWAVYJWrfV8XM5L6kwu1iUsl79oK9ClAVYIUgvDyl2XYXVM7QSyKZw0h3R4
gnKtOW+l6ZJwZMRot9wjnPeUA9TQtr6eoSHFP57GA3EZPsjA5Prb0PKPDdvg7auhXwoFas9O+z9u
7rdd+aHiPR6HnonpJMtq/yaiZFHHei1/1Q1lIVbL/qwLk1lB73BFG1HLXkOMQHEAudI10lIlVoIb
l5yKsemrOffau6Yty3E7eIZ03mX9YGhsDxv+K+xYr////sI9XMd/+9noSKDT3RR0MSj1lLI+8/l7
qFkpwSfyaw2Xs9/ryZKTzI6oEXM5ff1IIUAC33TmwTajox92j+hJ6vDiAiO8sJblTauNFAt3S/yD
VDw6EPf3sanv2bJjbhxm2xf0g8j1Ibr/nkTJ2bEHFAXSZGGz2gv2tAh3Apc9FY41H6naZ/si85os
ZmT8Y6e4gyXf7v9mrfmnwh5euClzKdSM3ZP9jJvm/MbLODfX2XEV0/5X3+mgiMFW1PAxgT6WQwMw
3HUJOlQEdg/s8G/snv7istsUyga4PILYbMcLCjVva1aGK//Ccch0pbIFsQpCzFLe/PVIZD54BE5Z
b9INkcBdJC5IAODcjD995BCw6Bdl4TLC8DWLVeEokoTfAvUtJrbfb4Baba/m8lXjAL2nxAyVgq8L
yqeerG7I1rFJv/RIYswOpHUhmlk+tHeQBbqZ0oDEbx+lLapC0RGG2fgQOx8V3M5waJZjJb5cQBgr
TbwEE609i3PWcFTAbDnq2LZ7r44eN79exNv6mWgd3KJ23NIOXQ1X4QoqpIz9dba36VCk2xoQddW5
Syt29q4sRqHmSn2sgwSOgWfWzvxmZgeUz5i4WMO9yf1Wa8UJBhGJSi9vLXiuWQ54Q79bsrdxLSSj
AnXeIntO2mOhqTD8Z743zJJ8+9j0z6A0KTITqUxzar/mRimOSnnPqw9p/TFUmKdPWEMDbSLUKbUm
mkVUYCgoCARV33CpkCDfFfKKIC8JJOh9ACvVJMhwchV/jvvj/U3yuWL5nIek/adJELUyBU1qJF2j
cmc39XbcPWKOiRXmc0d52IMH9v1BDm9A1Bdv0VHZelg5vVw/nDuR4tuqj5ENgNWvILIdszPbF/4g
FYuEX1PE92vzkUF1gMhKDr9iYHF58yvlXx+FyZIt8ZZv6qtqvHAnDGGxN3SB67g6xCh6aiXt48kR
eTGMvYUw9w2OGdL9vZvsbGjNfPsm8zOUpqqSENriV76VyBLDsLnMxF/HAQT8dfpomFKMU4Ycwazv
KVjFsOFR+ma/clCAasB6bNRqWYMEc4xhH2HHyjI5zbg0nyEyAtgly1FeSva6WpGe076d7rwYetcM
rM5Q9RTF9Y66At40wd5klBmY+D8zNyZ6PwTFBIhVHknlKrLBUA0iS3ubGGot9Ps7JCRhsPRI09eo
4pwF8RcV8fUWR+wBD4z4jWe16fLsLzwEpNE+sCMOf6tQeI8FJDY+LePwur1EBVdBfqwwIH3twTLZ
oVRKcO51jOZ6pUOOWaSw78OJHZmSHEs+PymZmuf7BiWoC+uYXLY9KwSX8tgcjLimoUW6zlO5lWAv
lE7hYLqrltVxnAob+u9kgnYt83ik0PNKb5XrLcztbM2iMkoox8XVPMOnEQjprIVVmsSQ0RQYVYGZ
2Fasjt91i65SytBIGKEYZcgk4EMMJUA88NeDQAc3fmkq8Gwk1NHPXQmG1+y39z02jRyadm8QTB48
aFgjuG2E4XugdtqowLWa9LnAGSGYrX7ihCZqzihhRpl9ll6fEIsNP75sQAlwAHx6KfLmEuSoXrIW
T1pvSn+gWg5NajVdhsT4JHcl7+IslC4YHNWqyY5n/E9xDO9Z+RhqQTSOvfyf648SQav7/unPsOgh
0/v8m82dzsp51WymCivhiYMBzUdCxm/nIPPqPnoiffZK2DkOfiP15kv7gaqArVoNlI5/QO2z7uJm
crvLVDTTOhgNGqiKhazRqu7I2CZx1SFzPnt5ZgsPQZl+kwa7psZL479Io7X4NoCsMEbo3zciGReJ
zE9XvMl5I7fUBSoG3EjK3d7Nv7p3FPu/9vTqcwI6fHvLH27ftgWTTKX9QwgQmab6otI0GZD5g2Tw
qE77bCJvMkDUjCFCGmfYLtA8aQ0Buv+fzzhynauN7gE0zHYZFIlD+TdAtWTzwlcIYf33PBfQeaYq
I0pMQdckGUQf+ZWoM3adZwk4c4s3+fVXlhfe2MFty9avX75saq/EPTd9APZPd5PwyBwQ0cmDxDzN
Ampk/aNc897bqq0Ed75rILd6zoMABu54Dj+Bw3xo6j9Jx1idSynI3p++NouepfYXu/4ebFvxFbsg
S0/sckuGGu4S51F1rskgOsZO3gyRoEDQe2DU7mbsUthna25xnJoRK8e5jEz4xjtZl70mzFVLA/j3
3wocPgd63865nmJzWMITXNUMre/1bVoAdPnEqMZn+02dlsPmTnfiAZ866ekdDIkzSgx/yRHU9oAR
dTG1mXsS4/5F3zlu7dOgEI4avqAQ5+eqKmc2uuA4d+W3iYBHtOzbvCTqyz+qT57JMdGEGTFl8Rjl
IhE8ppZoKlwGA7q6Ff1sbmEwFzQvESuA92Z9YnQAvVKd5I4Cf5AnDdZBdynxvJ2Y0VlMp2Glg4Wy
4kQtg4nX71EOtLqhN0s2zDHktEkumSsLfhCmoRUYV3HVCTWpmxDANY8bNdherf3tNbNLfTwIyg9H
Ig3KERitv/3FF6dwM9f0fXC05aCMkMGFnM33UNxYKZhvAD7RIFjAbmFXYzjNP26MFSuMwd45t6KM
p/aAs/QyCsiJQkuMHqjh4tDwwFT/aLyp0UKeTMfIjT5aU6pHBs0h5oiuikE+zT7nZACegj9S9yZ+
FNxhw6H1e6WAiW9AKDGGx3vCPOefDT1/hF2gPuAnEMyrA784wS/qrsl/XkozjYlnhu+ic0s5EUAA
iqiY9dy1xkrJVbL+QMteopcw9CUI8NXut6rajcFEA4TOYzbK59HCftYOff0R+vE2TPmbSP2XArry
mhzot0CJjPYuerVoH6ef6xQeJI5/Qazf/cHDqJKGPR0K9+dqaYRnjPFAfQ8rFXQ3FPrlr9kMmMbM
X3PsrjlMT2lz2B3nwmerEmq6M4HqIofd4LsSt12bUY/dK+8zZh0qa5pZZ/vuaF4jMffWXWzvtF+V
q1syGWolQKeaQIulUkI7C1UhIgGfbLRC6mVojsllpmqCkElygiKa6d3oHPOopIwCWNcvHxQL2tLi
B1puUPr5wnj7a5H0eRDU9Uq/hNI6nf8BQUlFUpcLUONDXEucY9kbqd77M0onmPVN4H1zFhR8wf0e
dPM4VTZzd0L/WTTZ8JCT3uW3MF7c5jdv60xW71qlaJvEVHrn1PYT/gxBs5S4pka8rDtuoz/ufaxK
tq/FjjKiuRjNtXuIjrhwU+Ew30aD0hbKKTvCd+e+RaGKM1A4UfhiXJS6RQF2tZVnZtccXxS5dNIs
mgP52dE1hyBoul8ISrUD+soWWiidLyKCOMsL5Knua/k4JI1gw2L99a10jDYG98ai99JtVW5koMe4
aFPA3JFTOBXPzKXLpF2ZNrPIqQBsjiJJf/ABACIJEn+0Mm0PQ6mcWSMq4fNO+ZmMZmEnxvI/q+y0
zsjVQvig9+DdjEXkkO+iBlU7Sgo9NUUNo7HLhHx5LWB7g2XPaW8NaapmgVavp6kotqaI1w9gS5Eo
lbJbOvlCBsGgZ+3m4ws7lNY8piXgtnO0i+DfxZT/8UfXX/bVuEbC9IEHGHzeIfERfXRzHAE5WXOR
iNjpLO9/R/MgJbwLGkDBP/pYHBENmckGiu+pMNk1guIIBhRoqIk6m2sxaKM8hYRgd7Me08fQ4gMH
b8k8GQn/xGE4yUdEu2UeUwG/KBil761xEKd//fr8r2aOxuxG+FyjAqeRHSznNB/uZrS9+pGS/yh/
AOvWoRbZR9+383Jtrlm3bmXXdxb1W7AJ3miWuBp69OOm95K0LOjOG3cxDDsPz4Ba6OVX6NTalYnD
qT0rThlxhOA0/Gg9MHsRsYxULlUfyrt4hK+sghLz3Nw6Jo+mKn4smrDgQJk5dGiCpDSn8FXSkEzO
DE62hiJU/7aKs7tzFxwhTIRmDlVQNftGxE28V1hVkaYPjjfPMkiuep/HPSMxTBhLqulVp5eT6s8Q
3hLVqJeZ2j34pEUZLu9cqmqgccrKwxH/ln2C5vrWCLAu51aoz4SXHpEUgJxQ+ef8YvmJfa7iH89o
2NBJzvzhEAw8XiY7Spnl30pho91OV0/O9kPKIcB4p/c5+gWoBgZrW+9PZT9QGS5OMH1VbVc2s3D8
Oo0hy/LHSs5hPvyVQ0/8wSOHdTHKixo/3kW+iGK4xGz4pStCK4ExgbZX1/ThEJTaxm1qIcZLbxgG
4V0DRyPtE7B43xzq5HtRocIgEId1OXKAbD7wcd95LYBcd5mPpoyd+PRyf13Ju11kYh3cOK01SC7L
Xtu7QwwQ1sQHaP7Jfp9MWVR/dOjkv0+Qy5+vI3HAhihvngHh4ebONKaDW1g4GnVpyjrmV8Fp+9yx
Rz5drTzSekTD5doJBXr3FuNZhpwiGspcVOI+x6+HeteO6u3T4rzEMdniBYs63mho/10MKBq9WIx4
wo05P/k/9twDVxH8BrXUDVSQ4q8QwrmwZ3UZZlt2MQBPoXnuhb7TALfGNy8qu4Fbvay90L+ddI2a
6+1rELymsGChH7Jg1jvesJcKXp55Td3q27FBoXqM7LEnLoEjKgUFHawEwBACb/5mr5o3kOodFUFj
y2r32wfZNcj08KdXDGv31hRrnz2IdDnDlbTOicL6CEhfA7CBD/qa/1ZRAAw5EQpC2xhCuAs3Xpl5
mJFknNHwlL9jX3pUkUMIoPrURLwbPecNdpbYtA8S5VPs28OKglsDSg1SbPp7btxBfrc3VSACwOvZ
84Y4/ayfh6CjUybN9fu6ZXsJuelZJ2hAwvbYKx4ZuvVTLsy54oOqxSM4lhWIWwX79mlgED3jXjz9
b69sROkroDl6pGgrYtKkpXIi6mXsLsMvfGuIEBudE0mMjyB0yHq4BYoAS3yrd0DZFw9vIfZ5NbVm
okFSat1kagn/wElwrHA6+0Ygxj1ZFAUuOZUOjziJqp24byOef7MCClHJnfoEvRZXkK6xAxfw40Me
ueC18ttIiOKCT/sUlN8nJol6oZihnEzHcd1sdI0rAI1zPUlbZFblLgcZgtgBGCLmErfizi/LpF2A
A3uuEzunaeFeotIOpyAa7irTJjKgnMk7SdKpYv+UXBb7w/S4pFJASXiASbe2IlZsDi1GXmC9ak96
AtuV/NfAV9wUCkOEBdYOfZdtMMN/61uOOIE8ms/sTj4t5PSzFzLJLTgt1f3rAz8XNLSNTmquiyGr
nQGJdhamIVK8/cIJFP8nZpbiaxjr/LCB96Cw1q89UTnf5hrzw4y2ZKXrS25XllhSQ9OWRc/LyWjD
iJTO73JMutkAic4uj0RZzJDg0WKM+PSbWe1xNuqOGvp+kprlzy4UxO5BuTHyMNUBOcQ54qziJOus
IINY9hfJBSJHfg7MTYQtwAPGUeQhF3DvtoQJUSRd+Xtjhlli4fKhStDbcLEKXV2Zia2CJ+tBTwtM
9eSg9qVHJ/MysnklkA0UXkp+MBSdI9DX+gVXEDtU+V4VpYZfsSuIx7sqYJLtXrLkxiO39ePWrAWD
0e8kLRmS6EJafzx278QmSi9QMYYgdG5SRxRKd+f+Ht37nlHHjYOaAKoSSr1eu40WTcaqLkA5HRpI
zOo0eNBWHzVZbgu/advsCNFAPLzwRa2DTT3lKywR9kuQcugWKngxtBG1OP4t0EsXlpy44VyQ5hmi
h3Iv57Hv6+lcFZY30WqvUie/zmkygrkqjkmlrUlavGjeLvzLfJfyeDlTJy6zHl5vuKWbHohyglbC
Kk4oxT+0ykynhz20ziz7CCuUejGYwPLZUCJDwkUqcqODOWt8GgNl3ws7uDettYOAYLak2g0UhM31
ZwipluOCN5dDauN1E5DP2YSKLXMwLkiUB0QBqlrro3mE8LvDhtwU4qYSuUfyseY1FnH9UdZDTrPI
NBKwamRa0LxWXLucSW4Ar3XK8i5gsE5K0HIPaqgHCthzuOPqJkfmRCb02cgFJToSxDyZRT2HS91h
QSvEGJ60EKX+BqP6cbujlQDRcjIjV1PhCPnG7VViMNluTzjz+QNiiy7JIgpuE1K0fNJVZU7lCOAG
qCVSSxMVvvxp0upHk0V2TKOf/nsmoyqVTiOx4LrBFZQ3kOEMJSYyrhfpoNaIBE6wSryfEPxIL/NQ
NR4RhM0lxF2ZRkBXtIc2YurjZYPp86zuejTI/pOwI1CFG4myP7X0KqJrboYbTCvdTM3FID5ulgah
flLPP1P3MKsaiJoWrjhEsZh5bV7MbmHhp2lFrMvtErn02PpD0a3HFLGiWTqWb5kUOfvunJtRlnQw
t5lWufJet7SVY6hm9gbYnHGhu5XYmO6NmJZ/I/drd2WJzJN+PNSblZTXWZ5yWxUYKCla3SxDoYzj
9ChGUZQ/oEHl/nHuJMT6O/CnXz8nk0WMd781w1ZqRjDWckAuK9mVCSkTdtWUy2x2iq60Dv6N2IQ4
8b+80bzpJJ9oiW6aanBoKtukEOLewQLfS4au1IKIhENrXY/P3myjBi6YXB86rQAiXD3BvPC47Hsn
gu+AjCraAXCe1QuE/M/C1B+23VcIY1lFbaoECWmwXH2vsHy8b6ilvJiZkNkHapuH/SFFwy6gr3P9
AvX2ln13xU7M6luGAdcfQlDlqzzNyuvbmo+d1Mep0FIWI96z5QKfWmK0CLgz0yCNJwcK5IP95hGP
aSBkZ/45+9Tvwa8jy+4AtPcUvAVz/9W+DEw0SwHk0YW/NAxGwMDcemT4Ka6q54eTXXYxq64EoV/j
4sZM2HTJoVlB87ksUEkutcPO755h41w7yih9+BcZyzfAAEaECxsPAtkybI5BfEzLXZFoQ2jKpm86
I9fpomWCdgn0RLC1BqElmzJnK6Ljyi/yJ2itsngsgnt7AM+ZuwkEJvmY1jLGqUBFelNY0nSswtYb
XheumY2Jo1beuAgp4mZphiBl47EmrVC+f0+7hiHpwfK7NwhJqzg6WhElRuAfW/3pknY+x0Ar5Sly
3jvFssT7sk8iWYFmG5V6rtKMZNf00Uly6RREafrQ2PONygh83L6LmN607v6Hug4uuNWINP7HERYH
qvd030Hup3jmCsAHDW9RjzDCvtuGJ74zOCNREo2dR1GDUaGW860elh3Bcmf1000BkSzLcXas4LUF
yOB953jRLHGfPu3MziPm8SjG+5wAUH+mecMi98ahZR/mqEwTQ+PMzuKK9Giq3jYRDdDd4EoyDavc
fHZLbxpAg8flI96iv6HlYVmjxOsxxfoTr8WTFjA6d2T9AxqiZFe0woh1MG7vL8zYN42tanmn1go4
WefxQvgkXvwb1JVsr9JfymjZjNGid+28OZBBKz7ZMYFC4QXWjoDc68QKliiTJu2+Qg0G1MdcnLu1
Mz/QCOCI73we/645h2gwN/BtkD0FmjswmMXRpBOAnLf34B/EDtn3Ja258eFlVGhSNTmXyVTc6Zf5
kFRq60khew/6RGxVyUkb8Sm33+AEW/s4egbmvFLhRhTZzhhNoRj/IRUnhhVhenuv74zs9lvyOebW
woO07nis5H7hRm9N9lbi9TcrFgKODl75S5mYEceIPisYbmqBim4Ys2bNSr5xGjNI2BNj41mspeZ2
zQ9o27vA3vkXUsirqAbeTax+FUPUKufCdpGGGJnj4HXRg4dRqe/RXqU+OuwcMrpcK47ZLiOH4FjI
JY7/sAtzczPFegIRWAtk0NU4EOrWtV/ILEQRCItbALYimpRnjdOHs5tRFJeFbCF+B63PwC/KFXIB
NJoxN+IoU4EkowqmasMCKaLJK1+22g88LmmuJbLYOMqdeWDRES9wjycqBv5Y9OPzpZoo0psRZBNp
ruQdB33cInGS9VPfKBPcPFmKQ6NT04UUSytlJTOIXJgNGo7N/L6cswMzMJNWwllpY/HTh3awZT5W
y8pGI5jEu6iTJLxD92+zgeS1UIwlkN0xRz6kqPICfHNlRFXd+LGNiuYyqfHQ5aJD8S6CUM7c5BpG
PpVNYShpxcbq8tciM2seof4ZkmQqHPfQENoc/j5FiwiZQq6CyeiQawzMSvZsns+XI5tEfrJ8KOuU
gpb9CwFpVeb3BQYYIUejVQte2byurwVbAKHZt2eR5zF0rojmZtSrKm4b4BqUdDG/CmQZ1InvEQ/Z
bFJbZoPAIXPUwYleoDxAcU2QIYsrMWai+uB+om/JtiYOWkTjx2Ki2VlR/RZXKDKyY231K4/8yMOb
reC0F0zQiFjUvARrzd7Hdy+Wpt3Df+Bh0/Sis38U/NKKCnIzo00amSb5H/tT9eOQa/OUor3gE0J8
sWSVXkaKGv9fEXE0Tq1HPZlHnf5ALJZ1zUlFfajieEP61teMfH6l35gqzVO4NSbdDKkGUi7ncsBP
iFupY2miczJWX46FqkMtTuIXzmLZnWGHJwRPMSTsrg6rZHNc5B3idzusA9iuSjOVkTfOVw0mZ8eQ
g+L23AeUUSh1emQt1TeVcLIhvz2reIyBSgolQ4uFQ4UZJFQpgaawilZEud7FAtbQXau0scu4d5fL
NGIp8zY4Fyda7KlEH2ipg5rwxqn7bdn7rq9AQP3v646Q9Gchn3fu5uD570pR7MJGe0eB/8tVAW9m
nbyt6/5IfJIP8k9x13umVl7GjN9XTYoBhvNhbEBXO0N07F8vlrjKi0isSn97mWXJB5qH0pjatWz5
y7bYvD5ICdn81Lnlm3/T7L2DWacXFi0bghCNmtwQkvxKf9K34BZ4HjNqRkPO0sQlZUzwwyemPC8B
GTGEs/0EnCYnc3deqpGUnsn6n0BBI2tu5UVpajjXhKaXkScCQt70PSV63ipPfaBO/xZpHJ+hOANl
TM+EUSOJnZAJbbZ977jvqTYgVu2SYcJ07uwjMdjc9Y8pX0QhKpnTxKGdF4yE6RbAEE0tztwPG0pp
hWVbEPJNvOERRg0y2ak4BpEWzprtMFSU20SeAZhs8WWf26adVhlxKDjMnYS1HYO7w/o/MnV6Wmvc
Frx52m7WQgBwEXgg4QodVZDVMf/nHAVFCOQQLgKfyTakUYYB/FCrFHH98Y+6x9zkp1F6YeuRr26/
nvT3gN0J4zFvdzLpFSMQIjoh1/B/3a4ubp8w2qCZfDZ3HKWnByrqCNxxe0pQ6QRwH1UuCo0QeoJC
ZNb2TvUYppji7YDETMQqvNl1pWtGYVjOmDFLqH91k4FwvGHPIlesTUEXSRA2oXseD5aU3b3HSrop
CL3VzQ7MLi/3na2QC/m28Olqu+p+75ki28Qvs3vvQWH2UAA2pmR/wz0CSIIRL2LzBOgdltTs7Mxi
JL/M60g1ND16vyR9MG92XxVAnUIZjTBa9D1PNvp4KSh2KAf8GIFLcYDSslFUEiyeiAuN6uAt3687
JIWBeuZf7jMMgVdYYYESFOP4OltQ//YomNY5/W34z4+3lE2+sjdmfxnFHeWbXd8bcPJ6vdVBaL4i
zX8OV3goHgqLXwMqkr8O1HqAfDkQW3mR1PAtxCBoZFrqRjrRRts65ZLgpqr6fXZ/hZU5hgYgN3v8
ZTCIufPH/N2l4Isb1qIZu7U5fXbcDKxO8hwP2304LEzHPcIACbWyP4UkEmZd+HfziISgBWOsIe3k
GYEH284IMuSKwn3V10LnhI2epvhkxzI1oXK8DTgvH3Lv0erOGjd33Kg4fk4RBvbbfv1L0Co0nRhs
hzr3P9FYjhWfHfu/QbpvobCGiRW5vxue+90HfiY2QpmnDrWezcBJfnFH0qQZC5ov3uspfOQpvBHk
4RM45j+pmvGFVjPPEHR25LXJ7seIFcx+WSuAiVNNiw6cGbLdMH1jzg/7c4ndjll8MacAQik5V23r
FHqxpqfsloHGNNm0Q/g3RznKVQX4EjzRf9mpZzWpMSOKlsIP8uH+ZC19uhy4SoXgKLesWKLYf2iG
RYLyM1AH4TAFxxqYm2sQ44MuiC85Any1oD1PV4UiDJ4amFZLkctRoxLO2U0r7VKcWaFaozLLNjAh
3QgCN6Ils36nfqlXNQb2cuybkr0/8G2xSmTnLPw8OUUlRtoLZ075sdX3sdb+T679X3Sd6rjryRWG
daDxPsEkIX2yDRbE8lkfLpMd/OokxzmnE69N8eyYq3KG3x6FSvklJ0c4etj6M2AM+cjYKzem2Fud
mCGRNvMHvOLGSMdJu/4ix/6YAVDzaQ2jGuGUw1c74OB/Az4WkuxB/HXXFXm9eqkNd7low/blpfG1
J1LnO6mnuYWPHTtsMqgjFDuG8eYfujiq+HtWvnBKyc3a7O6jJmFv4OXK+aE9wvK0p7qGNuO0XD5D
CUsxhyANKr0JxU+P4dcxBxzb2o3QVZ1UXwMkOp27S27/UvbOg8h1t4EKMMjV0Y6iJqwiR/CdtqaS
d+RqKDQcnEKFXsfs/m7ea2wgPboE7LFsTo2GMpeUkIXFlwOf56LMoKSzrX4J2QqYkRMTM9nwWTlx
tGF9zxxop9SUuj5EMiqIBzizS+Lw3NSb1JoWa5794WnKa4mSln8hUo+Udzc6WRmFQjbk86tGB+CA
cVb79ejrte3aNNFSP9pwrNCOWA3Zq5xkbGgplux4T6QPHbh/ArDwztEKArYK6ms6OQ+Pi4y3Fi26
6qOAN87JLFMD2TYCb/89dt/8Y32jWrfeUvUv1/nkBB0mqPhBzfvByzFIgZIXvGP10R4BcSin/Tjb
aS2rr9YC6ZnADtKNjPiD/JUuS/OkMaLy3+YGRLGZ0HBqelyVhfGcvfWPLMGHM/V8TAMDcaycdnCl
P8jF+DIH6ySWh+bAqejZSusewrLgaGLhJjQpfjNJo+pvV4/fP1MTjA5s870SNeBlevNBLzfRNHUQ
k2UkNJBMnAn96ulXRWTUuySKVNBdufzZxioWsLNk8fFnmPUvrJq5jEx4GfocH0evPK2rK7CgY7G4
Mxtuz9U/q4WELXQQt4C8tsGlSkwiDgxnnuihbtkI/fTSitNhxq2MsdTh23GQ2SbiPN+La6b9Lwap
vZ9cigg8GOmzS0kOQUzIhhSY6Yh2V0+O6pHCWnvYOIBTaUFZGdO2swSmaGtD7JQciijpLNfmMtyz
xUvweqf+CnFNKWL2gr+QC2jqossoI+97SJYO8EWORStegqhiOcSYyPFhJCkPOWSQ8TJRVqBFD3E6
zFni+yB77yAfcXRCO3U9Fmm1xpYM1GoiP2y35b1e3ss8tZ/haodHu6q3H9ycN4JfWJPRGhvEQWV5
H9kujGK+rusGUvb5iepGkQ/Adgpqltt85dyRVuNFIieizyu4F8S8334k7cF7U6u5j+ZtHITfGpC3
c1YQT968jvhk80v8qVLUABDuTf68M8Q6tnSDAbdH/FP/l0EuOkpy1cRcTb9WzPwHv3ARHq0p5BZZ
ppZtv95Ny5VFlHecJ0rdPVj6VHfur2nVs0Gil0QeV1glSB80zY6nuFGdi3a4V3JhYdX2J5JkSkoF
9aKYtJSI0QExqcXk+U5wT+9gtEkjjEWnwW534McYW5dm/ER91UP9oVozEHXNIm08XGNXHdzDe6vT
vOUhSlpZ266mzAbEufF6/rLf8B1ijG/K38XTQURzglGTHqhSsFdacv0uiIvSpvF20efn2mtfPBTw
cyIPSqIaRAQkTmqXX/b9dLUOgENdwovQEC9hrYbv9ivYJ110yvsxG1oilavMoh0dawLC+A9PKdw1
VdlOWTu7rIihkCXk6MR963stpP6hJVdpc5udx0SUY5k5NxFnIaL1eoMaZoO8XUqytNUO7FDZBySt
rGK+8qlhPBVDMZvLnvzk1KkgQlOITNcizF+o1rk5X05i6sNy0pcbjavQirv8riyCkajFcDmgmTRQ
Wkew6l8V586cp6qFSYwL76Cmunr0EPo4SXtda/vAvLHaBQZTTUniVkoxtQPQbhPZXbLwgblwyOev
BR/2djMlS5xUrJXblC1XfULFsOZNtOFbirtFsgeof8omSd/Mnl1/UXaN+QLTUYiYMyC74KC4dl2g
cg0IJ/ftH2OagdKrmhbypvCLc4aw5JBHjZoLTTfSccHedaSYbL0KBWfdQIsrJQyn8FejBPgAiYlu
A+5tr82e4fPBFFyC7YeQdcrRPB5Fsmkrw5NXg2tN5W5cXFsndK45mbOdKeqDe7sYnuvprlMEn48V
qjoLpbm7/B54SHeo1SK7s5McCoa67J4rzJAKLQpbEOPPzTidvPXcRjzpzAjEgBGMuuXsJ0hMDeQ7
qM5YYu4az061tCygDbuDLvWg5apGM0hF13PWjBqgfkoYX6g/5NORlBk1gTNTrxOu89oZD46yhy/2
0k6tYKdPZVzXRyNtIlvQwwOc6Kuoh0Xma0drg/PqgSxYoJ8JQ0YaA22IZGeWmVm+UDEIfLCYGHPp
D77UyAccT8YK/FuZiBUpu6/+vB1XM3eYXzoL8QCKfu7VSDQzfK2eqA3xU8wPyFM1vlKgH2LmexU3
Ycrjpk8yaZcpp1xmquXD+POX7jtlB8ti4HvU5TRPUp7V4PpKaxsClJCa31I4v2LCjYg9rdLPZszu
gUDcwo/bK5m3Cg16UsUf5A6gE7ZM0L53H4JhFtdew5D8d9BDfmD/4ODyiCS2nl17G1xklWXySUyG
kc73HSjdlrwmF2yaI1R9k3N5ANq2txt2JZqPXl5QMh4HhufTme5gyGFCP4sWbeQ4473JS89aXwvu
nGe2fIuo4OF11h/u/XWL+PUXs8GMhoEpHEV0KwbW2pZVB76Fklr0yvdyJybvtKtVkxO24pDkRGY0
ktYf7TWgj+nAtMAszutEDB5XatmzgQpHZnhzp1jbX5lMPCS2g5Fp+RFwL0rKS8BAW2ZRp8kdYa0F
FiozsOYbrKyMFoX4X4bKL+1x+xQ8t3EZ/JCmttxbSJxbnpSS+XT6xU82rf94W8DFGRabZA+Lro7K
huFxXX9GMmx4PuehgDtrjOObZiZ8hI1tDpsZfPr74PEdFeStzwfAY5qodOpMP/zexhM66zsmNNMk
wqfx4ftgo+eYr1RLNKWioMGf8t4BZM2hgjik9BLHUP/yFCSwUtV7WjZ5/QuL7ZJwMjfJ2lXoARW4
H63dbVboCtsjZrlHDwfnjCDKToIhUe+qiWrP+MXCWmTwJXCN9cPLrJ6VGWLvdvCo3nRaN3uVNzAe
PR8GVMinfIBdCzbRr1U/zfW7Di6Nio3wHLwXub/s86VABrf4roZtZ+1B3fdD2oavHNMO84YqNz0X
r475/0sFtk+A0aLE2+/jFRwcsFxRWEakmw65ER26U5u/oAWTZj3KfbjDeX3VquFKFUnVADp9la+K
pPfwtYOyUp27GHxgydZw9e3ZBIqgpNatzwZySkeENQmBruDoivqv5R5FfZDs3h8FGlzIgpn+Tq1R
nJiLtVtMBIEMZ/rJPjMgEY7Ph5ZhiSdrD+fgNVl4u9mr/WjSS56gChRVmBvaZyPLL1QD4ZKvlUwY
qGZn/mCTHXlXAp203cGa0uO9TxFEQGiaH7T1k0FeCzmhyNhSV7MmucMaSgZwrEXF9VPMjRGX+cag
whnMLCb7pWTL2aAV7XbcxvwB7zJNyBqNaeHJTXvSaOY5fyREXb3ewAh7nzYHa9ZbtbOPdiF/nde+
VkBEiOOcIBzD/4sm6ZXN51Gytnz2RezKbLjXpVv8LpmgzZx4YW/kt1g7ow+xiTJX6VmK0XKlc5g6
vUlJ36Fs6nFiSCEs4LFi8zINNenJ41qGQV9k4V9gX1O+cEzQg8UTi502rl82SjScRG5aVCFJhkVt
EnVU7/29Vwl+pgVtvoCnoXRuo2FhIFPTkGqTsYhcfUoTxw7hJsy3+j49XOPa6jxgCU18OUVESh51
NZzgl5ZXnFWmocbJjrNKW/tsbYleHYuQrOw8g3EkHclWtL5FKYOA//2Ssi+IvdgIjRAYOSdd5StK
7KkGJtJYHtunmwPdM97c2OT0j0foBBV5PnGZW6qz9X2lEtbqB6obrujBnD6+EbbZ+Rd8sxSTGJI/
RG5h2SByByrA2qwYVbnsOwck7BZtxbfG5scjvRy7RudKDRw9ihvPaEwNl+iFMRn4FRbnw64pPKV5
eLUmRQIx2sLMW+rQ8H+n2vT6GiglISbIzlxtRITdw2OvDLs5MpuqtsQWqWxUnIrtesvPsMyrrYK5
4fJOQxqS7WehL8jq8JgIKi+5OoUuUQd4thhC61qdcXmBHdBBiEQ8kHc05kXbRT4i4b7D887VpAAS
qssinXkLJ4dK4bGJV5OtyLuoUf69GoUbZ0eus+178MJ5JL2t4+YCype6D7byYAx0rof8F9KnfVwo
BBIe70TbtmWjJRoaVU7Ur/J+LGykWyo2w3mKnToyZVA2wraqMjGIopgIRnEeqFQ0lNQFhhX5X5GZ
0YsqeIKCVYojPOWFKR2sPaM6lYD8tg+hJDIR22T31k/yL+jdGnSnh1jKskopZRhd4pEAuJ0APxPc
RA8DUQ7naEvUQEYqGKhKzBDHu9Q9BiEwAqySmrpgVam0/zDPPOZY/RD376Q5aEQRuqY0+fZ2TpRm
q8l09BbTd/WVm0ya/HmuKdTu+aIsNS/15rPQ5w2l82DbHNRc+LfLHkiwWXTNvt99g1iD18WlcIU5
0AlIq3zSQoK9Hukp059/gN7ku5iwxyRY/vc03tcvFaB4C5+Pdry9dAhheELJXS6jWhJzBvMvMrd2
ShBBDBbF5WfqNJCRHZuuqtFZMss/NAM0k6OVaHh4tXPydOwrCpuIo5FjtRW4mr/7t6sCv31/7Ppi
08hlXAorqLbNZ3jFluMYwAu6pQAOBs3F+u3b0yZoFOgbjziWtK4BkXBPmxAMmS1wDwKrzAbZ534p
g+1ND9MDfAiRxKF0CVPAsEUix2qbTMvv6od16x5Orcn7stX4LiBTgsLYPMGEvz8gFwA6D+YM7k7L
T8FJWe1YPQxKozHLJKUfBifR+f9jeI5zNx3bp+jv9ImasIchhQhdeySCOFOwQxr7zvTkiQbUY0No
Di86TY5o6h9/y2vx70MeqYlDKPLVWBlXNX+peLmseCYNOOeCrXENZEB4i4oLdQMh3qucrnEpfyiL
kH4Hqgwa3poRlz/VIrUVb4BL6RptvF8SxxzTr0cENesJ4brmqpCAj3E3fQdBUHQPFZKUqv83fmTP
0IL02ULZpD/DLaXY71fP5fMs/MFIi4XwTBEUBupuRyLhBQArJnUtHkB1sc3KT54lJiVXC9fweEvX
crMkYggNwbbZWmB7xzzyLs8RoIIH29u8QN29xsgG5UM7JyQeDNZz8z/VVMH/ymZs+X2ZXT3n6vAI
aqvwq6Pr261Qz4M1Bz3f3AcB/BekLTmGFpuqkVe94HnIdI0O/StELRXSQPuKSrhjh+ncZUwsp8Yz
tyCavUnlZV8LEarJeBKkNrU0vjZTSnkMPSyhx0GLDUsGI4+AbmsUaxspWK6hHtGgYTqIhI7Gh0AN
QMaNIx7NTJ9mllZSsSBkueS2Ku1S794sCCteSDAkL6jvui1dRoKr3BFOnsCjJQ8SKPtKgqglB9P5
Zm2nu1jgHujlIs2fNFNB53xf/ZScTKJwapeIJNGZs+l9L1putlsbYthxEyImkKVInFH7/wXh+KIc
hxDFCxV6M1ET602eWhpwc5kbHm0PzyAegURz1lc20pDSbQEoh0cWSnM7ds0VeeQf928r8wIHBWJB
xObR2QTJdC4jTM929SzpAEmyzjGYn78df0tkpcc2yx4dB3aykR4BFttwh66iKIxBkS2DBtnPQNhI
IRMcOTbldFMprHOPibmJCLBmOXOl0JVfNo0nOD8FbQl+JTQroeUZCyd2AZyxmPmgKymk0YsvNhKq
4HZ87tq8ayYU1T2AKFiEJHii1P+ckx+0yvLCvl2OZlRL9m6q2W9Dewrawy8h5xunEZBoR8+sHZLr
ZdCirh4KPitdtjSMyHOKUzZ7kZqEdzNosnxnzRSJ/aB72PNF9dhooKbP03W+bxZ05yT+JXt9f4PV
HeT28X0HkGE7RYJhzn7lqIfmJcprc90lLsZVYikXo341FvzWyy74DO0hg4bvM4+7ZwarEF5PKC/7
pTG+IMGeHBefDaj7w4zgFHVT8WzaBLWnHhgb8WWkeLxUE6CdOgHQ3kg75yL0o4pzpIk3/XSgZ3j8
eiQMsTN9sR6nMDhDuVlL6pUTFds8da/dUXbli/3jPiGidEp1DEf0bsCRF11zmCR11EUorEW3HXfb
FiqZPXMeom3iK9+LPzg5h+p+Xl5zELFPJLl9zqR0QIACSovRfW8Ncbqr2Mb8Wt5VdNFT8a1azZ5U
x5908/IpNGsiyOnvvz//jiL29fKasRiK3PpS4/oqitf5tn7LKK7ziwKXnmhqIHMuHYqp7pLtH0Vv
hS7ZzxqcAHtVnQVpWNdhYQxZ7YnGUZnfQ32+ETfUrVC1YyuCgpLJgcpYDSOJ6dleEufYlaQrpgoS
LUuqKiPsxZWVSxNNwoeGLRtCrIKus1dfdo+qNv8P+ePFefA1BTt2s7Q07vPUp17s8oiXMqwsM3HO
frTLAxJ3MfTlJGkEpWC4rXX57gyS9sOd1Zqi3/hAF5S8nvJTj7Yoq/4d6GxiKH2IDfwRfMxAGrp4
K3zT6hRSAEiIpRDHVJkf1g0uMn/fluubm0ebrQu7aqXbkwhsNaIYkIIT0gbqIjhgOjJYS4XEaGiQ
IQOmjfm4Y6w/FvQwW8uZcG3txKdbYXEtLVw2tbdpRINzk5R4Ie2fg7eFBe6yW/xGyZkqaPPOnmLg
Juv0ZVXmwoRmWxFP+RE/b22QJKIJEUoUeBc4/INKht2BFS8a98cgHRQ4G2xPwT06Kb3XqsdLHBtB
XIHGNTHEKclWbcihXpA5OpgpQTkDsqA29Lw7vFWX5VQ3jSKCN8qqHeN2lrG21UE7vTKNParzeuVH
QMiijsz/qGFM51ngwsfp3BqBeQs5wK92KECTjvFV/VF1VP9Vqree5f4C///b2Ms70pov0HlP7EMy
sQ79yJKkNJWrnXWko0XHaB5nYO1+xbpOlQzUTTUbzw4FuLub9uCCzWoJqdZzgMpR/N8L/jlw97Mi
RO/kI2UBm9UDSo1+eT3VQleK92ZZlQ2t4yj9/TEFPwXxcYU11N2I042rzqH/ebJAK2pOY4mmGkbW
G9GNEXFWOxbKsNYz9K4aYViY0tlQqXT5gBcEDfj/WZAcAZXcbE57qYjFDLkDox4Kbl5QdNxFH9A8
NSZAlmbuUGvBV/b9RDNOj3k77kmV5UMr4RmF7l0ry/jj65bsqpmB9TvReIy5ma9GG3L1GnFnUmPz
b4ZOqqIbj5MPkf4bqHwhtsQnbnwB7WTiynCB+OdEwUYqgrVpZQBSwhLgFjSG2bUoO2H1u/GRMYYu
C+DRqKk4QHAJCf7BLAkkMkXNprj4HdM6j8MLgten7hR9A+MkIjAdABvb01d6rSx6yUGm2hMKglvc
noO3ZGiehpDRSn0vyEcL0e2IgUF/hup567XZlYZ1xks6h8r+K5LqwBvyyhQvZ57/VB65MMgqrIgS
vE3jFtixsnVmbIOeRvyzOZ7SkB1CV8X25WgKdLrg5BD5/WMUH/RKt7fRXqBjpAtMf9ju2CHJdnWP
4c1U1ex6PnYjho1jgHCtmKxuSEQNfvuRZoW2wk03zt4sYBHz66+IbGTKFj0TbmLzu713u5zXOLUX
3C49qKbYIzkKYBzXfctLSWlAlultbzP0/ES5dI3PDwEoXAPDB3BAs5WOxy8Jin5coOV06fi31kSi
1jXMP7s9OcaYxIC9Aaz+kfW4A5AZe1PQuzPjNyKVXREEPBXc8pKKjY8+Z21zuGRCezAsNKfr2Hc6
2vSUYuaJFJGm5Ulhs61upNj6zAxFaZBVE3wO3rUNEoBzwpkrWXthEZ0oD3LEijclAjygP9SjQsiY
AJcnSpVY2Ve/QORYimt48O+ZsBCv9rQuE2F9aSqTxMgWjwImA0E5alx/K7sKFReVonFv7cPkk+xI
EfFEukLxvrtxH2/EXUBWid/ya7WfMnLB5Mgm5oqvZLH3HysgszhNVlyJHh4yjSvceKRASphu8heX
LIRI4QK2VpxX7JwW93r5NmSBtG7E534tyVpwQkOp5fXcdfy05PABNB6M1Xeh4w9Vta55DagyUnkH
TuCxerVKw1/iC6/2BTOIxLAlPsVJUSzcVp9Z2O+KIUZGFagdtCPToAf5MAPacnsGnWzluYARHB9U
RkRvAvkbdhZaliuxHLj/Rjt98in4Yd1zo4GCuqh+Pw7/LtwUOCEqznXX7ZU40XF3Z2uYdtXQ1VcK
LoBZWwXAQjcdeXgST9BGrWQqK46MBACBvWD62aeTA7HviDea7r142xr1/GkyrpExuKyCc+EZVTUa
mAnDPaGckK4Zgk/NauafRLBmhhJkEUWfQvZ7U2ITlaH9cdVzz/3y1Kvf1QQXvmCPBEBl96wn1W8P
ae9nl2X17DFpkdH2Tl/a+JDvv+DXSN46YLMUtTikByNlUA9mRGCcfw/gpMwLuofjn2IJQJHXk88v
vdm1cQMyLcrbL0VUXKO72fEAH4bgbASqFVHQ4OE+qRS1+eKkf7zw4Up4f8fDpYh0swhnNi/Ph+Jt
WZdaFT2xUp9qvTvKi90nymD4ght9gviSC8KHzzqbI2YoB+WKmb81nAAFhEY8yMz1qRdLfLA8jkgo
APtooSYgFaC0+/M50jEyYQfndF1VeW1lewiEZQ5e4Hj2cgFzm4cqOFro8w9Krr8Sf6lldsUuvEL6
cQaG8mcFiyrLwx0eoCRujL0byEN5McTS9CyVrF84qHENmGSDVJb6WVmT0BBrCF/uLJ3O7Jz1Zo5b
Mh5zL8MH1n6isfJnLz7X7eDt7z0wrSixlQ7lD09s6EJrajeq3RuH0VzxtQuUGmYtl5De6z213iq2
J2qt7D8SaFfiyyYh0JFeRYGnKa+CMPyxOv1DuFV+fUV76s9LXS+ewm4hznBKBRRGXEky1FRXwkz6
h/35KwnQQBC4yfpdoyNbZ8t+wbFvBvGf9A522jH/NbjonVUr4BwqzZCm/TG/NT87ZISwRz967JMy
IPGa+WNyD81Gp/vtTHMc7p85A75b/1Z8xRl5TfzJRpLe/KJaooaczhfxoElg8ykHxnlyiqfszdy+
R9FWk63g4V+BQs3FtJID5gMQSrPm+k315juNzUmWK562Ux6hQ7QZ+3n8oktYG1f4TbtX+41WrnaF
YIN7M7PvPzi0TQClCDcxqoWWcqG4aQnR5tngFHedLWkrxUPncLgL3GqLD/+A7DSQgwugaWhgfshx
+rvkNP24/KQk/eZsrzNX0tlAT2w9APJS7ZkQiPjCcTExaTgheTu0C2b5ZQjpH+YUtlSaJBNeByQv
RSWhSgBQlaqUUsUve8pgpO1QfT6xxd/knXKlFDWri2Le5sDxJXovOMhuBe/2bNoyQ7VMbQTd0H0J
/6l7nEpF1HzGPpOIBg9ukS8/OSFr9f8dp8HKKRS00iwOPgDl0NKxk05Vp0xeIcc3k6U0rWGBxED4
C0eoCLx022hvryStWv1RtqqfwaL/DsXKsRlVp+rQJ7s+/U2NXmQUsjTJViDAJ1Yopw7pGJlH3B5u
jv7xZ0dtYqhCnyn283pjrlfMjzizab767LTWWRiu03/+0CldEVoLcHNAMZXca+WJgmb4djx2MByF
85vELMCdorcJXU6r4tk/7mjHp387YRei/U+XuEEayMu9J+DxnrrsmWIeTyV8NLv2AgQR/UkLGFRe
i4tCSPJYKc0L0qUPx02TWfjjtEYbesokDXR3w2Uv6M6ucQVU+jNXs95Sl66ewNAREdeOiItPy9UF
gDlNsg1tDrUB6kgXYAhZSsStzYvtIU2GP6wEeH2V+pay0hTI68NhM+MjNZ+a6Ni5arKE99NcG2jc
AyMyHX8ZoDXN/3HpwcvrFTmD9lzcxfjRHpWYs1si5JmnCDKHIL4zv3UpidvqKTQQhZX0KK6WcZXv
r7vxuNR++xik5nGc0Wpy6mXs1dAxWPMXo1ExJhDhnUpiW4wPfg07qDOeQtZ4tiXLXTwo7VR8XSua
dfi9SCGr8vyFGCnxwfrRuoN92SN58RrtJXSVX3aJdSCA74qragkL/fahAFZnaIhR4+9NOFpy6SPM
R2bDJs7SeglKXd6yS0P1fvDQ5L7RbUCjB5sulBqaZ9ZlhPwiuf2kybxNA6F/ZVjrgplVB+Xh1Sdy
NWORslie8ZnAMZyTu8qhgt6qFFA0oQJdNLW13E+oE5STLYZaLFUehs4qqJmEojwhQQlv6JS1ZKT6
fLSdyvtqT6TOFC7vBvrEVncdOvlMtsI4P+dX8hNqGllLhQdiDEmLnqOM57R1u+cTzAhRRH8l/0Iz
FcivCZjTvRGdPj/M0ClndcY4pp9epwLJ+Tx3z0mdwQ2QdB1co+JpDRswUeEpxmK9/r+mvu5TJihh
Vyv6PPu7UW/X+Wr5EfdkuV6NXUh1NM9Gxrt2m/WHTItne1UFIeThm+eT8KzHmdlCOzUSYy7ahA7d
v57RE2c09f/K6su8j60GYqHXvtLowuBd9XxOtRKolcoQ5jzKpno2dAsPUop7B3MtWzmZeS7FEcv5
3Usj5Z2BYXsFoUR5SAQ6MBe/PJgEq5YnMz7Ju2rIIAPj4M2NPfXE1jmv1QYUsyPBn6eUEofRq7CI
AGSwjVqcej4Rht1/OJaj6H+lae1zttXWP6pXnxwg2RPsP8BTHYT3HKlTQPEHRY2aAQscorUsyBLV
xsgSKmmDsefdeIduLmGtat8G7WRYkB+euqe1JOtQyg/VtSzdzHUuHh6AbbIT7JoEwXgCMqGFmE2M
al7KXZNR9TGcL0juGOCklyQQbW0PmNfdaiaUGuTY4tIJpVU8JJUN6SM4jSXfH65qi8/RVQ/pMoSL
Q+3ufne7M/ZwSKuYRVC1702hlOQ9GgAFoyRzXwHqzZEWQPE+O+tbNlMYfWPfB8cgQhF20VfcnAnm
+QSlRyb5kNEE2AyI5sbuIT4MT6RVh89ikbOnuoD9NY3XxN+GKgVi70Cs7zEuU74KYVUtFsH73zob
25Tav87RqxiKfs/3LoKIyn345osEncA/QVhbie2OtfgfdXlQc1Kub09IZuvhIQtSvZyTYKai9Y8U
bnkjFKJ+lel54socVZL/mFnKhfGscf/QzeYTtTJQ0Fuk1SFFnZonehVSvuxWPcsHggDT/1WUg+ow
AlEsUJ/KCImailhvSA3DnU6AhBVOIg+v9cmWMDAObGTwFKTD9h8QNfzpeEa6gWsliSIjO1I5nao5
CbwpUsSCZZxqYUlu8QuyFSaCtGx++W/lqUHv2682dSq1wqWvBCqF8CfWJeOnjHz2FeIIUgBVj/0H
l8JMSP/8Ac83xuEMPF7Vjco6p0x37wXwkbhYmhN07He7Dv2DznBvJwPZ2HUtkKSIq3tF8ksjyxrT
2i1KgMUiLsvHLOWv9MjDnMkLLf9ivSDyJHk7nYv6X/uemUUO91ld7ZF/F0gaSgUryO+K/GCaQeso
ICEKoKpgEgIjnkiVEJHR8Woo8eTOJTkJIyeVnsINm9NP94sSgYWbs0J+KlsGsEjGLQa8hGwp4LX/
q5/CDdllBeK1tG8z4qF+dso+KBLIBhiNopopJicQFZgvsOAhP6/w8BZnXXbU1m+7hyCHJn/Agd7Y
HQzUNnOFjwZC2MGkka4WHU0rPl7CIT+jWc9XZjah/KCT5ZjnBJXU52RnOD7RCeb+My0JDBDpj095
4R/8W/jIzb3oRQAJzIs5tJE0Sj6cCEnzYejJTr5gbL7UhHd70f6c+Rny2p6upEPC3bhi6w2aDWb/
TIP7Dq0nvFkTtRsNxOwkeTNUi1W0FMyOQ7UxuiD76tB3tkfMk83MP22cKG1gUBzaI2R5mEMMRf5I
rneqRKtaPCXfm+bRn2rZDbmPkYo4AsCHQlEbc8XzcgtkcBmsYljw6tlNd5qGFshJoFKxvyYlO+w5
9tk7KqD7DMe8JrgXJKdZq9b1v3sEX8BDT6xyQhlrTlfSC0m3vqACTdItZJ5MW5Y8igI0tE8zExlp
zUcglxMLWnihwnAzNDqlJSWgBw7IQ4UoQyeVq/3BtFgXDlFGiCkuFpboEWZBTaP3rORAkHzNOcl9
hmVhuVvhh4j4xJzQdFmBFW/RVLxrQfYkfdEyZVbe1YnzSIXTKkbwmn0SAgabqrDAKMMXNZYtteZB
D7Ef8LAasynM5edrJH40WUI5wyrpWkSWFTTlWXRTQzEe9No9eUBcY88yoXd257bc8Fhg0cYJfi+j
j45NPuhme9pU5H8+ElljF+cRSEpAL+D0IUk3ONWF8mSF29HxlhYPELViICsIwGxXxYrT3QG9mY7U
MPDzBaKG/qTJAwPYjXZClx7AQduSYy2afkpVUMeTfo6IPnkw6uFvCOoN7odYUlFj8Dtk5z0RfreD
S4k+mwG9w0akgsNn8+q8wwQ3USZefVnJtYkTDXFukXhD/h6y639MQWmj+PQLryCjZo+Ese8LIdkK
69SZ5WJAqUgVuGpAgGsC3wdoNSkZKN7iKT12aO4LJeqk8LqQCmAX6bw=
`pragma protect end_protected
