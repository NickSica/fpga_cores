`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
R1WqgqFekyFBf+R1EmSjRCQxUuOx6MT9aQyodTNNebOe0CK13nDxh2Wir1luIC2E+1RiIa720P7G
30ynEHVRjA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KNMY+1Jln0fE2Hw6EJV59uwRAjQ2BHIWVdMuSpeAltv11pWP/JZCrd4z/uZcVTngSRY8jZzhCZTQ
WJ4MxCfVaXUWBZm7mY0qLw6qcMnyzincQFakqwRdOx84IckfsGjNGJ3OEjUVkf7dW/J0o6KJvGRq
A/P9gVOYmGcnWb2CkLI=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
sL7gG3oizEXkzDHancu7/45cwKfdv4EnXAdeK54QMEX/eoc5P95Q2IxqcI+tnVljSH1drXWj0Eb6
Of0W/iXPKZ8OP77HA72GpMs5rDnQtlgP3rECZlxuTJ9RMJVfJzzO19m/vMWeqMysX1t8PW29rrsf
0Tqwcs84OG2uxBTuyDEWCBSCU7Yk0aBYU4VmF2rkELqh6jo2Q/udlKIUXrwoYSdX0O9uon++5ahv
mjzu8SGK6zkA4uqzG9ghLIe8qBE6KYXQuzvdlMdTVdy8eHbCbzVTNoB6j51Qlq+S5oMMSQvxBaRz
DIAN76FuevwCbX/XKHESsvee5Sen235LJDeW6Q==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NTwqMfOwske0aroynepwGO4Lz00SLylJkTISN8LAcq5uE8ZoeT6aFHS3yIuZsI6EEE3s5mQQ8Cob
RXh00Ler2BvOA4K7lNGJUpMzGqJI7MZao2GijCVpdWL1r0vSvaacAIY9nlusgQmU63NqWs7cQx1t
7NMmVlpgPTHr3KxO5lMNWR2EuXJ0I0zOxQbbrTneEEip68PBGwJFyFdSjQNe3iwSj7O0u1NlI0nF
01F/RGHelGngznubnZikT85LEu94GTbx+WNlMlaxWaxuIaRvhH8UG7MPhsxH6x7sS5ZS9GHBkFDK
gyo/ARDW7a6331M9HUgGOcgw3trs1/Klf0nskg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
F0eZzxJQxbI/Xk9S9oAxZw5Tpi91CrcqL3BrQB2lyqn9Vl25Garq+8JIOwcSUfEju0nEdI9Cvd5l
ooe0NMs4K3iY8tnE+FiNZhFGnmyV5djhXaAeRPiaySzeXAc0nSnoahW36RgdEHyPbHBrMfq1pT3d
S/0aa8cloJNV0EZcGFq/QrhQOhscPpDi8uk4IV75ihx4K3Y6D/SPBsIijokh2lVOyPsWt72NbpFl
R1J6iXczzSEND79HNenePfXgQ1Sr+h8Z2ujGHirxn/++xFCAHxWZmhGcFFwVO7AI15b3pfNiyQF1
2SACCg7/b/5q/JpHGBLoFY5e10UGMoGkaXNq2g==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eShHfvBzKaZ/Wp/QUxGlK7/6Td59dAgzaJsrKOgtjc73r+sFOocLpKUK8YR7XmM0pkfLOBkjrXYq
jGiy10qSwBo8l2eE17VZo8T9nQ0IB2FFGgVl0zNGiZaKSzE4a7K5so8c5gtUyyVlyHWXKqYAj6Ro
NzUEnqMqJPppbTPQbvI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
VtDvfrNdg+YlmytFZV1nO9Ch/hNzGllGY3c+wOLUGxBvYhloxzDDcAB/7/ljwrwghZilvxZm/DJg
2fzdltt6rugwiyCDZPTj9bYqZhAAM0bSdp5YpZP0gTz8EvbCxUo8+Op+ufZee7A2QX4lG973f4tu
FbV42AkOjECD3RCU/zC8zhB5kCMonmYQSEe1sGWBe2+Ga49sur53s1VC1GSUOY3PQLHNqtwSq2Ra
owo+cSlmwu7mHpq7nDvHG8vWLm58VKt4pglBRfC9BYdbhmSQeWT4IcMsVz3wzwUMY4HmFkj+0Htu
JAA3fKLFH4/svF3ilwX+klAmiEhOn+ftw2QOyw==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HHgo2A7au8S1PE/PLf9TgssZhqFUk1LyRHoBPoQd7KZOhYH8iTwJV9W8hjvxzC2Na0peqSJ5zF18
7DRfKJ++XfNw8OtnyxfjOhMGRjIzpk9/xlZOxoCpZPFsl6WTW8CoN0RLlh22HuIAeiFQu4jBiY8s
f/eG3F7z8aDUIS222+2y8Lc0ifWDx1YbNoJritsavlDA9L9WOwq+EXi3pvUCyXszhqfkMn1JVCVR
qUhUx37i3M4UJEKXpk5rfAol3dwNa+jlOtqwiBj8/VnhZxY2i53S+bX3OP8N1Zx5wRoa1UkpaXLd
9XQOggc4VKKTgU9CJZPlRk8FrwN41qv2G8xfRQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 160960)
`pragma protect data_block
eeCl3Hcc/V4mGRBHBrnlVN1dv3CW1AdvJGIATgJUUEol0hkfOJc2B5GKyha38a/Olk7VLganWTqV
HlFsZE/4kRSZJDl1pcgbGBxlLLZbGdN4xxS7J8zAfCU9JODLs0Pz2FttjmU5gTnEjPzkS1P5YSOz
ZHW2Zpzl45Lr8S8HKDkqBwE835P+ZCvGRdawrgByUBI9z4GXqEbZjITN1TjoTw8Qkj5URfvMhADU
v2gXGVTpUnXQXmlcLaMoEtbcKzpEFO9nMaKqXkyLSIG1p18TyhfdEX9qmLyWBWOeLJbVhKq36GtR
q0GeeeE3jlNI7xoqM4Ff3tOSmUNfpDGytun09XE0wNlFvIoCEcbyfFvpU+OgIQihDS3pO1Fk97bz
eqH5t/DggQwKAt8MDjMXjSJbFzN27w9H6XDSYvh4zWOeAjGRwm4ulEsqG3KXunF53M1r4x6r1DMn
lohVTjhHTo3i4pVqH6ZZYYtXUL6EbNx3w6xPNyyBZdSYC0xH2KiGkm8+Pcf7szg615CFJE2QJ6EM
z8YYXJgle1UOP0hQHaDIIrqJgix62tOlx/lszCUsH/I8ZE3BgmWZPTPt2C29vzJz3o+yAM6pmwED
URTS5hjK4iwmWWq3kv3aqxkrAakLlI9PfqJuMxGdRDjOU0/DJwLafsmgGpWal4ob1G0dYXaypFCe
5cUHC1wDIu8Ff6y1n0GxJb85LP4I2VNJNfD/7vd9s+wfXeJpXjievsxOGQCeQr7eEn05Y+vZwH99
XwtiAYZxE5/1NPla+6MUnr686OtTCll97PaviXvFDrD94TdLK/EsCnIXxsutLtxnRJo+iv5TGx8y
c5e1NBZGfyTBU6OIifUmilBNkxNQEkEoeTEBF/cdfXo7svnX9E1JQ7MU757HVZVzRRzHiatkzTia
kVF2Tek1i1nUnCuEsHbclIbCd63l5HWxq9dzSM+bOt4fLTgoG5pw2sDcEjbsHgtKgZvQq3wUYqVE
TQ53/PJu70zOqvY3nUmlAMBh6PPuqVuEgk8w2olRsLWdXpfr8jcm1Qtr5xHOv7XK58/Pyzl1CbGS
qWJN6I2E7qd7a9sRdntcCM+3wR9q9O/tx7+aVeXCveUYfBVbamZUE9/2NfeGUGSe9q1CqXlzWbrw
9Mz0Qp+TD3opSX8znR7PVMvuOqdx8xLQxVqafR15DPEMpJHRuSrB+1e14GLs8AHP6xUGbg1IcDvt
W/UTnzb6yvqsbQ/7kyaAHvsOOajwat9SkV3wJEGZC3iLgdrGfkncnFAU5Bdds43yaHUWTrWi/eE3
fZqejcQuHqp5dxqq5sWYkmwbi28rzXo4ukJC/03/nUqs99CkUUdi1kocwytKo0yelnTx0jgX+4yp
1rB/xY3W7ir0tAPYPmTyYoj8ji45MefTqcAWt+9G+beXKFvkx9rsLpTxb8fQwCKfH2jXawIgwUjH
jjjwuKjjUr5s5l9AnZOtptDrx/5kp/j/zGxQWsKJqfFibBBodBOxn//zW5CzL4NHMONh64Vv2Kuo
UonVl+QjkOPe6fS5RD8k+QXlIgJvGOVGNRCfU1vwXUXo0WSj1VktsKv+2cv7JIwHmPDP0YTW7NsK
FJkkIWksOJPRn1RR+IrsRUJ6jvvb8NSORRKe5lsSyj36e2FFsCJC5OwO8iqqOSpgK25NyRcZMHrm
56kQBUsKMZBRn6uJYJC6jj++r1HJ0Svfa+jM2LMg/sSU6xSCbJBdB2cwQmq7/REv3BCGYJCemsvU
NKm+yGgnkW5Mhfi85cI2CvEpaGpf6ut019ZVIWAEIcIdy3ak+z/KMDmHNW9zLwvNF7Cci/4bTeWx
Gas788yjtmAR/cPvw/toMLOEckT9gnOqtIkAbFh1B4RtLM8EvDxVpEF+HpScdZtEZTDoJ6LwPc5B
uW/5lfyaA1layyLKhrMg8PmilAqJXeP0FNok4tWQmjjIUV+TJSnL+g/amYb1FMHKqkLaezAIoqH4
4HhyUuIUDQfF00ByKo0DAbC4wpip0AZJQ8ihg4xZ5TVqd+n12EVzp0iIjsr0d3K9vzXgy6UjSOCq
iA6x3uDBayCi2AYk+H34bQW8sZDHFI5g/+pEvmDSR6Tb87/M4f37D2p3WFQ6WhEXlSNy/uaCqVHJ
fBecIODP4SFgA8+p8WUctZHVM7FSdq5ESb7StWhxHvGflJq6/cdmqQLwjmgbgdkiWVUiwq3DtZQ2
TuB5mU7do30OZbPEGyXQ03s5jeq+JXdSXTfYXGmsIm1iTWIo9d6Cg2fJUMzu83ZUvUdfH5qdhMH/
iJ5xrpIBmI8SF432n+4DjAtv0TXvPy7fUgA4cy1VZE+hoNLoYidy0dBVIYolei0TpG/noHyiCKzd
SOCnOw+JxoPr3HkGwMVFp8gWmFRUOHlmD/b7kJuHpiCADOtl8ifxjo0/0GOKk98mUMfHILo2SNW3
r16d/xzAC8UxU1WzJCjZu9Fz5fk/0O01WUNfD0gNmGBCgWfKVzUcRjwSFpeDRprwdV9iA3eq3vB+
lXkxs4d2Xt4rg1eJMMmBP3wV+vEKmg1cFGm4ocmRCOkmozwv0ZONstEDUoIKrD0awXynqeiHkTWK
ucN6PuEI+EYykampz7zdel+erkvIV+nwx8vVa65H0UmaX3YZwGA53RQc9FOU4Nj5ZgHnfMXEoEEz
8OF3z3LLFNxr+8osftzBXn37q4rvOl9Ag1ZdofWQo05GpSUlOrjtp2rQxuOeBT0SLXkttErGyHJp
EBMoTlhzwjDhjmh/4S7/6Se39pewgRFD45fTEWwimVrVPpDuWO7A1trcqg1sv+BqiVESLlrXCqzY
XyBhUHBiiySw2MHojF8W6UKSP04bDhd1k7MoWsm+Me/kB7Vj0r4V/0ImmZw8RwMEeSkr6cPc5rrM
E65wCtLcSQwRm7Ny9psF//WT7hwc+hncg/SNfot1w55a1UB8iFlELQG75vSjaVoymd+C7hXYrdPA
LI1S986DxoiZwXIt/rVeHE7wmD6Ky/dsA+29I3lxaTWiA3GzG9Cd2i/vdusqCIp2VjMF+FiTKaC8
NjSJBsowbNk1QNaR8CLED7Q4ucniUIgt/TpgzIXN+yMyHozxfLqqa0faWaGBzJJIgO6SWL2y6tc3
AKOY7Y7fTVj3BjiQrHydqDyVF2UbgUlLhPwgFNHhDz6k1J/Ll+yEI0anCs9MLvWLvmPUc8ZSJ6jm
2a1ltXoWs/A7FPdAIXM0BWySa0sseuSzVR2XofT1vxlu5Je24VJYzbn8DtOXosEiP5u3ie4Cd8N9
3FYpyzFFqTbrvHy2TVREHGqfUFkI4gjd5FHl5GXv9ba28DzTOysUQpGTUh5nsOltKDkbgXHDmxCZ
FQR0AlCVBUle0AWE5GGiNGhUnAeAMOItV8cEiZLaYpBM6ekc9ZwQrFIqZW37KSdGb9Kt5UXAGS9v
4jSnzkoVCFfypfzrol0vJvzEaoGdZcSsLKJtwSaGlxmPQH5T3zJ7SVADYIKp/GEr6tayYeSSi7Ed
PpXIp/PptJvH+whqSYgz/jFxXe9yAfezbo586e/UT5w3YDwI4kmPjoLYhO/E/jeBgpF+GK9U9bqL
w2Jfi+InRFu8wMENYByqvk5n1BexKSp2ivCqrAOLbwthnRiE8HFLjVatM83XFF+cmS4JF6bOr2cQ
pE9DbcArZx2sUMMP9zELHet2ee34Ug6BzYvTztw4tcz71a7TF9T2F9iUfo1d1GBd6gpQjbrED9cJ
X9P+WO2DN96QriaRQxDd0lhD1vEfAwyBU0OpZTrXYx/9UMxUutBCiEnQQXiUI5DJudfUwooPHnY1
yBcEyPr6hSAzgdr5hwBJBRlHniKlYWRp7Xr57IrJt9RhpxlLjdswJ6eJ2ryE8Q1HWUq/9nagX1Ur
kwDZM1AYpGX+Yo0b9WR9l0YLqy0WbvophzIWzowYZozoXcNHLw/HspIDvtzQEde6cBFo5pf1fIji
kwYVICmn55k7uEo8VrUGUOCc9Jf6xVymPYWU0r5ZnmYUCD3tfhs6YChd8ZobLvMFpMWHpQ8+ULJh
4c8bg0Odtdc85jhHGCo8vGuGeE6nixDCj90ozSeqIL4U9W+5Ybrq6vJDTzQAAQ+Y5kQ934KpQXVR
dpO9c3kFNucQbzF0/H1ZiUxbFdS2rqvZz38BURjgMbtVD+P/PxoBiw2iqekDzOAgRvhRCKFrhkPq
wnupSHHPa9X5qlmNEK5fdZi/NTb5I8EgneZJLcWHAJ0VtQHHr96qod8W795tTaMvKaqKu/q6/ixO
bCU1AiTS7+a6bdd7fH8OQUqrN/H36lj84n4uA6mqDmVkWQPm88ai6T4xaPNwGHQf7Eo+BfCwe84o
ij6vPiK1xaLBYfr1pXyLvLNhmXzM41V9GbJ/AIZziNr731Ri7jWmn1FbDgHQumN7BWaPgQxxaPVE
3jX2qBLwueuaGBIfPMRqCcgz7Ar5jvPyQbK3NfgctOBuaf1UCmZ2NgqRxJ0vw8J8619brhIM2w5H
N8kLzCyyxZvuqYv7pXa6BwYloVvE32PtObOpiZyFPWWFr4hdfgJ2koDSdtX0K6R6umP3s6JV9AeO
sBnda8ylxDRdA2mScrfjXbQ8jXByAWZ/hf1rh5YkpPRqokqLDK0JY5x1sSzNidkZWYBYuBRlGN2e
uhRkFrrWkNyRw0BGeY6ELH2XhpWkAP3I3SYnUsJ2VLGzxMQMrQXNEb4jo3k8ikkhFWmZ1CcqXlML
yV3RseveI7q/+bBJxZKXgRFW2JgALygS2mxoV4S9+sRmiAun2PN1IJZlD5mQhCfozC3n+//7SWdK
D93Vajc98nnbp8HHT3eKWGXy8F4AvMGZ45YyKWORPbOy7M+VtpV/ZwKOuqqh4KI5ZHzea1PlS9zv
KryqXBpiRph8DzvW0cuZFp8nzfsp46qZ+jx6xfdixkNfntlUfWSTmIyiZUUlPFtsfMYLwIV5ndt9
DiRbNVvBGtVkJ90vllzVGyuu1uwGEhLXd4EafrWPaPj3NoI0nYo6OCGsLbRnIr8po/1tKXnV83IQ
UeUvEIRELO/5fZ7pZvKBXU4zJMbfOftBHf7FudlY8fetLzwCzqp+As/zI8+o0ooAFTCbLXJdJbOx
fkHgzFsEXiv466vZF2iZD5l21UVndZHQ3onA92jpKI0yFm9hn2a4Gl34S6xfv32eD9Oj6q7PS8Rz
NkM5oj6guOMQFsOoigENQlCkqfztUf5VUjPeNr7X4zpr/cmfWUQLwPNTP9B262WHdfot/lWoxir8
NaZeuzTrkfpjDX4As0/qpMS2FgxbV3pTeevgWAjfZz7xIROmz5bMpDnffp7bqQHsZQiaWxeTeO0A
z+3rmAxaXMcU0ooqurfm6X10ANDi6QWXaPJmPpaWAQ0aoWmocBWbzdSzcD/F7PrG9o+Rc584SwZ/
XPBJEeBLdXo8yToFVk+psDCfAo8UuQkZGSFXYMY1OZD0xCGNkM0GRSR/QzQCPsEqy23JH8QWopUa
QMCUcDumZ7IvllmJsdRkFkGnIL46kfmm533op4DBKhLJobZhc1kI5q8yUup/gA+2VyQNIHn6VADN
FHqXn2nQvM9DpYGAnKtyz7XT+yBkqPDEvqVtzT6FKlHR3dJdJq6aquPEQosj1a+NiX2M0LtEKgVw
4cc+hLE8Qbql5Qaurqw/ArZjInQ7p/PNLL9nJhtkGBNcUWeETROVViWb9S6L1tOAgQobB+UlT8mY
i5rheRm1otc3k6NhgMBwDNpWyUgtQouis5k0Uj8wsxhRyhvVZ0Py07xJimBEW3edIMFhbHYk6GNZ
KoyeK2DbBR0n0Z02kgfvlY+QZ0XYTjUzF12iBGQseAOhfuh/HHPJdgGxEd8HktwUpJqPOhOBs/yd
p/euzq2sws/DbUnNRF+TsqeWEzJsIjH+EAXTmGKf3ZqIetr1TvzE6XpHQU4QjjDCJO/ofjLu80Jz
cMffmGcTfv06vRo0aGoaMq9JLaJtFOMYXmoGBapey6o3j+IJnL8mWzvz/prmz39LmkZb/QH5hj2B
zpyRba78C0mR1rj0Be3yBYMxiz5A83GdELwd5WxTEvz5ex+haUMLK4EEru63amDidVLJmHDlD+F1
3kuoiXUz7RdhleYRx9YaPp+KJdhUgUItM9QyECX325+WI2MBF0EBegyPRx+Ed7FAeOBbpXcOTo9R
dqnGiMwYJ7rRHrZo4RAG9qed2+x9urjttI1gUjn8L++z5YoaN0EQ9yXR7pVw1HdPpctRSMb/v0o9
JUQPDW+4eaCUQnRTsf7HZUPALIQuDEkp5q/jVahIDPnsx85+2ug6t+OBVVcuZEboKhzzgDv33R6E
9Hqet/IyXkJPJlWnDesZOpkVOvb1bApZCOON8nKV2YsOYnvCv0d/uwbikTLAJgRFk+5uJoAEhSBz
kDcvEosjHxmNTUbW0VnGtr3yXpIa7KRswdkYF7OCjZJGk8Gq9jTrSZeqoVBd2RJRz55ARrqXCQjV
BuHBDuK9IGv9bSLewpOrSOvw/Dc31Ocvv0k7kv4NLVp36hh2kLsp4eBZtnkuWVIluKLTbG86z/s9
HNZKMrkXpYFvmgddlMGwRPUCvP3j8y4cplH2WAPTK+hbqTvfSIfrCgPweP4zACwjjncDPwt4RgeB
tm8PtKW0pV7BpQ6Al1OYIhbcUclRHcvoozH2zp0sTJn/eY2XQXqHaEDnCVPnFm70caQnFBkUkzmP
44y2rn3GshGyoEPzRkg9XmLyIR61XzFKksA6TXSGdQ074dF6DBYDbhVxSG/ZVKgvivw2k3aUhbyb
MD4eT/nUw951X2rptHHjB1KXtdAKkB8LboKJWv8qlXQieZkftShdrex5kptOG/G/u3o4I74VZCh5
XVk20x5KgDjxpp0cOhmDf8EW9wkV1y188ztc0pn+l4A15KXC++T7/yW9FCgjYWzg1IpQmdkDSgfe
oN5aUvgCRhDwxnreZbDersxk4Z0gkC2M7M/0nKy50uDVnZgSLQJ1YqKtWO9cwtwxlQj9BYqskzZu
ymfh0YVAsvwEa9sIf1TszcSg1wtNdK4XzGAkZvHOEJyY94ydPIXYc+YFthahaGaPRVMALqaOvNMP
juc3+BkmUVS8r9eC0lfp8DcQ8LnHzZZqqTP4KOy9ChCp9uq76pMnCuAZUb09D7EzVgrOLmxYi/Me
fu49UGHG4oek/CImZQpFlwXRyADhhmVekfd0K1GrSRayEqRC0DPPphSOXJZFjlgyNGor4xEFPP9u
/THc5biRcqloqsKw8pBiFdmP6NuhoSvVYcq3XfTJdyK+pcDiULlsfjlmg1vXlIvtFLyuN7wQFkbv
VvP/6aaSo/ZEWC0qgFkGMtR97yY6JvAuZjHdEfi2mQq0TFkJ1bicqmZfbZjOwfQv3S97qSDWwUMJ
t2HKO58ABJfvhqcX7lj8r+lod4dL36N3dq0eJjSFdTC0Jfay0UE90NCkVZl9X/Zig7wi8fe6WLnm
hsXKx3/lHND+iL9ziBn8H5CaTK5mqwL3FhARsrycsmliI7Xcb8rIorqxMbeURR5NR9qro7+/Jva+
q/gobWKC/+f5VHeHdxyKsEp6lC7VnW0mO7vrj9PmAsqHCaQNhgPDZkVVHFHNsVJTp39wVTaqtZmF
+NEYJNo9CZA8O6jj2UolpG/BJ7J53FFz4bLYBhk3ibDwJRoJ4FfCBJuuJXRQOwK93Go6+DccFLE3
PgxXW0uwFNPgtsAscXsG6NE1kSD9L3WhUwD3MJgeXF8s6Z1PYYTmigxbO4zeUs/m3soS34fNLI3F
MPqdr1yO1eo89VbC85K+xhllj9RzPDa8D2EXZwQqXczCqP0IYkXWGd+Ti/ysrCQgnMJIao7/sgcQ
2z5w7oyVFNEQRQW9kKZyr5enhuNr+yeIg2TZwVSffOYHjBgJsTVN4c+ak6rj6YqxVJg67R0LSuOY
51Oz07HRqEP3TJYTa4EIoCi7tdtLCxXmIJPoaJfwyqt/GyiAf28brmac6MPnsPHN0D6t4m6mvNeR
4AwG8aAZ8o37ta642JPxftTSRSxNsYsl31k+II2JWHwk8nQpgLmmD17byA9RaIqb1l6KIgkE0ZSM
1q9dVCC67+MRa87cQiCorCXp6Eqq51Qb2mvvt3Ix8ACPrbE6zJQS8hBdQM3GVE+dwSSxNc+y+P7e
0LWQOl0thM6rCobPFScC9uGOO5evMZG3edMx010iFDTd+NsYkibMycevQlDV0M8G1/qJosYA1LW0
l5KpbLzkaWFGBdEotTTsjFNQP5d0Tm9T3uVaRW3Z9dFqr2J5zOw5QjHFlZGsRYkmUVKQCxpOAIlL
z42ebXSq6n0omDf3omd0CqHOJDJIdSvYiCjCOqHT9jdcxsq6T4OdrB/zRs9ydjXdFaJ7uEjbv1jA
ETmxpexvxAks36my9uCLpYTVVAiT1LZUPHDYkMJ5WL7h2BN1xn/QeIWDJqScsEIY+l5XQk2FFhNg
lyhAIISOKg85gSufx51wrnRflG5VuNQT1D87kdWGd7jO1pycGm+iD5QKrvkVTGsPvLW5kzBFMNc9
dyfBt1qXgXK7ceh31JPtucyzblJhvIoHTGRBseE71WnsApdiUereI+T4OnQfLUkAsTJUbu6tUBm5
E1jKHMGBQy0AYL2H2JsdNS10e53/IKjDMi6tUm9EmUjW8vKFCOUwWqffdXkDtS8BjIop9kKr29HX
wnqZVJX/IMP93rOj9zXHcj5Hn5K2GYGeVoBcpIA4Vs0elLilL4n1kaDetjvNymuOoS0WQEPPQNfY
o3Z/N0TH7Qh3R0FYU/o6ujejsa6eJDi9z5TOVhq0GVBKVvNar7jQiN8eKEB/XDP2TormuRC3XwSJ
5AgjDTcj41Ka18P9V/Oav7yYjPojBNVPqjwI8715VswV6Zk53JbFMLqFtDUpUtw3b3tREHZa2GwK
tVH6362xZBOE7q/RPf7qAwSrCqxAz+5FBKiQ4KapgRY1KsWxnfO3g8J1rK4+t4yWyNqo11HW7YKf
zz6gl9KUmvqz2xH2QMbKgfUY59gG8omJJNUSVqgfyEIxdweNSZDIpo7fYMS7XpoZe3hH85SpNs3I
nS3Zsfqzywkn7fPKqTXPx1DPCOwyu/eBjEQy0ZvtdGOgcYyiW3lXspW5mBnKl8Mi1ZTxmTLb3Kvp
0eg69siLu51dxRF/F2Ol1Nro5KOHTGdKoxuTesOtS2kJc+bJOejbOlgJvJeeYPzDoB8dK2RFXNHL
jpQiQg5CIiZRKnZmGChVTCO2FiOgnrQYAUaeLRDv1pufModa3kAC1zX7xhcihWFmkHHzxBEsADU0
NuUz3cqMDndzQtLYYrkiBlgH3XDD7R7xPLoW2+yuKr6eTtKp7FjsJT8GRMDUw3k0SZS/3VJ/rG7G
tZ80G9VmRVpj1VT5RA/24DOk2hWZiTp/QF5/Y8Zz5f0xdDe4yBCZXjQRGcq4KFKhCk23VbwLibhr
J3gTEPko38yg3uVc7gcFINXIubR/BiID83Hx3ucW6J1a7mhTFH4nSE1mNXR7F/WJulQyo5NS76Si
0q98pUcAmt6wMpGOrrZdpaQ6StIIGrGWFaEpcUh6oS8/yWvwYfEg6Ot0BejL2hZIuBzE1IeU0vi5
Jd2tOhZyL+4/LjtpR9gsqu8LoM5ITo9zCYHRnvYcJoCNCztlmgCOyyLilH0OgZ1z+2vAZ+Y9asNX
4OkVz3HxUgE0UMM65d2AjmTQFbarm8qlTSROwEg1/HEZxejYX4KQBN5UY65v8Lib4hJo2AkkXfX9
ACdzqS1XWFSB0YB1JmvPfZdbcnxsNvHgrQhjdPTKu6TJzXgUK5gyJUPQwE3T58TReoiljz+meAGk
PY5ztk42LOISXaayjo40Qo1AcGIAuptci3E6KvpPs4GXs3tPKPZcZKS7sbFf3ipi31gCY6EK4eGk
h/q2FBZaojg9+cXLWcC7FBRRCdMkxb88GzQ61sH8O6778eYpqxBuqOBN4EUmvXmppNYPCdMHNwYr
IJuVLp+3/4NLyPduGyl5ifOGdKcNtVjMdDAmt+KaJXhYRG+PN4o3Y1ovV2ypk2WJgxAnS99W3YPg
GQq8OMJOQvm3jZafofvtJFeaSZQarlZkv8BBOn8tKPjj8fky+yCBiM55sRNCzFLRdADOjK2Fbn4z
CAGYkqe9EXeDjwUN6hXW4mW80vo5X337R578WOp9Z2DGtK9EfPieDTFvYzM/6b4iyvTvzedI1Zry
FMurL35e0vZ8rYCokx5mJ71/uqZ3jUcoWsvv5xvZ/RS9tTCpAa8xrDDXEZGRm+RPJXBM1DEtYFzh
Ew4myp2Nw1fPf8PdVQxrHc9G8PeNrda/IrKV4hX5FpgIWYWJqrW2ZES6tCO9FMIV4KR4+4Hp1wX3
hRfDceg6l1Qr73c5JzXDV0Nn84lHbD+h+xw5EeAbcBtJa3/YdCsDCjHi0GiDoEXhZlCX2ICKZIms
X34Rhtl5+O6/PPuMY1FgXnzMqyzKfpVzhiiIaLDwp6bOmPD5oqfstMyljDrbY9Qzy/ZYAGblE4Lo
eRlujfA5T5GUZZ+WTwdYKJKMUaWWn6J3X3o1U6ItwtfcoX9mZ9j2xriJKM92TivEUZ7T2Yhzb1LS
53en+Io+2tNBcytkj53lFN9GILLXnmJoz5UNf0e0k02S1geQ/Eyi7xCWBa0YecPlzxi6nGFBNGwZ
SSvKUcWjjZaqMSa0GtXmwgu1/fEPEr56dzbYCOPLqC8G//hewQ5OsHqHfxtz7l5PDkQNwr94UDND
+cRS16nwbVVA9tCZOrf+ium8CNDOSbaKdsoHosywqjEKc95KqlB9aLFpmGKzqF6lrFRtYK8RAsgK
+3Wrua97H4YJpi4tw5KplVMjihRvEdZ8j55oE0aYWH74VBZCullV2A6oBsmeuv6OrUSQxC01xoN0
QAWE9Sp8vcfuofEKamPJUGlEY8RgKMVpf3xR1Flv1CwaPfPtei2gb3q9sHe/boaIEoYdUuZHG4Np
rU6JV6vV6WuyE52elfZ9t1Xk2QpnynOLukKgPgqCbNa1Iat/bHeACun2jdW3ATACFUhOk2fP6J94
DCIBODnSjP6TBY4aL6UAvfc06vDicbUI12LRQ1wyIqAbulAVMxI19JD6if1JS22thi/y9dizZGT6
fj7svMz4RoHqOXupgTAQDnthVpoyHHWqaNQ6ZmwD/KNjfbjFzVDLsSsQ/Stnluty9U66SzWYAfeY
zNz73vu3wldWE/+gh/1XeoeBpGvvxlkE0LwWqA9DG1G+OE0kX1F1kdKaHx8yiVlc/+MdvaD6G/Ac
SV4tFW70Uv2nlwsbN6SfG4kdIs6H5P8GcAHWSY8Kg2CuHjr7mfJ01hDwk3qk1YW2KSYrfXD3fKIW
+UWxnsv/a8DE4dHa7c0m/isnRtqzvdQCY8/3bYamNCtXRAvAel0aKVInBgeko7PPkr/eo8VLsbjq
u+1jZcC8p+uJjdXoNJl39FjCy5tAiGGnIvoqMm+SfU6wGsOl1T6rkhq4175Q9dMHQQySWt40xl4f
tppeBnXGsNjJcfCNA6g15ZnYnJwf0A8ij+ieW3JRHgiw2DGzTVJKyOPBsAPyRnn18WmqFWwnC75G
YsrV3P6Cq20a2HFTOCrtTARQbciYb6aGnonXohRAxlEp4uPDgqxcBtvyzlKM/eYaCewnqrH9GK+y
kQJXAEl+9SxVwY9WQp5E32tcum40YC6W2OKgGQT2ZJ/BGrSbR45DjrgQLT48EPoRgUsYml8S6uGp
Jni4YunzisVB5pYwfKVORmy9oTXA5Mi+1XrEOLjnpXrCPVKEQBV2enNxyKyoZxVBnwXxW3g4QSmq
o5FZzIUerIvN1Zti0sQj7TIh5wn5ZTEDwxpvu17nLoXJkWwglRolCq7ulVeEShM9TX0OQq+TsgdT
JAgvqI37/SLxSg/Hz/RbP++jl7spndTrnZco8lolN4z3LVPQRQkHHtKQX4SkqTUHGskzkVqlMETu
slW/WBzA3JQ6H9YayTEkAr/u6YUMGHBPhX9QXIvzOdNti+rw3lLpmJiLgk7RQ050MThlQGQyb0or
HaQrm+duqZAkBRyWeMSrCYwKEztqm6m1kUJZ7QJ41kA0PXNAGIcC4vX+LuO4HoxhStUShcRkyDW1
LHJnt1equIfWhdDB2n0p9eEqzr/cYt3jC6Q4dQOaj2zZT+F1TynWDMLhMAO5y0v8fqAvAS0Dh0OC
a/2vgq5cTG3ivseDccQL7fzvFJctRcYctJqYI14Cv7mOznPBoKiyUKNHSh74Y42hLwCLfB7kVyLT
4Ag66C0Fc5qr1aREEvQ9pWVpOgh+Q4VcGaEiysf0YqjAJiMsIbHUEpcsDPQ7nssYhyXokKoIrtCR
k8c/S3xaHvDCZ7syJRz/XGN+vvyx+gqM4bDTtsXoQV2/2XtDwGEkD8nS4k2POXNYQax+Wrvhrvmj
xU3Zh5IBdRsq/bIfI/Dt3Xb+crppKmJl0inbNMrGnHmiYJU4EaTG7CvjDIsyFxElxPfHNJZQEyQj
yQTr5Z/oB4qYha7jyOACUmi7X9s7g6AW6XKBC1YJ7ZhMNhj5wuHbkw5KL7gJMW7hj+mYmGTOS62u
0EK6kGTKpoNucml4XzWXtiVAhzz1im38ydRC+jQbc3nRF2IDJtjv9gbmK5haKxeGsMY3R2LdY+s3
3d4CcGcXU59dYIBiGLbM4tLMpBf2LjtlaG/VSmalRedNRIrJR1GQyo7kijUzmQY/ASzZzwsJcnJr
DCCxMLLY6QuMWh7OwnvSr4C++W4/vfBEP1EC5u5VNG+q17TX5SP7CVoO3bhi8JeALR1qPpZ2yEIm
PHaHT6xSzHdlPp/SCGC3PZaQWTiIGsaf/TWHCaz+R6RhsL6OsOVD6mYdMTUb4aA6vm8GzH2Qou8w
3hA07Q/rLkjd7tI9sOOEifAN0VYF0UPTzlBmXgbTOTVV38KHFtdBsbsO2iD1944MESLkDsaQsX1f
MVKoAWcXRIIe0ZN6p1Qse7CuLsvRnRKJ80GaPObL3pptd7IabZ6XbXwYiKrZbuu39ryaGHQNcoAj
wdCoe5UsMCJVpvxNPKQj4j89FByDrS67XrUGdfGi/TSaQK6Sm24pY3N5qOhexb+vZlVFU+t5uJ+E
AuWvnQJB1vwV9tFg2v8T1Z0EKYQXCAI5u+J20Altyb/3IIBZYufiLPkrSo/DcXUosJLmX2b7+6aj
oEv0CM0nAz7d6HrsuP9WkkypZjh+spyiwkJ4dN3slKHTUEkA50NGfjXXxPkugQJAXXB0TKEfvAR5
E8/v8Mv59KCeowpptCT59KV5OnZJpaPI2BarMW+OyQCr1gjzy5s1fPcR8aN4K9OfelO6sHKaoB/q
zIHPZHD9OygNQ9hMmtt4bqyShMpeSlki1fH+qsfaFGJAF8seIDe4+PcYjPrj7hE2sO7RHgff773C
/XGdfeHKALfoVaIKcvj0cIz8FC8ZLtcizWjhFmWj+rYpD4K3AJjLUx1UEx29aVDWVWMpPnsTXoi+
xnLT4K9XOKFHqXTUnjkMju5pDfExvZuRnKznl6dSvSYbJkHFPfFkE8Gv7pq1lOLfPU+F3k4gNqvp
G2N+Wyh3I/Hv9qokvC3dye7UF7p4EooTU/iuJdnVMNqzeCus2vaahSkTS4rJHq1VDsVb4XOVbVRa
TR99+5tIET6WOMAhFk6Y6moQo/G7JAGHSd7bDRpb02smIhvYxdL1sPcPOOyun87LoSgNY1TMvXpK
9jPWvRnbQG+xUV2jmTRETTFoP63gaE158eneFQZDHluX3Z+AGnUMyljLWve5xcUFaqba7cCS9NdU
E0I9FXoLzghLKeH7yI4rl0vxVhNh3LerB1M7nYexf8+p9syvaV689zlo6+7H5jNtWPyXA+MDfnv9
unqFuHeehq4mI3tzDxQpgLTq2TU4v/GE7n0Y71pJ5IpqUSmPK8uBlFk70LiWmj4AC4y8M2HK7vyl
7WOKaJuuENPa9UxNaiZtCLgd/HAlY+Xj59ePz7itQ6VVFglisme7jbGJ4DsicXldHuvF+8TwQ9Ow
UVulqC79+DI+Mtt83BhTB/bNzsKk4Q79Q0Yl/1b40Pmki11pCb1Aozypu06/MLL64PsJq2hHJuHg
HpUDXEo3n6tYQXPvdSed09JZudgyIqIh6bQz8UMNjDIwm2iRBbVBYMz5+AFDnW63tYGbbW4G3Ai5
2j2KqGsk6/we/QSSqTl6PZZJZRKzqgW2BtJdd0C+AHavXejiVXRFCxJBI/p8MZz7fO6lbIl0pWLQ
kiQdu8xaprIQtv5Y2kowDah70MU7LElbnQjxGDg+m++ogTBtzm+gPuzvX6IJKJqYhfki0WYqWflx
irG0CGJL92wN/UOMpRIadmkMISnEa/tAZldAAxp/iNJrc1vBr7tOmr5dMbybsZXfcf+svLIba+cq
lP+tw1fvuNzB7UovEr2TIdHRrfqgBCgEaHALo+NSHpzOKMZONpFudpjSsv9EgYI2PFN7yZl4PWK3
EbRSLe++jGSMdI6x2thuMm/Zx77fAG8Tu+KU+Cqsi3r5G6DVdcY6IoQLnrzp8++OtCHdA2joQfL0
h59pFteJ1nIubFAVhFhq1aLSdkIhbllj16UsgxQaEvYxEeKu47uud57W2J0chKe4NmBFCmDtNb9z
6RyfaG8dI7fPTiMJHivoOFwVsOHxLivYGSfM1gx1xnlnOdUatp/wa3B2R1hmG2g8ySSmsJhf97/x
0kjCc59zWSLDgHvsYy0bzvj8v7p+Zx9GOm3DaGpHPgxJ9nMmMk1OYwUoM3OJ0EYJRhnMY1QMNDSN
eA64gvKbF6xjBTTn/6Kd/fdVd6HLBzevQSFjE0seuw9VUPqynosbFQIiGxCZ07XN9ZYdqSqfDENM
UV1By67wXgmWgHM6x8Em6pJx2NMBX466bM4PfTu7yBNk2mvRfarGqMd79VjYLW43ALiYkn8kLg/9
fjSfcIEL0Iifpchhh49fZ+szhOUJTNLuixoR346IuLVR5b9pZBDnHgfZoa0NMGiqfpYEb1JzS5gr
ya3gjEA95UweB+Q12onDcLSqIu8Km2zFBsihaHfqLCEd6N/EqeYCphhIXy6gly9SnB/jBjQSUnWe
ai8I9SjIRNDSQHtuT69yRmtd/GxW+clcU7pQ4nHuoXQN7MkjeP/j0zEuI+zG0NLMw6WeMY9N93dR
zs0D1aAWeTvnONpWiD4BDi1s/lYTf2DS8p4i3I0dPTJ5VCZylhnNeSORAq4MEpIRw/bxydsg1AQX
lbei93i6mDXWtKQjZGlLSJ76MXV5vrZTvwhiMTWdE/bO3LLtAjLZc11OvquJlJ4RWke7RhoRSnvV
ZLnUsGDz6rW5q3UfEqeSyjnppzPRh0VajdhOIBAuFcIFafqtHkIgBEA00+KX1vjtSrASMLfDX5Wm
+cYF7t8dZxPmScBMLzTB1cnkLXujkC08D3IXoHv+K48UaF6VQ9ZpfujjYR9sxd+QlKeKatkunvub
6DLNGUOS39B2IIMdZfDBJQhuyOgfOeFL5mxt3F0jS2GblogYvLOSdEm7dmjZhPYzLFzZuPYSRPzO
ktMN72Q7RAYTf57xCYTF8e66jElf7ogJkALbt9yC3ybJZr4hz5BerwohGeZDY3ylZF+wmL4/NHsM
7dvJ2/Lv3f0NsPFlxhk18ED6fSO8NaHxH93PoJitfRgxc79VrvtI244ungD/NikpscPtOo7b21hu
/uqV26MGc7N8ZpE/+mNQrhcYmBMie/ZOoV4nsrbcnlJLX5Z7ml8Os5V4tVcFYr8Y9ObOfVRzeE4d
oov6JuHo6xZolzGeznVsgQq9ZHkDnJTqDsSXWrZzqIOzJGSEEzcmMq511qqVZsIj2W5EHgBdpVw+
L8GJKPCac46moAIlYL1avKN7VloGfoQvZc6rkWvaUuQOdAmAPBDcAsUCfsrEBlQD/1M1Vi4EN25z
DN72EjwRNU1cl3+SSyauynvYfsC3TXLH3yPkDuqVW2YqxStxwf73NzmaHSLdlcaN9zpysF5u3fud
PgrLbXkQXEEQ6gjwWY/lB1gAHxQ6d5o/dw4hxO07NRRvpoomqnh7gvfCzUIufnVV5+V2FmruRQtF
TcokPNTnr3B4HbtdqkIHXGJocHeN6R+ODlD8VejeIaV+yfkLfmTxH4diaf5LxdD56rGgdWTPmfZm
m8FQ6ZAuM6kcR74oadPc+FeqO5g8DU7/eUHd/i+Tl/EEESt4S0nso1sr6QcZC3awsMvYp5tg/Djx
TK0gXNTbb6yIl9oG4XXWalmV1bImw+23LOhbXJ5ICdCgz7ZZji3t2ft089Gkt153uDZnMylJgcPl
aFMI6wF73SLhsfHKBV1AMIYuhz5fjSii4vbL3jH3QFRrZaiDrL3D+RCAtdcAP8uBit8vtBV9Sxgs
w/6NuIuKlr4OvphXRT2ZZpIMLnjykYR5WEC64BiQJ2WWmEfwF6NFz9fmUbAZrdgcrxay+nFw1H4Z
OMPk8AHi1x16RSboGAj5mRa+jntIT9lXWpicORPmZMjlcbuiBpP2AgXtjTA5HAJ/CxChVPiVYxOt
4or+MJhA2NK/GqbpAysMP5ps/j6SA38XYGIMuLexmBvvjsayRv9AQY2mg4dydJsOYYUZ+09zOabv
oJGpyTc6eQlLNf7syIg0TZ5btUXIcMuAiG7yhQHn/YlZqG5gbJ2nuwhquTdhdghcnWvoOTRkKofE
Xz5g0QKXA3QF0whFWURsPR6ESH0GnTr0F4fn1ETTPuI8oLkN+TLYtc5Zif99RTW+YppNeAS2AalL
XzBJlpjSwDjhzR2VK/5BUqcxVHk++zE5yVPtefaGHINH+jSS6gRTiPEL7w4GAsmfAdK3OCJroWiO
CcQKlx8qJ6pR93NJ21QN17HJWZKTilGKiLLNx85AerR2FL2YT7b3q5LxTYGuBNVNS4xIr0MsMRi3
3p2fGzMfEA2M5JN48VHCkw6w9/YU71KGy8KiWpYOA6KG1KkT7wllPWcJqNGtXHOCHh5/YiiWKkup
BTQdhfHqO1Mjo0alJXB23sgxgTArbNEyPhOpNM9aa0g5VpAzJqDjW1xFVWNAvG6rw7remY71VAFe
FPl8ulpMLMyTyFV4X3mOKakI0MlbcWEpku5bcWUany0OWM/5r1l/lcMz5HcYoGBN1VUGj0UM3bER
TDpNWEqf4aSxrqD67fpOk9G5UPsVLhwJGoRcFp1rpjymoptFB8OblGkSygLThwkUn+EHs5z4NaQ1
hMstlxB3f7pM7yu8T/Ehvlx6XfF3t+aVY2q+h53V5cSYF92BJLQabHWsDiHYe0Y0yky+56Ip23Nh
gWIZz7djkFjvQR5LCgiIJFA7JRUaQeJry7pjh5IWlCiutb0EgSxEb7q1+77xEA2t5FiXNDHeU9R/
Yfqi0pB7eF1LXQlrtqQXU0IFwqtPUtvIhykxekRhmqWohBr/oJvd8z/xRqGjEkncloqD8rYcxcvm
tW2rhNuqf4S4mXtpPGEoej2mnoPcRDON+s4e5uqOLph6dfF0GBtB4CB8tux2r4sqOKnxEk39H5bf
8AbycbjDNlKntj4vvf9aDQyFu4n6nE9nefuhEW9rCjxIjTCH8wLv6Y32EOiGC4lzTQRZHW7G2ysV
cPn9Cz5R2q7/VE2dacqJWA6P5Q5koP6fQI9rYHnVu+XKT3vv3ppLm1Ag8oRO6wPyzHhYsK7tOAY1
oh8mz4Xna9mn8Wm1OLwzuSIw1rjw8aEweQY2s756d2UGO6arxBHl6uJKhg08SavoH51d3FHjBNJW
1ygcnthINzm6p5YtAGBKo0yX7xEn1AVd8uIlnwwhI+pKatue9wl/HfCswCkQ7YEFnEEHy6ZKaDA4
Ls9xqZyZVwpxmnSNfgTrcCKcnp8tPRuGaJN/Cwtxo7EPFLoQpdjlcAUascEcCXUamWL6y9Ox62AK
H2iutFd4YZCXq3R6nqhUT8a9ycIehs02G21F83eR3d+mWfmYuDLe9c6l17kjt8Elyq3ftZorOTwt
7cO9YIu9ogWI+QseiENDyFtYk7wobIJmXMF6PskjpE/RdYbt9e/uPwyLnydvmhz4lj6BD/GT5uFS
rVupgiQvQL9Oze/R/jusw/cMzCddC+viQWO86djWGfSq4Y16GY7f9u6Ir0oamCJ2os06N1D3VzNu
gEAJEczshKzqImHwceHjWG05FrIzy0RU0gFas396aoUYba6rOiyRGQrhEeZjDc1YH5+JvJu3xMSD
NDj4EKGcmlj1V++ly+2Vz1FmOMLZMcYx9mCOjav022zJ03+BuoD0/1+nt8OvbeMEv/LdacoDEk+D
rwZ91ivexfD0Mx/zbD8BsMB0cs8Jp7vI4a/tcjC5b6mqZagoIvr8r32eNGkrFCZe6LUdR/H70Ooi
D4Th1iKF3kGXPk48I+1rjSknBsV9YXFwBR1GeAEbKe6PfOERspm7reAiY7FU0JmARMu7c3LDFbAa
3Frr6ZT6HPFvF2BkYu1JZkPnivSE09Wu8mZMwLMvsHkZo7nwy8+rXpvM8sVg+eY4MZX6Lnmi2qSH
40D9wDJiIIuST1wUMDOOqR1Q6UNv3SSMwtOFnic8A2JhOL8HtwvBUKd+MRpXuamzCccxOhHv8kDv
HoGR9no1iY5Mh4ioyv5S19SeErt0hQiQCX8GB1ta5Zpwf5a+Fy90vJGLxMHHbnByqzBfo2JNkGnj
wfhsPFf6M2wbjcQMHqg4oJsJOE4lX1SPFmDeVbw2hFkp/GFM5eI0AAlCDSrcKC87OCHkUeafYPTj
tCXDvHJY3WbZD3wM8U3lURICsXHKJVP3dvhNXfsEH9rkrHnMiyEIdXd0jWkp9maRoM6PVwhHgUgo
8ur28RNVeLq6o4PynrwdAadim6pTIWYY88mNQeg1iWGBFVOQPMlbNOmNx+wJsBliRq9gsRdtIeJb
EEx35MEhUvK4ZWXrnurowyF9yRDzXaxEH020TVJv6SV4qXadQwLp5vNxJWlfBAUgqhJoTIgsOOfP
0MTfKmKv8RYaZ1eIG6wSK0Mp0J6wqN59ZkIBhOeDm2Bnn6e4NO2A+BA3/qUsr+S8knkx91ucJ1iu
w+pUZgkrmrb8TCwj1mRjpMGkBKQA3/tilxMGcMPcUxUlMO59tby786iEkJa0f7xcNITpiPHgQRmI
RtUxLCgjIewglwnxqkuiw7SVLjH0oPMtcIriDZ7g9UV9+d0lrsYVRBBRVjn6KrtYziMFNn+Q8lMr
/iDXA1nKQb5W1vpS574fBBz+KgvvVbWXLznZOXgViyOqMukQ00ciWUSBBxinY1sgl/e4cIGTWSOA
y3k6pA/YxKkpUgzQNrr9rdGYTLzRpXvVOXr1Rmu7dwLpPml1aqM/G2cj/+qGB+0PZLGHY3ELAAjH
FSjvf/sS3VeeLV76LORwVZMZ4/txcW5NVc6hkmfMS8/Uj4ImpaM6VQziAxy3f32vC07M+TYwSpXx
f8GynGKwFFzl9B2sP5SHc1G+q85r01OHbA2+cxRQEXbS2rm7U69SdpaJkDnxEpIimZThejH9Rizr
CSr7oM5iB8bd/2offN6GB9emremJR28r0uRDpwDEH3Z10d5YHlEzYYZ3aCB6A1R+942pk5Y95BKz
OcUooDQZbyURbRWTyOetQMUKQKcAoPEbMjGlhMI6oDAJ8/FsCcreIjKqfpUuh5BoDEIjeiLKwX3X
pWmNtO3zuWpU8h+EozsT7BSM1NU6wWCl193jUKS9QcXhuJ1JoprA7Hvi6Wm1roB7CrNd/HyBfyG6
lBBdSxYT2HO/CoRS2DRCUCbuyTvWA4im+/1NpZ/+0o3Ny1qb21ZjZKSR6B8drNx6jdb/qgE2QH43
qPLt3wy1OL8EHZ5mqOaPCRcuKp+qktp83Sp8BN058L6feREoFbgOTEybRZrqRS8WSVnlm2jklnGB
VhOp64Hj1/d09Td/lVWPuFf1Jx9RtS/OLwaZlotwwJZmMnjUwafNuaP32tPDMr/svz6UKjRtuBlt
0ZyU3ZiCkXu87ra1qcOZ3+JGK7htGJBprrYnReNeFaTo8lxWHvIm/akfHKEQqFBm9MqKMC4LzA4O
xfY7iah/4AF4TQfwufsUVZN7k5oSr+Em4TbVkueZAiUg4ciyQiPMeHhgUOb7RihnzUS07NjF0aCG
TNzbXTGvC009H1Vid45hdiQtBfmFx7QQMfJPYs8+C8cxyl0RTSRWjFPQFkE+LcMTacuGbRBQaDoq
TRI4SSV0hOWqAkEmesRFWPsA5Ojj+xbZ0himS8ZGbn7UMvNpmsg2lNItzHTpdisNEBuwNt+OPXK1
QvgVzeytA2RqtOoWQPnnKlT3Og4w99ajfISE3t9SD5JDGjy/57rJH8NfvD9cbq/rSlZkTZRccUNL
r57mHNDtJ7NIzxNY9SicizBSlCFh78n+g88VWaR/+ZnJoUp4dbWXEdUpUsnLXf179PA7vULwdyN1
gA4zyuhs2kI5n+7YTe1xeLTCkCmhwBm87A6CrVBZj2Kxl+bQ/0WiZKiGnwiCAHN68H8nhUnW2+vX
RNLZ5dy7SWGIOtKITAP4rbOohrL5+g83QEMlcd2TQCptRAMtB6qcvLc8xzO0OAPMoJbo2VNcJO9s
Db1QYsgqmCweL/tN9uFJ8C5dLwJC6gTv+8CHv7Y4pTBRiKJhD0+6BP0Rh0gCR/EMyfW05BTUti1L
u/fGzaePifJuHzUTluaUeGMU9cBkN9o2tD9wwgn8eHPsDg8qZmR38WEg3tCzUysxo/PmIya8C/I7
Mhv1qkzmCTnH40V3Zp2EQNOQNggxzfUL35/bjls3A8gYk+OYaz6ouKwwqjauTGHhDkR9DcCtrpkA
3rQEaC/I3qDK31O0o/+BfkjWJVVfw1VNKaZ+TlqUuqWGs00frWQHJNhNi/KChveTIeJ02wakQnyQ
a+nXreuY80B4vShnodyEit+4w3g4W+dcHVtnZpVH7InOMTpsdOG+7SU3XXqYDJqc09SVIgC2xAzg
RRH4g7uM6LwL2wC30koi6pz39/rzzBbXGyhTbGteEHqOfXdNDb0ZYWv9EiBzGBUcKXhkDo6LxopO
GxFR0SGK3SNypm+nAZNCeri7fPhpa8VZDaaQ0Ernf73f+S1Sl6E0eZql8U26SyCef50m2V4BbpP+
OhQfL3AHJbL2qpUWvsU12nPMISJy/gmoc75ZddEtd7StGxQJZ9qwdMEGZQF8U0n74FO+/eIGH8mH
e9HETBFr9RYhk+NAeOlRnBhc0Kw5sNQnedSEb0uCaFxrRxyREsZwk6/6fF8FjjdIjXx0nQrb87NB
4EXnf/i5F15qjlek4DpO+I7BUXlF1JlicXwi3fCng2ynEg/P/85oOEQRMLPxCBivfhntL4h/HxgR
h7j+npigaz+iogoLty/vQFBSIVpJSgGJq6moDOl05bEZGAIXbaKIrB2m40lS3Du/qy18c30lsT9B
imt60067E6EWlpGqFpxkQhvFEOVJPGXdlbQdjCOz1zfG5nBZ/AxurhvuW5Sd8ps8t7HhvAISUuy0
X1o3JgWp2Uf9dgfm7Ch4x47zengje+6WuEuaijUSggPPRV1Er+RnL0QCmuisKrKqIxrapl6HAX0L
cLOY/3QC73a6vP3Al/2lh3Ea2chy/uw+8mt+HA9sXYbYBB+sYIS9EWapolK8kcg70ZTGrZmYdTlz
A6gTrYqMAaM8sr9ChLNvH9vp4Vih3CPhPd/Hj3Dj3JCkNvkHdSlen61+yX3qS+lkpoXPGUW4/gEL
OXZ0+A9Q3qmlnGvlhr7YYyB+24xtWxAoRiVMgfSpu/OU+POHUK7IDu/vVWq2MZeoiZNhwkrt8G36
ipCLh15POb+flgL/p/626K6O9L/9CEloSd9IOwx1d8gSSVsG9yozKSBL2CM6A4ntGns6BVmHh2bG
x0FGwBvV0l3+/MrZJfbZY5t95/NY5A53MXClhMrPg8/D+fKGs8ZwCZQgzo5YiogjEzLLy3vtLzYH
c1xOeYCGlCm8uhwnDn+Ky6d+LBjk0qV7nPppXRIoEe9PG6VNrOdb67ltgRRrw1H8ZENjeSj20/rK
442XoZmZa6qquR2BsAzWJu+TQQ2mo/b91RUEfnEqNLjRfT1rC8Vtw0riFfcwPzq6xuWia656m6Xn
hzMfOQYZ2LkmG8NL3xs423oSxrfui3C4bucPo0QJzpFWZAaTDjhtBuqbg7Ls6d+MmcktaYPo22j4
cRKvOrrHjYxo6G8KJ90zqvsQo8yXtwoy5XiaeRojntoQO4a9CPWQuFNdYJdEClDBwNwNgd+cvjnv
6duYO5wyfr8TfYlq3SgyZzOu8uUr6EiEBorjm0T2ALdhwGzTVgDlg5WWbSHYy+ObWSYDpswl2YD5
ReN8g/UywjT+nR1/xRwXcgdZD1hL77m2WLOJAehzVe2JsHgrpisld7kEBixzn16F7ziw6T/HhA5H
iYFu5q4eDRQTG4y4L/RFm49MdhIj+dSSvWK5+/JtruZpFJ7sfdmB5ZzAuIzUSyVK8qsAtqGvEaI9
F7V8a0SdpgGgvDUfu+fipaezPlplzWYtzIHN8FsPZRzuLUnIL4qQNTLtJPxO9tpz7BJTfo2OMXrE
8va8piNTMNkEht0V14gI1VVOveVG16UbsnQJJw9vDKpTvfd6bUtuH/McPraTZNK+fMHS2KFKqZsl
cYEJ+H8hAz8TKz8Bk/meUTj3chbBG3d8/t2hYBJ21lK07jW5r6+MHi3qh031s+zLG1UAXZJRRIu2
jiMJZ7S0m+o8DlMhMumcShuFSJNbXiC+/vAtcGSvzGZb9vIWh30oQIYWp2710XES9e467U5PbNsV
uE+OTxj2q3/OrdNw7swUQ1EZOMxGfqT+35fbPDePhajL+QZ/6/tgapaOpkEOxgHUamLYXaDPIIoO
9D5wySuv00a6ZwLkUGIL8w/I1dTpCyr8WIIXvCo5JH5qHzMyI8n/FieT5dm0FQd5DU+sMiICkrf8
MR5zbI3CIHjAqDwbjc7UpkuTq2mcCGVThPQSrRg0dRQfoXwHNV+RXZk8Vbr0kDgYRFLi2H4HtGxp
3Tr9hu4P9apGmG1aXYjMZVagXP2juNuiP9btwjRojkVTyyZg7C6kXIFWOZ8s6pphRehbt9SjI2wG
0DmKXocj5egl77DBUDtBlFwFCyVMJAWS5q+ymtLuMYKvtbv7kfYa4ruyA6ibPwU3bMdwCf9dAxCN
5Shb7JqJPBVcopMSAG3zWIBLGesQgwO+1uZVXs5Qf8Kb3ewin6GCiuRjbOCGsTM5QbQesct77cJt
mTwyQHSe2OR/c7JEkhjopqvmMkoToBBm4zAZuOxLeelrBxDr0Ueur0wJba/QSUpnSoxhf3/JegBG
Wz+IX6qy8k58PpF8kLGECMt30EHPOSGB7sQsWmeJ4kpeqiHScMoji0/v4LQPXLj541oPCffxZ6ZD
9hyQW2faaxGngx9Y+MD1jNbqWSpQ4s//CakIWg7e2IylMyj37B1bx4JZbXbsWu74yKYDh3IB0maa
eXtDPiT5XEhY7+YHfxHXVStZdlcpC7BoOjzS5vNEzA7pCu0omsDaYai/xAngnka/GU1gt0bmmgqa
nUIpL9Q/86n8G5M+1H1oW2zQk6f1rtsVCwHlVJdFI5qMZsh9K+5VaZ7oIrdTVvm5mX0/Se1mCQS+
r4rRTAcCcKZXVp/lgm/in9xxSuq4v+WEdudkHYepiI+NhxtLmF53TnFCD7EIhJRSlZ1FV5BEird3
jyXXUvoNGdLcEr6uffkimi8lOLQ1P+oZAMR4VooApeuGXn5crrWPj2Qp8P50+IKXzWai0ou22G3S
VQ7MVbxz8s+zRJNm1sOp73NH2V01xG+50xwvdOW5DmvXmdHpf68gkSHxovNSuE/L5NkKJ2c9vri/
gCzpopA731KImjH/drRZRLlWmh6zO4a+iSQwFvvlU9jBVcIljUbGs6dzJE2MSKJIvzqAVJ1tcvM+
9asxKT0mngvD4gwG8zjCmtR1Yj92+yMVNyVRA++Kmh/0juGvkdZSnw13oLS1UTa3pvzPoPSn8Cf5
9fI4YHhftdlohIZFAX6QFaPtoikI1sEP3VJ4v6FGJCYUaepU3VFCLUhUmqK9Kp0Z6+SYMvXAw77J
pfJENw/WeddeRlFpAPvQbE91wOJcMBcq1QSp94FqVvii42AMvfbICti3c/81/qCs6DJHV4juqmPm
k/fdvgmzNt60t+qR4DLCGy6B9Rfe0AwT3WjfTk1DQfwpsjOVEzr3Zu1HWvb7MiiYn/F10AcPWAER
ZGytSKlKDQ8OmXOJUcNYCrSqYNAXlwe82iHvNHsXEtRzudLRkt9JohDsA/TW5h/JX4QHQu4AZy1x
Nkjc64hUABB1eb8kUTddou81vA+vxZvS/ROWx7jKgMtj0ARGmLb3qqD5bHaRWJtmPztQ6mIcquO8
sTB7eNLhCQ16G923Hf1IX3hvhOfXypS46TqZNppDfVhrRMMKx9rQ0n+3Rn1Bn6nZP/3gWn3i8d7Y
vWpX5jolu0f6MgL65P29iiY8WTmE1niUuWwzE672mYFeCihVxzRhkPxAuj25jfHiN1LwNdL17T0O
y++qUtcVyISm++9dysdPYzmhOaIVglbqeEKMrK21fyk/C/sNKnEI6G/Dd/OuJADG5Ph6ITp210JO
hz3COqHrOXwZPAAcLXWPYHm9NxZP6n/Y/CdSwGDwfCaumhjymcxUyi6f2W+TYBOOgh45Ss/VYDEF
Yx0t8ik9EMUMAxlYX+IFHuG9gw9hMAnRdrt7nTVAh5vFaqo+fSI4CA3auAk/1VttoTeaj74mKo5u
0f5yfQ27C2eZ2iwPwItPjFEzr6tFLNBjuecE8MdgbV3fg9+e0LOTZplmkcqJd/V3/uIRMeUn+CSd
OdgYuBqE8ZMKWpVwMt9LrPqkZRbIZgmcosjRr1LoEdRDfzmHTK9HI816ilA6VxBiI9OrfWTa4aao
kJMLoASlows7BrIf09FwHrxOlwQWDtwFjLm4K4ILMnMxGJ1LKm2OfYYtlGo2QScjwCBpyJ/fei+C
CL420OBleNYoPy0dv19ixHwemutChV9eltPDRW/Zah41vhUe1g22Uyxdoaeobpqg7/wWAih6/DaD
jFJOOPDl1VyVXJOMaQKLjHAk4CnWSRRCr6M5swS46gX+p47X9qKexTVKE/WHDiKUhRb84YQLjwlz
D69ifmgYsRpUq11lmsnLlp0cxO93B5t154R9VyPdxScMDdylnbRpjw2vjqXwoLuNwcW9uWHZk8G4
STcgUBYOYCaJiUhMPETM1AiA9/XJ+S81Xp469lXk+uASgILbOOuWL2r6XjMTOhuVboKH4eCUmpZl
kB1pnUDUh8j1vvCcUx14teBGMAO9BoHDiBUsZhm+pWwRmESKL7wYKO5MYsVs9P55AIZ4Dh4T9aDA
YAJiP9kVNfsjdnYuOI4K0EcsOR+FXF9f8HM+EKICIzIo3PU2H1Ls6JETyaaZEteI72+XZ69xBV1F
rYLe0ZDpBQuzFhomI/+jJtV9eZkXWCefNh4U/0LHq9unJoXvzFRmShwYLVOXDu6xJStSsZcMsZGj
72tR0OIPlaCKPRccnlq0KsJv7SfBmZxgZfS7RaDnATZLSLDtswz/Irtva3QzWrqfy82YjqM6bVPg
H1EFPXifZfB2bO2VWzR3RUk6n4GYjnLN1Rfb+bP1F1vsJ15Wn19XCCpU1oBwCRYfbbQhFDokDeIT
sZCwMEVUa4GhpJ9Cmt7uHYCoNC6JH9nnsG03aHf5ONi4vsFOPd3ZVdCmTaR+F6smNhjty9yObIEj
YTW0DQQrn6EqB7DlywCejqLaYGzS7bg2xCr1riI1QSP9C/T+hu03JQcre68OgH06Z/L/+G6Vki6T
0TdUMX1avQ3TwShm4zWqbwLqLUXaNN5dNATBDFMcaFedspR5m7X+c24b50YE1+tdh/Ek52SW7IxF
mMVCOFA1UfzF0lUlJ3wln8AY+2H8pzA9lXa8RmJD3UP1cNLjs39U5xG8sA3TWRGHLCWIbyDh9W4k
gAGscTyYd8k8+AM4HNZlewiVpp1SyPm3TarmgFFrawA19SMpDOC7vE/lOKO/2DFXV+4lIWf3glrc
Pm+RDpQ8BjuL4vTi57vbX6Ouoqz9/vvtzVJY3H7nhaNvpyMTF8RNfQsgiO3fYWT1YyyecaPMcpjz
pMjj+EF+iwVhnRBVXiPX1YxD9uaOl0G275cVBz7Vs9pHSzxJlkPAxtEe0GgRvZbaBMeuQSJwXkjE
5F0gni0lQOu39qX5DYC9AnG1tABkPhgBd+Bx8l97btgriCnJ5d4lOKr9+8OucssS1oGL9mCY4STF
Kd7616R/hoWv4fRZNueFGdL8lqenl25jipzzYUwWPnBEZHI2rdaYGu29/9FFvBgYzIjhRgqAG10F
AGRl1Y/DPMCVRofIN2cDemjT1FD3E3SQt85Xdjh0A9TctMqWfqZJePt++zExvrG8sio5EbdXbsAm
f7uemUTD6zFfbtF88skFho3ZDinvxqIunVRoro3LvrHYLHgIT7XbXua49X3EaY/krLaDhOsgYnXF
YRBLaiVA4LkwMLRjixkb/q6ZfPzQFk+k8vawyhnTc/kAmGqy2wAhyfwlisqynX68K3GNsUoaMO6b
2lEgLt6ZINexkO2k9d28hg1v5HM4q0Kuhj4UnOa+tqD8STWsqaNXGTnh27VWOdrhtHv+eQ9wtTGq
+pMlCQ7f13XWnjmL++l+2/GJz3Uct8djR7saUET85rVNm79dxLdedySs6yuR7gBAIckCzWTC/7KT
i7SxTO8AKCz8DycWrY0fRDmBcxdU0TYFUWyuhZ1s1x6JGALMURl1/NnDKleMTH/zqh0K1s4VktO/
sZ6KZVCJ4lqAJE/RoaRDocVWqNMeLR9GOmZkNuSvQx0xQ8+Rie6Atxlzs6Sii0/lCJTfhuk7+Q0d
YoAPtHS6xEO/bxhVxgM/5ZlNFsBxIH9k746oYU77wYuFXtFIVXT+DG33rf3YQ59/Zp1/M74BWmji
De6kbdceSFnCHVJXebL+Su0d+I9dwZYPD3axK4g87IhYMfFPUSDhotcKc81MKYlMP385VMF2mJEs
dQFXniwWiNZbfxkcfsWGCJun1lXObz1xLJ3fGB9tYOJ8STy/sJ6wKU0rgwz4yYGAiDCW1JG8biDj
x6D8szjFn5yt4feIgstWSniXWuIyhVK2e0KGIOY1PCpO6qzS4PwGFvDMzvTXIomckfRw2veJGzg9
8pGwqPMPRCIQIqb5n/nIu3OIl8U3Sq9bZDA5Repw1itvSmhzfqmx0b4Kdc6Fd8MgMjsGJkOy/641
wH1GMbc6TJjoj4TA34fQaqBk2LM1rlX4iwwC59MS3srBdKaJOlw5LKatdoMxYO8Q/FF0hcU6lB8y
IUo53yMF1lA6HJdrJ5IZoW/YwJPtLtTCc4+pj6kq0itH8yHNQsGxJi+gBAxY6sYgt3hVSq/NSD9o
c/c8ChGqruI9mOOyDQwbBFR7lO4EbLW53R0uwMxZ3ATtEWtKPVEgQc/ekoOnFhCXykoRGPhXKEaF
V+bU2CW1mrPZ7AAQLvnycIZQqJaSFn/B0wbb0o75889X9b5hjfpFooQ3BpF/jIMN3Vx8YG0kjuGi
6ENLkdn4s/Bmtf6YFuH6oHTStr8xCNOFiwAFwQUcqL2aohaYyVYVT06i2IdhR0IHbQrJGzHX4Fk0
Rpi1UNR3v/EUOLlHWFzIJMwxWP+xLI6UiDp3DP4dLcBfwJiF8AijsVQ7ia2aYnxH9t1ChGXmTak3
hID8VRDhqQunrwPeD5jqA/DZokjk0hhILs0PzZiZkHAMvN7KOeq+LUcMOaPyGSUsKu+ODi5VSt5N
I/yr0hX9FIu/dKMl+Vt38p4qE/O80nhL2ynxwU+CPMYYzm0jJhvtuX9gEUsyT4v5bp4HjfN5+Ytz
F73mrer1nkDjuDzcZsgzQZE6U4N02Y1JYyS+0gaAwLvACeZUakrkY96C70TowlS6zWWCvakRCUXK
rDo6hIBUwSvN7EzZyqHj/VqbT9nNr8c0JrDnaRliAagxi0pr6hhvYUHms9iqH0ztZWLkT8As4VPJ
pIU/O2sRZHiOo6l6mqEV//SOXKu62IEwIigQBhnHL8lhhto+DBGa2RB4OJQqdoviKwK4D0hA/9B5
0sVr31LwhYxKOZsf0k8qcTolP/veE80kcX6tkQZFet0j10K7FlaIq4QLqTHnortpAm8op+MrTP54
Evxe38Iu0y71Af3Kh1HxPzS+3sv2WkC0ZvsdvdtmaoPusTRQQUwtNKkKWLKh+Z0KUyrjHk/KqgZq
89JrnL7zhzJoHErL19WEnVe1k/Jv+Mn5ZA+qimzRqeuo7X4msogAVy8z/fr8xusfwFQ/QhfAfdRu
d4TmzZmL2s1zpp3AJXIgK8HoM/ylicIFYiRJXOC4ez0H5W/Tjtcyh7IFm4QXWvSS+ktFR1i7brYD
XO95lU9PZUEIIGg8OS4B1fv/728PoJBYB9y5bt2GuIgBJZS/RcBQ6uTUhtnZz3YxNZCqWz4Ze4nW
6c/JbL5U+FSG7dgWTc2DGtDKYy7yPMCiPeXNtu/oUWgSjTBPH54sYavA91k37+h7S/sBk9v9O2tm
fYg/tdGUfQDCSUf5k88lwJNVU5eBfSIxHSkBoRJzy4masxEHWbFtZrvxdhd44k/IFMPt40sIxN5n
DZGrnseJB42G0OLhzoCG6JIe6tBgGsB3CTl2+2NGusaXu8R72qN2RaFJggN3F3zr0Jfd43EsR1xC
UcLgvmjXGf8vhUqiWkuCX2vpLAMiFXFUH3Fclk8tA5qxCPECEBYjsCt3LI9nR5PbObym4ilyf73O
G2G47491IWZZfWan0nAAooceZ+bgxpSFWrZeC3hEqRMlVTZsJln+AFbDRwuc451EXMdKxGCcX007
AfH0aKuy+kk4ZH5F60wnovcpYbsqw678oVBSdXWGjYX3msXAwILoboZRkXX3T9dcT07iTbfTgdKi
xSEedmTEqrIwmJJtt65HwVSlDVk9iVnSu4NkQfu8OAnRq54W67XBKPIZxEEFKcGjVOfBgU705afM
lMS5yhSsqRTSNwOL0fmYf8ta/Ud/WbG3SOz9KHc/YoReDjGwZidsboRF5QcG681O3beg+QMPdgeh
HNEnaJ9OgONk0jMWIM05uCrJyf6Gygqn2XZKSylv+0p/TFwlsT0Ci2+OoDCYGeIrsYcqgk0D+HJR
9kXXViQ7sndLsUv1jjw4rt0eTxVAhSAAlMQ4g+e0ZzxU3AbmePDZa6ReCH6KBu0Pshx4j47Ngosp
zJ28m9Bc+U0uNJCSFjBJ217OxcAslE/FdWerWyQbzpPlNQArK4Muw1JdRQ3eBeI0A0WNRTkbx8si
6jrc6WxQ6g8vrRsCngqBkHJjNWlNBpo63h+SmF2v4OYiduIoNQYadgPrL2Rjo+ap1Pn8Nq7eTi3s
VUrLqv8SWYY0mHjDlYXXBCwy0+CPXZYo8VLI/zIzf/jxdnUfdx+diQqo29ebnRCMhCHuCHuVsU3J
bFsXENAFxDozd+0jUI39gCJ2WOAVn1wyuTcao0vrG6bjxW48KrKkmwCaRF900bPRxmp/iMQx6Apg
BuSmC06uTSRZgeoWPuUDB7HLoyPAkNF39itVrex0ClOM8/J5kDa7BLa6iclrTw3SsgppHHzeRcy7
k+CFGGR2sOd/AbeNZXlk95kDj40ooRuv+xL8MV9ElVT5JWKi9AG/zkFNz8gyEBI/J5PJ3C4SAXwX
5Hg1KplQQIqKEmZgjB+zUqTFGb2ftcnfsHGOlcix0rgytfGvLZw+SSw8+9PLrZ8nYkq7xTuLRykb
wsZtit3qt9Y7s0s91fvGZgEebVQu9WqbxV+tRiaIanJmMGrUc5wKkCkXhfLRfERu1ybHEm2fscLA
+yqKUqUyaHCHpGIpnhqo0EJIxKOF7V01nFF+9G3QfFo+oDaY9axeaR9MYpX/5UwXu+BoWJTZSDHd
yZpHQbBDZU4mDyGyQyis7wInYTUF6BFD7eKHgL1Q4ojzMCgdeUS2i/NncUyFxgt0sv23DhR1PIhw
B+JajzpMjScJCyon8j8uMIJq6WE1eKLb/eYioby3qCSyOTU54VbQ0p9QJOTYHuWtJ4JdXzbyrfra
uAY0pqqHsAq/wLTKiR815CPvI6tywiiu0VzSOxHIW6RjoEz/4siFNnHeVfEUwiLk5bti5N9lx242
UU96C7SrSHcXvp3zsinqQbV9SZ2Vp1JHxKmN4pe7lUtV+dBiCd2wrjyhmL+JEVHydga6DsEgoXdg
2O+WlnEiE5zVUOUQKnwzEANynb0DeKBKZa/GQVF9cBTdOJELDdBIHEu1uqRLOY+atGYgxjTlaQxN
FIscyqivS1mc4W1q3s1UbK2VAZXMR7liG9lSkPlxYLTm2sE1D7n3bK3sSHrOza1stPjUFA3KDt25
4V7RniVleEt07lcid3o97+ghp9lGe/heLQCTA/rbhri9Fz2YtV2EmEt641pQjPs9RNfnUfTeY9c0
n+UUOLnPXripnwIM7bAL8RhrcHzgjjDN4uemt7eLuLVQlfAkIaaQuKAEB34d6tpkoBHVvGzJo+Cw
RvdyvEnjSeaXJmFPQycnK7FEKMQo3dmXZNlBezMiZKJq0W7jLgbI10/Zu2Qwh66nZZuFkLO0V4wI
LTcsaaJcDMRrZ8M2z+mJ2YyypKgi3xm/ew6/DTFXeT/d3C5Y6p4kmtEd4qjRQbIA7WEargZb9G2g
YYghQBe9Krr06/lkraauiz55LkhQN9PYTIlhZwvDY+R1ZyXsZ0HAe6QnK3gT/PCgjvGdqXZtmS9f
1zZBDkiLlcljEi4SlmzyHNnZ/7oUFeJlbR+Gsi07+wUpsaMGUjyDZQyCfoP3IAVAJMAZcZc6FBV6
97lf7RV1bmBjTNVmcgw/+imazRnTrazx1Dx3kdKNUUDGlUuKB/YLnm6jllKgcYdYzUXMuGIsynm/
Ef/r5fXcPm19LwFp+d8C0UFJDltyMGBpki8qrdWCieqHRCjsetz+jUIML3DZQJL1/fFSIAQ+xOin
B4POwu2ohZC42iJxThWebOGxz5Re+SOqPHAPlAL2Mb3gWSNZ5GwVIxjuKJaTfLIKMMVluj65Yqx5
rf2CxdMkWI494c+VznI6D4uLgOSWBizijYagmG4+FOxW/NqwRcH5vxh7BK+I277EIIXLfh2FY12o
ev4P8llcZMo86ouoCX4BC2NR3FBUrV6ef/bp79Mr/3cnQjshDkuZ8n+LlLII5WuOm0aIfh40AgVh
n0oTiqYYaY82QIgyayb/3JOOEBlFJE0hxjYX/p7javEkrWzi6VfIZ62Qka4PLqo+/rNVmCUGLDAJ
EWad6Kg6xcepqg7bsKoqQiHe2hLRaA4VoS8NFdoumfAa5jXfebbB15gCkraa451r1IQSh8/EznQJ
iJBW+Lgus5+eVmjIEOjZIgILwlf2ioppqac1KhOvUOHnkL98+jo5QI11m1anPeZS3Za5w0EKGpH9
0oPNtrgMshry92KHLlw21IVWzWhZl5n9IgbjixcsmY5oMP01JMCl8se45S1a+AgWtCZmNi0CK9nA
iZu/AqUR7wpujPIrU3MmkD0KNCJk47pACIEkOcZAx87m14B/18yL8v2+vQImIuiBXm5DjYw/dBve
PNin1wLGa+GduujX21mwhBHqHtKWlgNYMiKkCk8jm5CEnmgI+LpJ/uhAaGnEyKyHznp9+OgY+9/B
/zt87l9ek1KtjWLZU/vNn56rKKZWWG89XB4lIOo2tFmXHjxmhRTLEFz7gLUYjxp3bzeTzacokkss
SaxKEZaF5LdEbc2PyoXT7SIn5fbhPfnkZUL/Y2l0FkBWj5XT3YAo3/OS9sABVxG15uIWXyZOD5al
SBlPxPloAKC8FLQQtdVKsj7jOxXmUiHPss+AgCb/lzBDgVkVp6vEuO1UefLn13Shxd8sK4zGNepM
Zn084ybXD7t1nxkFcKhJBwXjJi76gTm3ZRgoGrjEw0xvUQkgvoYNKp//HP8l/Vd+TdlJRJ5jazxr
/OvYluqCN0zgt2Y51ZBT6h6m9+sdDhsxKGw3qB9/vjH04McUmHFCVfF0LnQ/U2iW1BCPBu8n9Xow
70m6TnB1kAPR0LndFaH8gGwEYfIn2ALYlR7Ti7YFT2qhyWU7szAzyi/O0HhKvk3M4IvsC0xwqQn8
yrpwQWTGLzowa4wrkBV3YXa0tmFKoqWmazIMmPLnRReoOzeCXdUUDL62x6cmNaAwrntAEv+rAgpO
NEOzDtP5czVEXLCdBD3cYeORqhTkpC6aSteFoNGgAj3J6Bp/VJyRVfmzHIzwvO4/RcCKDmrxsqIa
Hb6k3jVhIUxslRvjk7Nf2LjmCWhZbRRUhw9abaRboOK4wkAWKfY1HcK4CJmausacjF+McQPclrYu
yePobz7kqJ3NrtHlcs4PFC8GmprUexmJ7kJKIUaIhc0ad7yZsgUeNm94nek8V6cBBOl3QeEW6odr
MIzG/HkVqaiVhK+fJf8nPQ3Iu8DCTFqwx+d7FyxeNn/XTsLotVm2QeO7QfRIrugALOeIEjPNq8F1
LDiTGYaGGdy8+k/UvE0OnNyoEiUU/Kg8d1zv4WatAPQZizB/nmqIwxGQo7sHDBBBPg5pa7k9uQoX
FhLAaJymW11QMr3CStpFM+JTpliPkROpZzQFrUm+K4QWMD+FwYe1JIiOR6RxpMsBwcSDMyWg2X72
aUQGgZBugAxmASRp5Rbq9FtulRV0GYdVKV4hHQwDAizykdinSGRq0E4vZvAJpiXKDOOZbIYtPoW3
ktpvUqBrf950tYrJcipNjYYYrTAzj0XGcl0tJTdk8XtWXslg+Rnd9BoHXdnlIbAkAel/LXzIYT6n
KQMDGvQKz+8VLgP9WYrZ+i+CGnBIzA3VdDwB0Rx10v3RMaCB1x0Qat/PTfsgGj6hks7K/YXrqAkC
e6bSeTkAWxMFP6B342HAgTQIZVqs791RJH4fHOWbis3AerxxZR1bJalqOauIAkMt2uo8cRMAJaLk
SF5Y/FdQgCprXWEdfbdAI4pJYQR8DTjhv7hhBSdHY5Po2RTxRX14e/fhTnulnppeFFk1TVqJ7BEB
8ThBpG9cuQ2NndgVIYBRvivssqYSILBSIrwvxpItGR105VvyhjiHoICreuUO1pkiFXQegQdHJe4U
8TX/U1AuyTCKjTF0Pd4MxDrLSGrlMAtJyHmJ4j7X4BohMcIDdhf+qVFiS2Kb3TaZAmdz7OfcJ6Gz
ZiNH0O6V/e00txzkPkTN/NeDQt1EIyKHd3o0s8B0My3+0D4tD7qTw2tYp+KQtNFZoII1Xl2XOj6C
B4EY7ROjH5xqwnY30RpUaRx17A+IzJPg6HDuaxQ1e11VQTyA0YSP7zi6tgX+42oB4S39eco7Hx3n
ByhQRraeql6ls9b9ijmt8adB0zzNEPDRM0QAToPAd0C/YRZhPMl3qbvTyBWqX19SQX+xVi56z2AZ
pW4RN95nZaazIbz8qFhUEhehSGEC22ZAW9o8eDKih5kn3IYKYh04Dyi7x3gh8BcFhDSWqV4NXBIS
o7MxLmAn/Vz/XGiXgvHhi2H6XpkWHtDXMhTwD2kdBeCCAviF2V3+z9djI9D3r/6kWD4edcoMZ33U
DQEJpLop4+z7m/7TgpFTzyBCE3omBtKCcEEW9h4qVeg7QRbcWYJdMjT9fLIu4RsTC31oS3pLTsJt
hGUKtdBnRPWiL6Qz7X6jcPj/26GygBMrpOzS7Sb1uhsis2ErfENLeo/Cgb2qQhsa7j09MLC9Y1sg
yXZoc/ry0wgaFAEGKvlP6KFbFYFnyrW6Xdr/7tVeckjY8yju8cfEyrCO0ThABlMxjA0DCS2mBYd6
XPKWY542XCjJf/imcdKlwlQaMeQzrx7mLrnQI14e2cVESSXVNTI7NHTm6oZxMNR3RJQxYcINwgfW
lbhEhX7yO3ST0I/csAMGw0PPbIEWHFT8a2lZlDka/Jhb4+lwddE5St6+M11xS4r7c5XjUvvzmeWP
ApCJ+/s495xx24gcZWBI5eanLOOsQJ4vJeauJxY2mbSOga1EraqPJ4kvtzGmMBtMpVkQIIGedHx7
Ipc+QnX05AYI+6L6n07QrL3KbcXZnjJxIl/4PCBEmnAJhk7VQ/vvEYQ13gqMhQu8oRclPRZKiVlp
FIzqisIFLT9JDQ98Pa6WU5F9YQQV1uQrXmBirxP4XrXkTNqu+U+vRxWObMAogK/RlrMnTm3lAdg7
Ek+i+AVjxhCkjtR1tk0v6tuvg8JOeEhwfVCTgk7a40LeFtT1vJil3bpHov6QMRBFQCnt+kLBhEtK
fjm67RkfAlmx49dwOMEGTxyhXgjNfAZ8e+FUpEsfXfvl0JwgJ9uQ4wQpTUu+GIG79cybXVbKSlDS
Qu/px+1U861mNtd7DCOnCl9brTp2p/nbR29/tjIMhUzXenBA7h0ITVWxavPwYl3+izeI6ZZ/gQmB
tRlk3Gx9Y6ZQIXgCAC3f2FkhoSUZXBsXD5osllIaXGx1lyw+Vsz0qNocC0qHoOIm/MBLMnJAmZHI
PCBnExTtWq/wEzeKz104Kgo1/aia2h6daSTNg1CaTTMVIN2apXKQKcvynT4JDIf2M10myRKMcOg9
PBSwqzXfYuCt2ZY/o0PbalQ5NsNXKpzXJYC+LTjSzQKwmhWsGK/Vd0FjutBjkGNjTgCKY/ozAadh
00t+0uHP99O45aWW8UxD+RoHw7KBNZsHQcjvduVJWinhr/wid/iHBinhs0j9o9OLOhBZu2U1dhf1
imMGmZxir1RhlRGE7JMTkAmh7UoWHA5NNRSCSPARXDZf8Sh/zHtLFWkv95mD9fgUo2pIG2DFw7X9
OrjeGqPi+FhEF1oBu3zxp4YGsBZ7ezV0oS47WTuzXhZYqH4deMozrJCXMNLEsdqDAlJBokBBZT+O
7MJASM3CW5mKfp9+vvgqgsQhvMoqoGi6AUDFu5xocjGSQGicuizStGykkss/kh4KAr4jMWl40jP+
eQ5dRDtDkAAyyMcHh7XvIupEgbLzpgTj5jBqsvHRJ7Vg+8LLo6DsEdqTJ+696xcY1//Cpw30OlMu
n4DdgYDmxT41JdtVPaxhyTcQQkrW4LzKfywF+oxwoBeG1j8AeqOQNp9dJX9jnx1nBORBVZg1vPhl
6DgRBY64JZ3rs7OzQGVfgiJVwoZ0yUnIV0CTSsSRAuiYD4VhYZPhSRH562Vqs6eHdR/vwvBUJ/04
lEcUkmuDHi46x+2v9YBCdi2q/G97lCEDfRhjDBCX51Ek0Nsr8uLqoNiKTh9N6Zhv//71WKmW2bLr
A0y7GhVOHMYAdx/Uv1DBGichU0rJFbz52BQJkQ+fT54ZH7pC4ShS3AExIJVHhkGX2GJuRDUnsF6K
MlYPsfM+TH/Dn1EQ06evoe57EIjwXSxDtmI86glIHSvVYcHUueOG9aekw401GWRBCBOHwLaHgxjz
fUYgH8pVZVUIO2XL5/bEu/GrVq2TNt5MqwnKyhHXgERwOETMcNwnpZnbBdx7vYz24zlRezoeVNuX
6uFaxv8GzVbmMuLgvf2SVbTs+7MxwQ3Uyii9B4kfxemjfKeTNqylG+LCu0iqkkftjXEKjHUe4naB
Nkq4hHERcN+0npexGzBx1YgUQyNeN8jVIXNHrtMSQSCkeS08XH09/8EFCkee5G+/+ctxtMzLZIF/
qw6Wuqs9m9YwMXoutu5XLtdNVWZrFSHtq5aJpb5tdlSr2sUZlNlJcTNjNoavRKM4OVKD8O5A3a77
U0vsk6DY0Fiu3EcU7a9QHApDFUhlk14SYUqAliknY0td9zSOs3xjuaOPV1ue/gd8wDujQMy+EpYh
dDEyvJCR0uDMX4bGsJHS0ibVBWNCuxLNQiMpjvgfzXf5BAZtTl0/h+TwwBR8XorN7djBoK+EQ8c7
dYYlhIX7GwPR0B9sS8Neug/oyuc2wjPBLZIJWckrgYjcDGkh4IjZ7DOofJMKL39aDOm+paIeWpGl
bBQRO44ImXMkPCJ24EsW+6e+pZk6aYdOQp5nHlbimjVb1nM/Yfsew3jODphIlgqySud7/ZtZ2UMd
/5xkvCJWOnIRyMgvPbQGno0POb10HZlUdEeuyFV5XnLJSoXSEeuvdCc9w0kiDI9+906NmAab9CgJ
PRNY42ki5SzchC8BVgdpzEvmnPCuk1L/A7E2kdN+4AbnrK7GWts2p4b6y4v02pad86noppmTc/ut
lj4e2qXg+Tr+PDvdQ6VQclPzMDEPfdDSIhX7ykfT/EXEu/z+fJuSBEvUVpA8oT90UtfuuGG8//Ln
XXNhnnvucr/l5Pq7IpXpbe6S+lLUG1W2izpVDEjCNUJMnRrROsmTZCZkJshEqIbcvvgyKLbvWCWN
DAboqzfH0E6FZYfo4m+Y6zceJs2AI65nd/VBbtHCuTi0jf3Ra7vEU66Vfl4ZR8dQKTfbEilWBVns
ilyD7Hw33EDoHX57OQtfyY2p0eg2aKrbJSyk7aW4axBuI2WGyg9wmInnS3TcypbHifnIiJhV3x28
erDXI/bIyZkGbmZXlqj7J4bMGNIH+1USQCROIaccaRvumbWmBs9mqHcMweiXwmK3PQw1o8mUpwix
x0eOgOkwbodUsy6247YyTSO9S0e0y5kK9a+w+i8olTAZWbNRei6HqE+qkelJTXuXGj5S6kiwiUol
RlPZKyQ+OImZpOaRoxuGKTufsRJHb9sEJ2VZl60iByve6TgdXfM/eWcPdc6HA0FAGLcXnX/MvcQB
gLUO+mu3F6YH4cOR/Sho0mU3fDFwttBYDiD0X9s3T+zb1+L0rp+b+4lxfSL4lwXWPHtigNprX4fZ
BtYErstAu8ZKfofb4GmtSS0Qwxi6+waMPuCG55WLeQPqeudE6HcLtQMXxMzxiHFtkCVNS0MgCn4Y
Ntltur99BJ2FNMdaxNyN++ulCgjY30zFK+tpBb/CF8jwU1sTJxYybB9Bx/FYiGW41x8jMJGtwS5U
OVl5D0pBNXPPNXxlUoemuN95GxacRR4rurmbeomkM2gLdg3huAwJslRS1t0exzUvjxcuY41Z6kfC
+gna1NzvCFLk+Az1mAziYtbmOqbgMtqQ4J4/2tuIOISdmc6459AjBAXBxZVqMUnguboPPohsHcJd
Z4cpsoERxQs2KNEE3sECuBRftcHQJ6IYd+QlGDcIfr89FXKG9EJw4Ryj5hnwt+7xgcP6rcxJfvIs
cSNjAwrNghOen7zfH2u1XCfcdscd9QmUwMJrCHfHusMXmyjkw15ywNyqGTS13PqOIqVEYnlX4BnC
eHYSh6Hie2EEMnqlLcIefbvCliRBBvNad6EEAxoN5lW8M84CxEGt5diqSt9z1oJv8KTTzMWsXZ2Z
PbxqJUEZBk2nfEwRtGxOK3OG+kr/YzoaW8uRtYMaWozwlGl7MrKifRnfT5ecNbh4aHCwinYY8I/g
NxTHP/zcujnHnOPDVZNjDpNFIdPhYUX3k48+NwlK/TPMCu1oWz2ltlR6ho797pxw5IG8W7KFXxm8
cHqVxkon/LRvHAVDzH/doCTnZMNLrkNILFW06GGZzFfuh63Ha+AvQPhCJ2wV1flmX+KD9ZQlOHET
l0uD6QHc66njJmuHcxrXfKlu03amwntwNT8SnCkrzIz6+1Ym1TStgvLqJAA8ifd3YOfUI7nPuMvy
osQ26TngT49B/YssTU+kgTkzvFhUJ1OZn1ApYX5Iv01qi+3v1+7BWTf/1+DVRDRLWRW+b/ok3iaz
4/K0Pxfo8hO7CdF4QXGOuD11sCvu1oihxrR1PXuvdmtkvHkoM9gRIj2BTbrjC3THW1FiFSL1To+7
1PEZRmsCmmJrSGi2oicUUYYjCxcRU5UBzqDA9shLALDaogKzkjcfj3slVz28KD+62DMTkm7ACZNr
UJnakBOceux5GIyn8nd3kFTPWVVnvTtnH9jY5Xyo9gbP+9wysDZ4JaMdTCJvfCY42f/M9hkCmo4W
xBTInz7xSaDPGWJJwM7/Km+zDKX25rmC+lQaIL6aWOwd9p50JQWp8MLN7dB9eaSVY2xlH08DWfTq
nmCMLcvzYxIdIbPHR782TFrO+M4kC+fRqYwTT2vwvUm4WIwkYSAnt5s5gqgd5iTNY1NWi99M3lC9
0lPP44eLBzjWH3s2kWndnCL+VRjVFXveYvs3FFl0GKmNcoJR7sZ4KDtMfbHIkO0Jkw0a1rmzWdLG
N/1lkprWPWjYEVQ5wLFexEClbmnxHxm+k/EbtvwtD0+hpNBIP5/O70zotFBThxxakqFmhEQBJo3s
hyO6SMQLFKizdYz5IZOj7TMv86eTlOmWDI/N81cPfOpHqPnCch3z+lmjqq/3r1lpQqDYaPh23zWB
ua1adwxpegEL5Zk+4veALGT7U3QDoaCiAFmwcRKgSNWKqK9y3b1cuRDhFp1kfoiVfmhliIweQpbq
OwpuYz3oNEiba7p68ExRWQU4oJaXwH65AXXm1MSMBBJS90g2lKtyNdEHUl9TuPhWh0FLIX7zUalp
+s5cmc6rOzkRtqE32KhAfWL4ZrCdk/1O0wTCf3Ao5LIB4wIzbHve9zxm/4SGW2moK5FYioZxtl++
481FR4GnbT9WUZq5Qln3Lr71HVKbJ31khuh64xY+5lwpYF8jHYSDebESD76UzmDmPOB4JR/OKIyf
rlwC2DzxG8v0fIEmwNbxI4uVFbB2xpis/wHKA5jPr2y/g/3MHGl3Ww4b0SPnbKpl0VMa9cuHAES2
vUKl26dQ/XUPILowp7DMevkSNJL15kZZPin/Jo9OVRBV6L7ay8QMJ18cS5Zo3S8BfooTFW6iWYbr
OoRcCiA+1/s6uRrhwY6udsu2S9+Z43rfrrdkqNCuWAj+EBdrz1jxYfScRhPoiXFS4LqNHBhg/LAa
Wtl83g4CZtO6Kusf8t6CUkWSADN2NyffIGmJWniL5k8nNukLp/t32jbzOy4ON5fRCkymxLSsR8v0
Mmzm5D4w4xogVQJOzNB+vmZ2YPBHOZiqrZ5ZTz+nWptzwRJ0mB/WudjD6DGkjeoPrxtqNsSi1juu
jTceIPj80BWStIOwK6IebtKQLF0uaADuSVANb/sSrLmoBhUKi9bt5lpIS0dvm18X6aYhoF/ZUIJk
TNhKZCqmjpkuQW1fFZRh0b+w2gDcN7+IHEGBZM+b5llzZ4HeeCC9TRBvgOzikaOstOM91lzAkN+F
9bKLl/PbBeGAgkrhtInAKpgDdcUBAHnZuO5nzy6UMlQGVFTIgEk1FVrfuHe0HKDZPWUUMws1wIiT
n1sFNIUd38q8f/yXpUPuHWMO6h0tB/iMbBQKE5DXa6vGTkF8ecDRKi8ZserHHCti4swMzjgDYUfN
W8yXYZgrikCRIuEvbfy4gxZsguKBAaifU06DuvJSmxyBCO6byiyFeVa3s75v8EVRSJSj8kQdkxfG
/SD4NSWlSaUvmftrGZmRv4A5G/EkPkbvybV1Tzgp1yUG2+r5RDwyKFF2bPkUdVW0ld2SR5B2eIAA
Jslbpy4Jdji8rW0vOqNurca0/IpszontDPO0SVsGRMeqbg9Xg1SsplogTAnUFccR89iuaVEeKiCv
Qg38Y01FHC0TQs1cqQ4GCjhCgK6b+KRz/vHfKlVSchqwEMf85/TDcFtkdF9OMl7JSM1rrfhhKAMy
iR1CiRPMikRzPOBptMDzE5x26sArIGdQNxgwZ0WKZsQVzRurq74JveycDMV6CbhLkQHlGdW+TN8w
mIN8IHrlYHVTs7wmoQed4PF8em75Ma5YVlTIEdDdf9nsnHF300K2Xi1oOZyDhhr2IXY/cWqVyJ2b
USevkcMNSAXk9cW1scyYIlMQ0Xsuw+9NcNpymFY51CXxKB2gtsxNEAJLYvyoxMvU26TKwT720OII
1unfEM2/bWxWJqiOJ09SmwF7H+XxICU0GAN58iXQ5xxTAM3/V/B02AVDjCBG33/XzqP0SCYgUSN2
IYW88f+Beq3Yc2m2RuL+GaysPglCQgBV+p7/dV3chsNnQzOOfzQk0xppU5sA2eJo9Max4Zqjrd+B
eOENrpxvBv19bAW4hLs2R01FJgaM2mGndaKJLhmYh56jsSfzzKt+hi6T5lQLfkVNGD7wiRgmwTAK
jgiBIeW3AMIsyx7ImvTLz3JrmrT22lT0bdifW0Fgpv9AfO8Mu8wdj0UospcSWgJODcfwneL0OI4+
Cnip4MAdAJhMOML0+BtxDPPMawyf9jxtZGp/Fy3WyUy4n0kfp2n3LYTayQIO1K1qVWMKw8xDnkkL
j1t7g4ekBZW6Ra8aqa5A4o0+5llMOvWEJbMBVO7Go+3gkW6KqcjybApRTxMlmI5lpEUhlnlc1POp
rw1YOPJP/R6U/lVPWC3dhGWfommVJD+wUY/CNNiE0iQL9oV0hxq/cpR8yeO+A4j8Z39LugVI3SZA
e64v+DRk/e2+RVcNiNTbu1S0VxskLId+5QewhsVA1IUvXzCzJ5O0/9qrCSwpsVQTXaI5JOd2LhTE
fLObjzEzxKTVZ6ZR2/8X4k7rvSltG8A5nREsC5N3StxYQwgEYNDtH8zptlMtL/7gji8nQAOBhTkp
8/3dJDSpDL2/WWSRuRBzem5NA5YTzQYyWQBvPxYMcwY0bOz116lvwhg4dcQ6G9MxsW+Efj3Y4OXZ
mDAMnTrGQh70FFxQGXwiT/spOU2170K2ibhFKmHF705R/PU4LRnrzEnrUo6tDg0BbL+QIXvasMPA
iHFD/7rmD6bnUwN7tTkrk8GyI3QKq6We+85/SDj1kLgBoqRJcI0L1yy5m2cxU9uJMzq27/CoG4gC
X0sl+YwLAl8ivypqbRnhQhgOMQuoCoLT8BdPjg8VBvDL4wO2oplzVDO4i5rsVUlqouKeNbqsbGRy
VnWa7rny3gZp2wJaaL0b5CbSp2awz+MOqgfeO3Tgq0ZXp1TsiSWmTj53wt7p2D7ngf7qX7nk8tTx
d2LfvDYzRhAJdobZVusiO1b8qYzc9VjO/WjndLL9GTmKWBCLa9OKmAmvsgg+sRwIUijJ9rrFrloR
GqC2F39JGBhIFdxkA6lx+2FP8LrSIV7zBajfDGksW0fVcRO2XTkaHXGmBSKFu8yoLhyy6DrtyMOO
IeE4sM+J/yww1atyjCN9SWOuEj+VMMbLbRxy9+C6GvWMzh5QlniKdvgYEGKZ1H7TsIPFZM2EL5iJ
eG0A8Llj80MpYqrrL/iBN1RMz0VV3L9anBY9oOPRzL9l+tYInJ9wupXkBPDSWu/wQJlEelxQzQZJ
ugZd34ITUCVdECF9KWnTVQDR+UKBmh021t44HuWEfdBEISCQrqDJWzL2tyWZvL71UPveo/ghyyey
MtFJBCuXWt8sb0xjN+SnQIXv6dG2xs44WTDzV1pRvv1I3iHDZFyo9dN8Cc0MyefxUKL8An+F9AtJ
FxP8dISLjEgdIW7Vr5vUsUageQZBCZ2qOfBAJm9R3jaI0I+vSYbucdIn3GUafNmaP/y/lsyX2vpe
ZR6/tUt2ywiPevlHcSjGECj0A4TLirctEdOx3Jpnz4e6+TTJaYDSFm+FCfSGToFjTdkRbH8sd6Xo
IWA3ufn9Z8//A5FgrrqN0oHtZzvfFdXsnwk7qulhBgBXJIFXbJNreWTJ/ZA5bLu4BzLmGdR4k1TY
37/gYOkdg5HS6xDFD3VVDQspSTolukLojnANwDCs50ReoQXUGzDvUxtJzu0rVOtKVbdE/f5PrMIB
WDTncauhsDTJ8c2ulBEtjz78WEhXG4wAk+vKa75BdQBe5TM+lr7wl9eavCN3GtaztpHHrqrWUL81
1R4aStqxcIZthJSd3DxICk73iNHzE1iV4AvDVC4XcLnLTNiEaotZFEFl5MBpcuxYfe4fzrZ9HDRA
Zkm4afD7R2ZsBtPmIDGInn5Loa39QyhY1jV76WeCXrcZWhr4JyE+ag7dPW6YwW/AqPMkfAc1tLCU
i9EXypPreh1ODuA5bW1L3ZsKuNSrs3UosRt0Uof5UuvCqzxTWINaXbS5J52PMobQQsQEeta2OiSr
fZXdwulQGRw/Kvyu4eiE9tQ9bYGFTYC5u+WsKHKasVnq+XC4J2xYiCiPQb4U3Srg++Ouvs7yQHLk
p0cfWG/QEEz/uGMmGA2CcpNR/+l6zRDwh0knJhYsKJQkIxZR/E05OR02LfPKEITyE5bEUY1EW0jn
texWuIM5dsxbCXFBN+V3JZrVV42pliTAS8cD6cnXh3CwgL9/Bis8XU8mQkNSXUbinLTnAa//U0Ny
gPLJY/5SHIet+w3hhQIbGC4RFK9v9yTORMESs3tUlx6iBOOIO1TmonJWGopSFpyKe7nrGAbBI7UE
FYkUoQncu9fdZiJzefHG2UpWaDjG7jfOP2HnX4Dg+QrIKUMCGTgYrY4tN5gQtf0i0Jt0qTTk4pB5
RJAMaVY5MetY6GOKtACG4Zahg0XHRrUzUJU9rS+09o3revuQmhxBt1hoXqqowK/iU2XjPbMZRzv1
76RaUXRF/MhLQnN4++lAuA/lAbS+wbQ7x896AYH1nsBiejtcbU6HgwAhZ1WKbbtLeiSJsFmj4T35
xgydsHUDefXh1aEfjATdI0zG2gEQZId7ZV0oir/3Zw7i+nGRbUc/XsSx/Hf1z5aDyBtU1grjnGWw
KoYjyAaF9nX3ceR4DaWo/edesFD8W6fOksXj6shA0v1w0w0RaJo1aKMyW5PS6gvKCnXVm3oPOmiW
ZDkU9X/xXP4SHIw7iQ7AWJKmGqlcMBnC3iS8rKvmjGi/tjXmBcx/Z/1d8yeDcmxEU2aRiFwXIPq4
V3pQ+5W1UhZHTDj0hnsCzYpGE0M9YgQX4nLTvUdcSO74mI+hEPsIOAKVhZuhZt6R5uQnRZsSMLdp
I6f1wzrY3/2A6E9rrI/cK/mShPaK0DtF9IIxptVkrGTncm17EOp9UHPbZD/f2MzCEwFXqmpI+nbk
aAMYflirOuYaX2VTfxVqhQZk862iSv17MAuzvNclZ1VD2faedebF7abb8r6ROQNGEjX1xo7DSbJr
U70hveVcayJhBuAL4TjUbgZhciJ8PK/CD4KlwbbrewuqtLkdXP3gRgwQ3ZN2u+I2MRQIBeDqgBUt
tFduRx0GvX+JFaoLtEtqFU0kswj4adTPccwxjuC51tm5E138UMc3aTD/gBzBBXnn4DgOF5KbLlxu
Kakh+aDXb4L3JzMbBz1YImAdv2A75gCKptV9ZhzHIG/mPB8jlJdDZxB39Fk8+wWCUy3GrkgqQRBj
ti0g5ZlW0AqMC/1mPj0736gE0ZJ6aNWNEvtMXfF9sudkLU8pixJ80Lnz0tbAdci516A9Ori9m1Sq
tzJxao2xfW31JB391mUoaCcm5TL7eUaaj9/Iy/s6edT3jbCIzLhpOGiJohPmR6oZCqaeZNHzjkQS
w78EggAdHUF+kvEFmus0L+C7z4cFU16OWMrj61/lwSTCruDFLqxGnfuxXBMPML/pBb3KQvzc/L+0
QdhLqy0siUruQTzLMijADAsp+t5PfML3x+laxhnRNrqTisoDlT8Ec7wNIq0wQSZ+cK8wIzWCuqmT
//9JE32WEW+ojqYGCaI1hM7//AF3zjx28aBFUYoFYicEBuFMoxNEXDt6HssdGlSEBzemiDSxOj/8
VpSZ+dTZ6A36XerzuVMujr2npXFljoQuFYIgHX9/EiueA3k0nkTwNspicPgyKRyrBIj3TLLf/hpA
tjOyc8KaI+8dayBpBi5QPkvmcUn1yCYgKgIsm5tDPirSLh5xnABJ/nBXcxzU1wm0vM0BCQ9Oz1Ud
CMsY3Cr82c8nzbNJImkkdeAqp5BUWrG2UXfy9b9QoVDuxyzV/fr2heWzF8eH7Pwip7CsiOURqyEV
bPSCLWkqQZsoBCf/MLOMeGpboJSk2BQXqIYDogsjM14GxKnLzoHFqextJTrd3M2frqAHpfTLMVMD
03oXSwwdxx4MPoFUEYL3eAICSruonpXsnZLecuspKK6c+px5fUddy1ZturpxjlNvICYdjXXbNXzz
62lXAkj2rrUG3de+cfytSY/Ru/8RWbffaVavOPgWTngRbOJXTG19Zonmy/MzpY2cTBdbkyJHf6PC
uYBzA6byoedvk8OWTaHF1KqKJf08SA3Sr6yqbmQXanw/AtVZKt6qOJEkOeV9Yw5+AyPFyAlLD9jC
kuxag8qQU+IAMLZ3e3oF3eNoz/Q+IOfghwxMAMuVnBroVPHO/z/GxIwjXNH24rlrxjueROXA0mNj
Cp5ihT2HBeEtEIZiXiYoA1iCfLBWvHPxJie2qR+WxyPs2pw1DokBqK0cT3Y3FOytMO/uFtSDvL/z
opnS22x5qU1WjPyhwLg17cRWIcBfpxWlKZ95k7HjGd7/PpwsUmu24PVCa+RDN1JU+cwmxkliJNMc
LxvRooyVKvoIaZEbL2l7kyKIuFWzB7uE0jhswKTgE+z+6ttsJGiDIZxoSKYXc9n1QVJvphatGeSv
xk1dcK5AKacLPLp3zh6R/cu6E7MQvUfrwsX09WqB6kJigkU1g8YqQ0nqlY49P3fncvhBT211o0eI
KfrseXrRxbjhUZWuJ2OPqJFYeJNWR55Ld60Jpg+L89RYA4Hn+K4dtHm8LhtPMjVaVIr1PAr2NEWt
BRfVyY9EUIHYNAmv8xwn/paCx1AJuElxlKEmnvMialRp6vpbGlg5lDdGXaNxMgaEiqPQjF54dI9b
jdzC1DdbnM+JH5TEwM7LKzQHxUR7SddrH4s9vvTx5HvE+NVC/f8YWoV6Fb34Fu2Z0T3xrW9BJXBQ
3jqb6QdEWoW+5LQEiCFcXMx4tuBL6w8a9ABeRYh4zm1It0feVtjgExHPGAPmyPPhQBtKqYSDdZgU
AQ09pmxAW0u+n3Y4KrORoa3JZYHhkAinGtCY6VS7bcQo5/+LI0CoxGdvTESy4Xs/cxYDPEFgPq6b
ebol0PofC3n17L9BqeHMo4Fr7vBPtdGblgPMEVD/RqU4sgtoNTEhyWlmlL/9D6qsvkSv2M3uNuOx
kXNoOoLCjMoDU2aP+mSfYT5hd2kbiebZ2iJmw68B69EydL2j89FnE4rl1/Fqu2GfUCiNV9q6YBW1
2/Q49OF8cXr1K6MG9TsknCjFiRDCPPnpBHfhwik+mHaAoF3t5aC5GmwuHDjLfB8yizQljghWmxse
lqmm87VNd5QoIoOZwWowWCICNoC5htokKt04Mze4MT94MEz/S0xSacWtFQ8ZQNqh0yBdPPHubjXR
61F/TOCXTJ1WUWJOmxCeVIw015cJk5PD/XcUAGiCi7HlrMkloluSKt5LPCBmOOmJpjhE3EEul1/J
V21TOM9aTn27vlURVz0L4iDHoN4YPTVwA5OBEQv/f/hAzFREut/FpNJEraK3ky5167Uu9vlLErxW
eIkO0Xkz6slDPUWdGEmFCKn+dj0TmAZGa4vyzfpVRyIEcDQ8pwPbbxE5KITQ7wzyk/7OGwSfOxcv
NbwSr9+N7fTFJhuVSVWEE9E1emm1E0MmaPhkdoiSSn12QSjEfqZKU8hV/+6bfH7h3/NjR+/MlVz+
Ko74JMhlmEm2h8Mnlam8lFD9ee9Nhn9+NQnI4LmL1rHqxV+2dmOVRU1hrqyRroPjc53UYdRG82ID
alYlUTMYaw7u1uizLeDceWk3Ep1QI6694Y7ZHlFmiyvuRHFdqoesAKgi75NacRFlxS62S4jLmVBc
WzVySkby+POZWdue3Oz+hOe7LwX/+nEqSs4hfDPns/jogvI+btqJjmdd50mQ4dsn4USXWbmVsQJo
ZXaQNgO/SDbFumxykdkbZWbUt0N2QABObiAHN08j/DJsLxP4CBx9hrA0VS2HKXMVYYlCHy4XPtAi
xKunCR6nupEw5kEIkAFAylTUdw7vvtuvGS06cLXXbQW18x3jzN7QigGHqX75f3bNAbEIuH39FFQm
sXaPdB6e4TIovUbRLGeF0JWfvEm1NEGiCp09WJH/0ZJPcqVVn8radTnMm466x4gdeD9zeWFUFR0x
U8egvZ6ODFf0P+hJrWln3nk3urxkGT3/o7boY4XZdlBovDLsd8OMBg6AN1HCQcrGIqPsGNZpDd/L
brtY7Ox2yOB0P4WqtyfTMRZu+OHtD7oDKjXfmnXoMYVLy29H2Ve9DZaD5O1OM4nMLLP1LnwkWSzu
yCU0t3wuJGh7OGp1DcnakA695HdFltXefmxxCwzKNjX2I67veWsOMW2ZJL56y3MWnl+yE4fkMUSz
B0repLlTyer0SvVrIr7lnstAvkK/EyJBvO31sQD/+wdKCEytDNXvbjF1lcDzKcW7CaJMC939KSGW
9/wkKQMkczMt4WCMEULOBnJSw5xb1RrcWeMwV4Vgo/X6Y14/sUVe6suLpm70P/adTPnuf3HsChrS
qa2hKKwQMaadRw1xftKCObwt0kEWebgPwgyB2BCj5FvUjoJMFXYij7JVwF665gXn7oUIcDgNQun4
yfcxUKOghZfCo+5X1s7Y0vyAxJA7kqWq6qK8ZLpl0NQXlhGj1LMdFva1TLmkfYKgUX9WCVI28dqt
LJxS2wwsios77XcKrIy9q/SAgruJDxBw+IS7IKcLSp3ywb3+L2R/q/cVgCCUYyMp0mfxt+ce5fjg
XomLqHc39vZv4xir/zTnuk7mLlmoGw7/qxlMrqa1DzQ5k23apbnfcx0FeETBJAEtVOjTnRBXyDZ9
3cp6JHvQtLdI907VmmMHSWg6K5A590igX0mc9czy/iza61XZ4LMgfGc5bZ1NDzama0N2XTGGsE4U
P8F8bHOM0fBkCfpPhzcu8SZrSGgrQLaNUS7HINuCnHIcF/tR6jKPVNrTkPqUaSjc6+Ts+Nfnb63z
ylbCDfCc/J08l2KTtscNIekUDT+BGGtUsEwuxbY+dmRS9k19LuWZ8nfa44tss73ykR21O1NPByp+
yeOQlAnWZxVuPg5HSaUJJDNRLPpbl9DtR0axLd2FnpHTfS1SQI533YJam5RpynIfC+Iy2366D43i
qGKigdE32ayqRc2lsKfkuhRqPRVFY5ifiDfyb6SvRxtVKXO+xpBTbj6LH8nXJWTsPNYIzOoT+Hye
O4kTCfhLtOgvYcwHTpRufxtE5Prb3Ojsp5UbxDJKatW7zPVZ5BgMS/KqgHXGmwvmBo6xRKShHAAQ
CmT5An+5nxmm6RETCysrWhUehXHg5Wgam/IzDZCn6fXGjJQWUq2veAKXxJdU8/3R+taF4TZJHQBf
nG4rSgpxmukeYY+OK3C0Ufsx1zB5U02I/lqVgGEe7hMfVrZkB+xV2vS4rmMVq1i3wkPz1StezJcG
i3uoQq53vuOBYCLlWJZm+9JR/qyuGqITTBphjZHvwxbS4LMEdlBnqMBEFrWu6n5k2MWiaAH2Y9QS
dB4HnLKUeOSxwS8RUVuwTqJrCSYht3DF3R/aHTPEngGX/lWz5PxTf43PqFoa0HkX+D6dQeuR/94U
b66rnAEaoCV7eM4R+Lw6gvFdHMpUt2Ro5uv485xppUFsguwY2Ty+J4uDBd4Zh9aU5MJoWomiEiEu
LUM98cVkruyQrh91afdG6DVRQ8xAZ6qs3f+eghKx8TGQ68dHv869c88QEjNBD9KH7WGSoFJT0qqL
+rkdNcUq+pj8ozsMBBqUhrShQTsmNNBgk4lerwRK8VFBSXAyGyDXRhYmJXQdAtVF5lt34N5kMxMl
rr4AzIjWchRnBgVFOjsP46JTWvEDKLwKEyXryl9Ny8OgLUecOyod439TsL5CmfrSdigVsuEifLe+
xOocF6EIFP+6JPH8xmz+YWgITCfnQ9HWN0tNdN61HHlvQQugTKSZvRIFcbvLtOlYk5kIpKfrzjCE
w0FDnhADmE5/vV+8hnGj4B0Ri5MgGN8az1JjdTD+7lp8oyqCWwAsS4gBz0ea1NLU2XUeWgvvPbIx
+B+NUWeTxP4JDxBKQOm6FfiJuLICUlCeGSZidJ+LuGKvcPcKNTimrcvvAUgiMGUiZCpI7dENePQP
pfA/z6YOcTAgVrK4md5gOfdUM70rvVyGPXW+JUEZQrHuHCh2steI2sF4gPS69kULykx7h259LhWl
rmFalmq/Z3Cb+nCVrpzUeBJyFnPxepjasExQin5YOnCKG6Hom89FymSbbJrQ95prVLMi/zi9J5z/
pDeZwF8eEAiHmfuU3GKB8UI8DWS+KArPGkY/RT8H1b7N848/Sxj3VeBqWWpKYvBzh8ydHKIS64ZX
TlpStFTIDtD5iPmu8gU7fUXXFB+lKng4oG2On3QmpO6ZFZju/LF8b+OdBhH1KVnmlGkQkGzXJldo
CxxRzYEG0pGg4YtEiF7rAfUqsVsw8jAYtDNxI6eoo7AC6fqRQXrFlVIARcps4rUBK8w60v7X2XfF
S9uvMfVyoNj7tVO+INba8J8yE87/p/vgBxwKgNgBIIfsY5l7dsGnZzMB1zgG79tKdFJ2EdsuNa5j
ko0HKvKPpyKgxrINg7y34sMdpFWcYOqpOaBkM0stJhW5HljFcnboZmsRLam8oWTV8LLVXS+hrDag
yalKSWHqEjjKRTdqnB2UP+polw3hKoKE9yOZdthPfijU8acOU/ft668nf4vTllsRW37GaiD3r4x8
EYI3Qq5ZAfKuuf4UvKb/ZXaJT3otzpNsg9VUcgxj7rZzaQN9vmqSotrgFWlJQy96SXYxSw8yXjVp
Smu30TFw+H7W9Uy7qayXvRAmziEbm+xtZdpnvuwUz9uyqxdZcp/6YJuN5g8C99foCX3XvfD7ZnzK
ZQdQrxlPv4My2jI5gao2xHwm+8s3xDqm311Nxyx5tb+iD18vVKGvSAHuyHbKpXFempyRO9ytxdPO
X2WAahJChMACyJGQA6Z1N5rxAaD4o0wLTxo8AchKQ74A/vtUgJtfaSPaQVaY15GpljzP7o56LmnK
5iVuo0iMyhjVoHvGGEoFpytlZLM8PcDZlDnsQ53kCE1+sW+/1h+lisxU46xmhVf44MTuk0tlpSgU
YX+3895jykQLB23J73Mp+fk/zlqqZbqy7xtB1zjwJ+ztGaWS1M1LNCbTVGZDZvTDJJT7RKPfBeMJ
HKktHwib8NkMJyJgsTAYMQXOeYDUvcLk0FlvjNpLUY+P7ItI2mkEjlN62wX//cQaCuNYbYmwnviK
oaH9YyeapGGl2rWuq6b50Qq5FMSKRChartGBhy5pNHI/+S//ZpG4HWj2v1nSh+911fH1UrGRkF/n
IJbrTu5LNNttRGlynkVkM4RiJG1Gnd0OJ0fccYUw6/rf2w8Bf5xN0wRy1yOtBS/+1/UO0xa4On2U
um2Is5nvGjKLltUth3uRtu33Q77Oxzj3/ATYxMwL/BX88eDCoXfZ2nvOCq5BzJGwT5JwXWK9mCU3
2rMsuh5WnbTlSIr9xAIQS5HlW0i4XpqwYkPqv4qjui8SK3iliFpB5bPqhXivKeZiTpZXwKtGNp2D
A7OTR/ElUwhky9QQ7pQpytNcfLr0Sftr2P1OMxwl25WKyaBrlnIsI41rbPKhx2thGM1YJ8qCl7gZ
LbCWng3JB+QCTJtPl+Vsm+SiaDeot6Hxmc2xyb3lkZ8U4eWrOB5grnn8kVrsdI+FPcJkw9P4v1PX
uCQTMqbbGl+aJUFP3GmVsR69SVHtFsXvdurbVF5SKZnfdY7I8011mW+UP4llp0OQQDlY6bziVQNO
JZUMKCdCmW3QX7e6ms2lZ8Q79bYg9YDRJB46bjP3h8h6Cg3Fs9Bv+SqpcVf5dkTklYCFn0EK4xCs
mbunJoBfkD0ejsm1A6n6TnQKWard8zwJbOTlotzJd283FOIT7BTwjitgCbZ2BioWIIivBf8sqTyi
XMiu+r1KCGtYNSofMNdXZVTWDLWgK9RPpZl03QQoY01pqBePhS0grfp9RnJ3Fk0FBDrtkTeHR+U9
1PtwqGbrIq6dOiyKis2eFUgJoGo1tbC20s0PAPx7aMbXWETXLfsr3SVgn/ZnXnvc4u5osTrrD0nI
vNxTTk17F9rYtdFokWKSRw36D7LEcLOuqbrubGFrEGa5UJY2kDNXGUWFePvH8DrIl2qaodYyo3Km
Nw0DyvNuxZESYz43HPevN9Ex94yLccskUxvDTgJg/UNGu2mjgJZ5VtllSFdIFfIQLAXtPXZ5IRLw
VYMR0gVi1R1utOQEt3xg40CRy0R0i824uazudFLcajvae5ZplYmfnPy/pvDlg3vnO8SVFmFL+j25
on3+R6EkSZ9wiVSvIBTyaZOwiw+clS02WjVSt/fHs3IawbZ2sxb5Tjw/KMDC1Im/RSTVHYc1h/eP
6vz2LpU0Ba+EXurWKw/WoLi/04ZjmrNoh9UZEUvEShUVarIjwq+ii/2HqnZSKnVGAXYEM+ZpdcdJ
HJ1tzScPEwAm7zYuXyeEsg/R0rnD0vkDc8/TUI1Y0CpEZjnvJDcSslXisEOUTEu7PIKiWOZxml+J
g7r8WRMw55nWrAc+/PosZTHguiOZQCW82r8HPAW2GRdWGg7Cl2BLd5XEwY5+HkhUQAokk3DtSHcf
1aw8Lo9pFP6jNI/rz2pcQFernhERGijFR61eaLj29ALHZV+m7znndsKnR8UEajotnWJy7sEjpB0P
ab3oW2rmWmh7CXSutyj6py+WmQ7/uKws7Vjs0PMtCq6gJmBkT1NAD7QOsxTawk7WJCXnplv5AynP
hQzEqwgR9swyGR+/4mssbgM+kOzTnGp2tPpA1AkLduw6VwU/Lu9c4bQrppnufJQau/NfzEqJimTT
U6E7mGk9NNRmrk56PorsDaYO3QQPIw629x7Wu5QLRHwvJ7qqL+wJABFpYyOdIUj8F1hiUxbODojz
sLnT2N9MROwcfY3cVwjuo7GexohL76aB4Sia62EZfaONC4FPzbRdQHjm6ZaNhyQnQ3oXI6em4Xsc
mhNTgGZBHemvFheOKWgeLJmEzifRM69V5gQQUwXqu7RzHF3e+nLCz+x+aIrYDlVYYmVkc1mdJPeB
3+Rlk2zHhwnedMr/z6I1x5HtucFrDGhE0YEY1MkwxPEEy/a1mu65tP15lu8taZTqMkMqisvtHuKK
G+Vnpu6dhLev9dCLLft9xGZIyix6Zzo1msFvZTc80Zfw7fZAl1nwXon+ft8f3qwXLlMW+0c6wwK9
RjbnQ6WEtJIxjJCTMYWi8MyiXHPT4mkpVLdoYIgY+N65I055X5yXJrQ9ejO0FdXWtxcPdzGsWS8+
IWSNXPcVzNHggc/XRfPje+QXnq32ZHD2PKK1UKyvX2TtOfGlyp8w0igYILX+pFlrwkcQwdCjXRVa
u3n6Ddxv9RmAlEltgfyBDVhNEKm1W5CWnDkL3J2D7hLM0Xh7QrhKuLR/0+tMRhFl0gNL1ia5cBpF
S1OeSt5Klb+NLa8fBTzxhzJdBs6vARfaJmTlXMWPVEJqtNGPWCm4o0gxJbysiNhfT2ux+I65G3fX
NrDRL5zdbP7lHtg0ENk93dFhp0oHRA7R8KlnYwqdNRV2oUUeOto1VMUQgui3coligMGjuoEMcqVs
Wt5yOOXPoFrI5aXbwS7mZP3Nl5mqE9rH4l3NqKNahedb09iQif6oRGHMSH0Io5YBmLYffisEZecz
+kU0BAnsh8pocsx37+qRaJZrqRWvHcggJb2ln4G8oU+hOyuxxCcN19xsWG29gpnoSvofBmjotJSs
C4rJ5aIBFOtRGdqHJ82G30KBODuX102je/1GKm2VH9Y3de3Diy1KE/nTTJxOQT2062LbyeVRBd58
q0bDCEYjdSg4jokcGwxzcEBrkXKGY0aYjV/l6MaMYABEhG+noTHWPZ9odoGH46fEH0loKmXHNDLG
LTVBOZVz7pY9nt8BrTV11sbogvDSUzjkIOoOZNfK9lKxkUsdabN7ChS4/vpCZLxNRihqx+vR2b5S
SXL0oRPgmXKOYGv2KuLRmTeQh4gQpnzBB3G3mUMXBbXl2QIPhOCh01ZK0ZMAlSumP1EIMmXVVy2p
ZRLnJAPBGcB7IBF1n3RDv+pvnB1p43Jy2OYu6lY1F/l02zBpDC2BauaWTTkaC0mEwlB8nnONuJNs
ez5032VbORxP/uJTShES7XycJ57+MN5Y6Hlde6hC/Ivzg757wiE+VAD0SN4N9wb3HwYw+hw+6PIU
y9srw3HmWxoh8ps/jwBfUJQJsZNStfTbQtkccpisAi5bac3I6WztZAH5wlHDTaXjygYJeRNvtGyW
c87topb/h+CYxiWIDTYQjk2/W30h8jaJK35y0qRowMFqOuYKoL4EiQahWTEnJxhfAWNf5Mn65GRX
BMuIop3+Hrok2I1xyS67PamTKnC7x6UY/6v1lS2wWr7CJ0sUMcszzau7yPt0+nHJ3wrrJJqQ/W7f
wWDXUEc5ay8iROUmidErRMMKflH1Owmc3PsYW0hBd2e9LQX+9//xUi0TKFnNrEaXEDaINnSBGKik
qH3SoIICBKO1AhMj6fhjmMU/t8qRuYSG3quXt4ucPIHx/izDrB/tPYFL3npA4VkrM0zN74KQRu6o
ONXpbriQNCdQWjma1lHCNsZIpN3Ecez7ElCre/9kY0NYQ0oLG6x4s2luqpZDk31usKtVoWMJ5vUF
0G5fD2BS32qP0JFtQdmeeZNxQyDSjgJcmvSNL8Oo47UMmwACo2if9RsHhuKEvcZ9PSpp+gTbc+tI
xKgP181cvFfWAulqNdTp1K9TdJLEBAR2YqujVxTy7FbAqOQzRUhlsUCjZqGfM15XHjX1/i13fPhu
Xyzv/Da8k9VGQiOD4Ag8JpRYEo1Hix2rFzCFnCfBiwQzZzQDo15i2HiYGQgstpsXQDmzigrxej2K
jWWpis56HGjktFjGs+0pf/VumiE9Hu/eFrNlIKdWXgC6IXSu4lmS4CN0qyxhJW3bgnHAA4Gd4bzU
vn4Y/UuvTQFGd0HojmIA9WWAuCyK9Cd/n7fNFQP7kJMSGeaTiC/mcNHztz6PXgje9HZ6gRCW5jO4
SvR2DJro3e3A9d1Pj+0DUFR8M2/YbssZRePE1WhPsU6p4FyC2kYaLcie6Ty3WSi1aqqDbfQyJfyp
5f/nMSRQwJS16DR6gS9KjfxHRBI5C7YbJ5FZjDv+VPuJ2GG4NTnqvhYIjsuVdiwwdPzn9NnjlUIe
Di9QGKPmwTeizOaeODx5KMFJDsfqVDkO2fmh7xc2k6s19mUoiNiTw/PfnMLeTX7VjjmJbKGY1qPV
3BC9XE97L6GrU3T8/8Kq734uvPvW/IemWwd5dWYdZx98NzWDCqaKpU+z1DE9TZNAtVxOkcDkfpdC
G7xTiZ8Bn8q+rG++RT9uFxkYfSlrAR/EGuVPr8kYfOvOCiU/NmopeNJv9JyJxCyFPLJlYVddYO/5
T616wYyEo7YqRsYayv1b4gBb6/VoNvPJ2wBAk0Jh/920LKWsp1sqYKR+9HXPNgdulhIhFF0J7WnQ
B8ZNS5Y0l6Y9vR1u2CobcEHhTwBcHmo3eYpgyFnntg0sUIWVEQSiARLgxhwQ6rh62V9TwhN5EQsB
aaYO4g9yS8TAsi3kHdJ6+ZN4/yPBN4xEZVPgJaeO8OEG3+B/KQvENW+u+0+SQdQEw5VaGfcM+gcX
H7UzDMgccSflwBCZgbyR/kPCJpNaVuH5a4RIa8k/sh86Gdpp15ash6nqF0CqgXNlR1CIMv8ann/k
a+1gq6yf/9FHQ8/jzzrH8LRRHv0JfbmVFHpgH2JSRltBL2TNy30p4BNuadblP870XtsyfWonU0Zw
j81U71k2U6JuQFyhZiYUJ0l8NlaFdjhVmbTg9Xdy6WW2t672OvBCNrMfliroY1SeDhA1rYxM6E4b
n3wkqdyxhapJKaWQOFHD3ouELqW1tHJixcCDy2Mhr7IbIFtvoGrYd74/p3uv/SCD2A2TY0dkCtTV
OKu4chk/BqLGHJTYMTbYxpyrboiVBOkIdYVlHEsKWHT5pyR0csso6vo2rWTlJvQQmqFZuScy7qot
78y6KyCeb0YiSCksbdVWyjB0Syf4FCXzlDvLXRpCLrG0VFIyV1y3UBtv9TsNShVv5wK/mzdD8SpW
jsnVPMARSnKEa4Vam2xbFdmwX7IP8lhnWda6KhS21z+POjvPTSj0+ceW498m14aaLMqPhfTgZ0vO
mVgPZXqB+Bu+0OGb7tvqCkhmCobt6evkygr1volTUh55gpOuLfWhBxNh0qHXCgMMEF/kHoIKIvCR
6R1wt6mSivoblwMO3ZAB6YGfCTeTrm5Eq2tNor8bCYHBJ3xjVW5aA4kokxB1ojzqm7wQxn+VWZmz
U4BynlGozEKTodyNdqn2cz5xcjlavi16WtQfwM3cBOXzopJwRKIQuQ4x57lH4ZcXKc00/aHgQPEd
YyPw7hnaLU/MCvA6h3Ph0FeCmcB7UjyWjgQjeqcfPnN8jEibmiSMd2D2rEyaF0Uuf3Pt05iPYrvs
rY8VnqrGRomXNDZE+MLjqOzDXojZJfrHURD9w7DceP85UCnJJOIOkvze9fqmRz6XBkW8Nrix9LdK
htxe8AeY7hZ+oYtwqLm/3iunG0Hxb4tya7ktAFNGMZtCZUG1UhdOzoGvVWBblFz48a733h6osG9a
OpcfyRzENIXt8O8ZYf1AFizFGX/JVNs3NCJk0OB2sAiclX1wjAdnwfZ0DP4riS2XUeGoDimibhLQ
oh5JzVmSPcK50adZxiFjPeZT6PvVBkj589t7XRBGUfyo/lrTLeWoLhSi2mzwI+Ykntc71qUmLdVr
aweYW4xMk0zj166Bw4aF41oOaeFQosjvDU0EWFQ9z+tdEI+AG02SjntcFbuxRt6GFjugac3bahkQ
rMSnWQOaJECFf6+T0PCv9RqbhEZ/n+9SoCJ8niACq/HEQ2JKbLooMmWAuU3iqFBb2YPNKV4L+Qcb
bboRSrzX6PuLsaY14CUq2mzXuH1r6EhtUVJeIye8ZEeuqi46cWXljvnVNn74n7gFV0tiJstj/vbV
QwnOjJM/n70RG4S134JHO+xSuHbR4Te4+TQ0P3hPLhkj+V0qb3CEku1PcBLfktdrmDUQFsfl3QXm
NUrPJdjhEvdL9/NplZ14HVCUDGvhhLSVB/yRAiCYNX9apoaU/qDDsUxI1eudn5T6RtCyG6g8K8jZ
eoGfgChe6+l/XFIcZ609eL/JL+N3tQF/Id2oDAHEJiACgWAqbM1cdkCC01xcq5oX/yUnF4KEjgaE
maS0L3bJ7QNztV147AvEGNUktWtjrzS3KiH6shTI59lgl37/CYbB79Ikdw55acpfM0jT3QGpmma5
B0lSNCVA8vASWwQXQR6Z24H9M/AaTpo/kngo8xM/dJ4GIxop97MRia42gRFeAxyPRYDwE4navOV3
CoI4ugGlIb4bKGayWTdHWrbmTRQ7C2Nwmz0f+eDrkQOaTTYtz9SU10TdU70P0NwMZBlnkasPOg5o
x7NDJxxqtT+F3jhNufD6hcPiDGisuDCbBd8rYIGyZV0w5KaT+8DHPb4ko5/RRATB1BssFzeIxGYX
YV+d1+LeQKyazCEaqVURZU1Z54oRFDli1wN9lZGFe6/m85QQzPbjBiEoWY+hLkYfEvygZIlgXwwg
0uUbR+w0k0A1yy+vi5DlwJGlimjkP7GxKXiO5vCXBXOd0+GAPBxLAjS7QKYEqItydPQq6CmLQKFp
6HRRphBt4KQrxyMJJi2yMuQPUQiE0Egx4C50QIn6HHTj5s9QBjj4YItnduK1xtEQf8L5Da8GyM4A
iZ9kdiDHdjf1aq5kaOBWTMidmAQnIF0aXPhawzHKHlX0fwuErlfa4pvbvhVmEMwvhjrNsBmYAFOC
MNl2i++Szpl8QPzbJABCUHAlSborHp0elGEfe0ErFxmRHE/f+UpU0viTZHPLMJow6+HOdYcMD0R4
d2GA+CnBAh38dIOLXDKpKpXNPj5qQRjB9E09m8HD91L3RriP6tG2MYds6SlEg4kr5L/2QLeVQONE
Igwkydcu7f2MMTHWJUhMUbrA+H2VErmMeNtufN0RUjHLTVmJpk2SLaLXvh8fkT8/BU5TniHm/zeM
t8hfWi6RH42lTxfqID6V5idb5ILZcoqbiA8kFPCEG2P0bs9g2VqCX9JwgzZWKJNvCMlfodkVaiu1
Kdt/9thvoCgPvGBVQwsB4OLkODuuwcKDvd13ikOPNAaW/vALiZeEJYHrc4KAaGXXmtlIK+YLWlHl
laa6PkUHPS8vOe0pwcckVQd+SrGqKSn758n4zg9RPw3oSO6Hw5qOoPxa+OqH4wsGX86wt/hAyNm4
fMsWex0SMx79CVzLdcown4+ExshaDmZqhD8FKL0poxLnTNrhBh2wPlN/h2Rlr5BgWEvpHik1UZFr
cSbsPUCr5NZ9tFxcbl1afVch9U941+kyixYT8yNgrUM/n6Sm3uurHZk8/9MriEijQrXuKM6ZiYr+
i9jlzvOlSa3o0ibp+1VJ35/cIx6KcC824dPyjTi5RZxe7VuzOAvJrDVVF8ef7ndR0LV3t6k34qF0
yh0h+kusYuGKVYhgJwUyRvnP8DJPWNnxDxOfV9YFy+/NCC5sHo6XyYL/4/rwMlnL+h1Ukb2bvA4y
6j7zq3xfunvg3a8fharGls4mbQAT8BkOMRlJkTEgxT7766Fj3s4qb2mNidnshMyRo043mlp7DDNi
3TBr+QQJIaNmn9vVlOtS6Mf8oYWU/ekSC7Gf6ZkXAv1cvb8S9fw6wqSfAXadi0KYIeRr+iacfbDu
4yeJ11HGPwRgZP1UjsVyi7cDYFZXSO1wSAMBecFiUohM/XJ8ADMeXze69f54XNaSB7i1WtASdR3W
/h2NzFYbHy6aVtBX44/ewIJ1Da7iM/rDJ0Te7fZdqYuX+fSYElQCJdBJ+sBghKbsnp84qizOFM3L
ZTXRhTyjeCQ3ZlNisD9oAAtmGiE+A6+V+HVxFcXGkVQIDBPg/ysbmb6QOk+0x0OZa1Cq/kuqLoFg
4KsPUGdb+kKzV+m1gafCa3AmmCW4/ROr2YjtFoFSPcfYJEXA40l78rXkMUi+ZP4iV8vZFHppc4PE
mARD9FgPUOaeOYAhrcYxK2EZzDLMkiCvVLAStK3cEohSGWEV0x0mokqt9LctfAwqvPXHIyVkeA1/
C8cBnucUg+wi58qU79eACL/xmt6NOx4ItmJKwASRarihQDjQm63QZF2XgNYEzfhEqjsQY65iTmRJ
z9mhMLfdwqiIPjDx7jnZ4oy5iwQnKHv8Z338XnMCcNeIq2dDEnIchqCp269R5kJAX4no4NjDXw88
L0NtuVpJNlNDKK1agnM/BB+ge45qcEaC/1XlfcaKvMvIxV4z3fdMm9F+6vTwlrqKbq3CWjmg/Bwc
gFIL3lsZdg3E+tJCRmL+uOPMIQwCBre7gdyo55oE7m+HGb9LsUyxtpW0e+dwH82g42QnK8YjJIqH
M+MJgItZmN7QUfXai9L6duJBFC+Twd1vGNdiD4Er2x4gmE6iI4oU2aljOu9l3yNY2/7QVcXUjioe
0QaPDaB3g9wrTA8toAbgVgwZGV+QEAUCYBXaKRIZiHSEbbCedU7sxgn+o4Is2JtWU8pYBEk+yKRo
af6TPnHqlWy2/091NzgoDCqj48MkqpUjLM9JCOvI9iGqH9tFXUxd2gJlYBWHIm/TWLUQPv8jC+QX
0akmDZRmbg9F+RH+TD70sIAun6wLzx2yIuQToChTAFg5SZEmWrBP59KZoZn7thpcaAWTzcgDQ8w7
vThpw0K3H2Z1auyEygE5718n+kJP4/2MZtQYwkMHRFRX4F9RWSidnro7rKB7ysD5Bm5wXzfjvXcv
VTiSrUfJxCFcsm02fF5DHeJE8kymVxADtjBPUqVvmE1Ro45DAUaKt8iYbNILNJFNcyKz54C2TnTn
XkyXCf07KRiieG4+8rgDgXWOTFKNDahfZiJP0gRJJ2/Zij8ZtgHnb0JpFa/roTfHvpLcrkW4+vx0
DEOFY0FPl/ctCZ/3269UFrNrRO71+sRouM3NE2e5HSiwhYeQn7/ZpsVGIHvxC4d3RuWFSS+oQg+6
0CPXkJ1zX4chsmzlr7C/gJWbg638cqFBhjam+RSMkYw+kAKJLyOaEWLyzwqyokhoniJ2yIFiGCXL
TJt7g11MA6xonkP/o9q5ngCibG15Eog8rJfXsPUK12Oz8e7lSwVW/clxS/t9eqMlyaSuYiUXY9Fi
VW/B486yi3qg56qTTZsW1JNpDu92v+PHqPf/tlWXOQbwA/YOM/acWtxIULnKAzV5sceZi/hc+FwQ
CTWeB/y5PQDw/TqVl7KRVdqFuIcR5/Gv3hPELGsNjY6i7njccftYTlJIpo9fhc9Xt75kbzykZbIb
FbhGNr9QnMCS7kiBy3KZWxNCSmlOmcUECH05SmW+nGf/G1vC9eyXNFh9pNSvEuy792hDufTpXYzp
dDoxsj2OKe5FjvbA0lFRrfS4reyxn1LD4/sj5XMcRWNbhN2RAhuFfQvNCjtcbLpDwm3olfVM1Kkd
woBP5Tt4iiGiwV+ukg+SyFvvUSfpXeLGB4biD2qErsO44hTjDxpDT0+wlbrtLxY3KubDquh7W2nV
u+P7EBs6bhhBz7VC7p/bM4vhP+SAeN+anOf+b/xw2nyMqc8iNLUJg8Y0ORKSBiQhpH3qQzC7CC4r
Wx3ZYrTMZLHiz9rjt7T6XJu6uBOLUfMxV5wtVmkn9ARIC7bMp40ABqcwWuaP37ILmLWmyzU/vMmM
rGtVdPyjppPKD8eO1+DMR0rH3d3Y8wpeWZJpV0X67afNdmeXQLaqpjHCJmjwl4dTS4FemlaJ77Qk
M+Nlzy33renr7R+8jFgA+R2Bwz5K2EEjBQCO4i2QGlEx/6eksfugUrP20ngxFzXLSPLL/5FiUebl
IeZMCx7UKl1iucFveOnUnc/yzpz0S26jv13pkERouUZ/M75F52fD3LWse4Dk12I25BqFQGLUMI5P
7bROELWFd+WWFwidU24+jcyXyFjtRIW/h8KM5g/FBI8rGFlvAm3WGo6BrtXPNcGj5lLLmbUt1gy5
9gv0rrwkFLCpWKgLsUkf5khdaROAkB2tx0war4avmFO1G2S20CPEMQWvTgEUYwMsAPhut7md/b83
wPh0MA36xa2zT6Fm2vo3glBAjTO+rMFgDiRjAfOiFjDZdOwGIifsjwlsbqkuImaSfoHcENKlMjpp
AToDNTsyG4MsJz5GTz0sU0F76q+rQKu8T5d+7TzwUJWzaqBh8oY6LCjzaBehapi/UBKUD78ra9nq
sveUXTjleiuoQbEI1fh8MpyKkk0/X7iLYHfT6BJzxX+pLJJcQkAUbG8pEML/waRDrQq1tLow2Iv3
C1k1N6eHgNgTqRPYd3pdM7zxgDWs9NHx6RGHARZAQb9A0TlCP1vckEsjgSXqksAf3ca3R48hzvAY
93rywJThqprj+LEV2TavBGj2own9xRsNTgvsgUQPiQTIBgLuWLcNtNhHawfVcUMp6oQKZbHpWwzL
t0+BETTtG2i1iyGcslpUXM6TCujD9/XETBmQpbgq7tqrYZIPJHXgGE99Z5DMoqJHjBlRbsgGXQ20
BUSVcXVg5OJruE+Oa1Hgmp6jnZwv38dAk2uSoUj0Ehq1xLANz3IILeuKba3T/MExrTKQ80BrEXV1
qwzWdUDgC5RNFPXhTXM2Q477m6QnhprPbTrN8WCr/k0ovFdr6BwVVMaQXty4BtWcKi6WtVO9+qMY
2j9ys9bdGrLggw8Vw9tSmPHdPBqFYc8rtsdGMzGGwZFR77eZmnQ8eRzB+ytbbo2qbTgMqPYfsQsp
qpozIwNJEWun7g/6B8/R3lY1kCc7PzcpBme57Ei6gIYOcAq0GTlojZKRkpSmKKXFBDcELi2c8xGp
PzcWJ76+8H2qgvhtwIbir5+DdxCJSQAIVc4sDzSTKQ2K/S6+93wp+BUAKdNechOll3lTN+cWK4bn
/7v6UKowg6Dbjchzr6PH8eoqL7XOFhI/suG/pdwgnW65AwvIN8vXv7kJKV4zx3jXjXMGk9gz+Jh1
EXY4Hppaax7EayIcfo7pI3a71Oe3wjcY5syW63JsGbneGGBtbigrqyIGJFHj/zFFe5v7U2Vw5qee
eVcs709/4QsQ/O0Yl50j7+UK7O9XDNmVrk3gqYZYVdC308gIkphyatTBXDISJ5OXhWCD5ePYSNC2
ik9wM7EKKzXAzthfK5FQoc27Qp/2DWBP+kGu5rOacSRPApQrjtK6U+xMzm0+yxbSsP1FhQKvm/Yo
EiLrs7hxZS+gOD/7AQY9O0y5zKQYH5qAyJMrJdfb7+VQSntEIAWT9LCGSneYJBUU+qBJq1CwfCvh
GLvkFzj7PbWgcngS/vSJljJ93mCtyruELDGNdthmJ1bkvjLVEadRI/hgsq3mhxa9aX1cQSS/a+Sy
EGOLOHBNLc55dpQJmJPoj3++ifcYees02kwq4MsreXqzozVhqCk7+SeP9MU3t8UfjovQK3S61KQv
fvcIvvQmq/1VjEO9h8LOWxcT6dSsI1KlQY3tL0EWF9X5Qvva0Cdyku9jpSiDeGzONFiKti6Zh2k8
yY67P88zK5xJ/7pkFvRMBl2aoaC7V7Jsxqac9VGypcVL4fSUZS1cvIB5MciWZTda+tuIOxcj/4vh
7xzB4Z1RAIQ+2tgAEFvCYk1+G1SBo7Mt84OtCsMqOjo3/zgYr3fZNqRgZ05xgJg2zEPMDq0hJSl4
et7m/H8Pz/IZqWUusSQYuZX0pMtpVVzZ0z+cGPfxPonwUxURhRYGl5vdY0qdKkxYFVdDhWXNGgJ0
xeP7zX+243zWw5BXmXGLhakiZe0Y5WlRO7FAVgYn8bqc5vxSACVDtySVpx9MKhEkvWAtnJnGfta7
nZhbZw5NSZRNT0N9NiFzWFM4nPg0gOlTFBOZuCsAsTDXSw7VWTOg+juG8vGSFKdvQBKWu0syt1aH
FINKS0tyem/LWmGIc5y5jXg/HnGAuAanVxkSHHi18VUq/fJNnZabTvNq5r+A032Dou3ZvJvjIApc
qwcpMTAhJKIdNEJir7pzfkMRJIUlGSRe1ASPn9ReoWUVR0iUqBmeZ8RXWaxX+Hx3z8ja4cX7eqau
Z4RmI4mvhZzf583OGIoT0cEK31CtGwr3bfnGV6IqPdUw788marZ9TH1dpRWfIXcyA0EbQcK87+zy
8i+48q0LDeKggdcYc1VMO4Gaz7Z2bJ/cuMuc7zf6OW3sKB11L4McEGcTIr4Zn5HF3eVyAWCJ3eMo
U5sIWLpCoAfgz7A+1CDYkJRxqVkg/uKea+20KEr1g5XlDMwe9l31gCy4qDT2LINHl48HnF54cgIM
4AxLAC++g4Oetr7Be+gCyx61ftGT/lWh1qgYPzuGbmbtNGsWG89o8wRQuM65+U/+8N362saNecg4
Q964BhJqEoRQ3/D3HJ+TzbWmaXNKaIrMv5WxdAlqm0/Qv4tNEvMn5mAxh/wgrL19VbcqNIP88h75
5LNghjvh6IqYVp2IrQgoMEMX+DXjTOAPFo8Z6l+L67Ds8tUFRlAv0SKWCwvCgz4oySAMsgE/lE05
9+9OVg3aJ3fSnsIoSmmq9flPLja5EpuGp/RgdU3kvmdI9zk2UMrU/XsXPRQ9ehF5YWnhUpIxsiB1
rN0G6tNfIMESzc7BvRKyXaIsDCmAdzdJsbkUQ5yl9+sGPIwcL2b7fBpytUY0+Pe3AYPtdtBjm2Ne
pC0Mz1BXHKS39dhTuW1FqjCiljllgWkOMXCE5b6oWQ9zmM+CprKFTlonTGzoZM034R8C5mEq3DhH
qh14KukdkNa9wPGRbyxq13WJ2LivV+jsaZbE7/4R4zj1w/5cl0KD/wVdFy7qi6iRz1OLA2N+oU/3
1UoE9WugtoyXuC7SoEghd/zqM0uUmMGxtimeonER63v/qRxY+ORE71T48DcqmdNt+KNzANeAHJou
dLQxc5m9hUjQDELewwk3OTnDFZ/z3a1BMoWE/E/4mPYLr2W4w4jAd1O5WxKPB3s+VjZhLpQCV2eN
oLIuWmSmD9VDNzK+9GBljNrEQXE544iRNqxNpuZ/eyw/vWUzleCgwqfGMyICdtw5LS4+IaxJcb5b
ZgYPn2JsgMDIOEOHMd1TIH/+mXkZb4GSYi5n2RwZSwa8SjoQUwzn/2JJ5yp8vYkWQQ9do82A+MUv
MwxVoVQx1Vbgl+YFyLJL8u5JdUbBUGnkoOBm1YPRKMspZ/iut6njYCsBErzrxJk1ifcRci7I+mqN
cwUMkL4nrsAp+gMYnrYOFMbJ/hrpZQl6OMJXrwvvvLKg3VEWAfiQLrd2XSBAWYNno4IfsPym8iTn
w8EWH2D7j16HTz7gvzxLl8wlkVNLU5ag5vUNNFpbB5kFL+d7gYG/nXa5X7PWjIdu/z6KzWWVO0hB
AtKdKPxqNLzUpnP520aUsk0VCQ1LsEIrfOKT1knn5jWa0Bpodp1+wHMNZ1QdONXRQhwoLovdxu/i
Rq058bgyIRAxd94bhG0OjkiIhyqymPPsRS//D/rdaY39mKP19wSry86hRX3jK6cEyOiHTKT0YrFD
Va4Zp5uVxU0uVGkMi+sEVMgke6420F4FPUH+UZ7u3A8tbTQEnz0xz2sjCx8CAu2OFTpCEmrj//xU
zZZaTg4x1yxUX5yb5kgCDW2x4mHwz0VRW7ljAJREIg0N+WGmoOE5cNzzpuxKBWDEFnlY60yXETTq
23X5bim4f3CLaCpJLmaGWEb+/QN6/LtWemtjQB3tncvJLbSMm7fRiUMperf7CEJz5reQAA+CyVM4
NNbnSf3rOZOtiBc5agSSyCGOjePSsXZ622u2+H2KN+9OdP64apscENz+YRlnkD8Vtxk40mj8lUpO
2MihUneX4nO2U8jRLLp4PX7xyVzPhUH4cDLn+NR12L/T0ICPu50KYcO8045LWhKDSkUypxGqc60x
Hpfh1rrSb2pNJbfz5BdCeYRjSOHo6WKWUrxoTmVOTzUJlyE+PyQsVCaKE1j+DByVw/Tq6hNygMhT
py7u5i1n9M4oGdOu798t3jQxdb2qIirh0CGO0l7P9zzHu2sudOigqJ0jOMswM3kF8hPbIGFtPTee
M6Ru3DUOMQF/UHm1r5hLYLB7WIkERJd7t1bv97d8pDqXRmw4C8lqiQjUlAPcDMuLPjQaDt/3Dt50
i6/foMEFeDfu7MtqwFjU/jUH+3U4YijpC3yxeob8Hn89fQWzQ7VFUL7JPec8KdnGkovJyV1Wo/V9
1VTxzRU0TJIG6kIRbNOsGBy3RPRV5JKphob3Yg+gFG4VRJGKyByIaX2a+oaf3RAvFPozDHTavwG4
wxlOVTAi38tJaVnmLIyxT0aZmzlJZKUtso+thiFOb4dhg6+UdUC0LTCFh8PVRDsfUK5sinh6TaAp
4GqnOqqKpcZewLx6cmI23fxfxwWmNk68ADacvLwYCxWj+83P3XZ+MilHUxObLQH9YkhB9apit1am
Boeo17oPEyyoYYpJbhcrscpClHLxC7YXFnBu9pI3up/r1LkX5x8oJhPddndo63p/7BQ6RaOHlSxj
KVQelpG+YutphGeFlT4zMPwP4wn/uz8RcbzsLe2C/yZMxjMzyabCdJNJAY9Q1L2IDCyAIDRdvZcT
ZsaMW4ZpJCATlwrwSRA4aFe6+TUpRsGJeP5juSo9PAmcTVCAcEd00t5MgcKA2Wx+wouSgG2b6974
CTSp+QaZNkPA34PasAYjJzveZJHaUp4qjsNEvRIq0kG913Q+5hgO+MKGqf8+hWLl9qdCtxr4Mci2
grNlrAnUvsZMYVIytERpBooPI1fQ69ry3IUwR7lYHf3gQzi3P5QwBvjqmYcFYU+4fbGUYdWjbt5C
99EQbY+BFzg2oLsXsF3eOq/jygMFBRiWOPKlYxvTI2uR51JgpN4ZPIKJS5LUAao+KulZTo8zSJV3
v9lAUIhxLWKLJ+UMS4jA3vcu/W1BlTgQc9PZru/b6Jg120i8joNI2ddoQldmIRuaz5zJ7sRU3n7a
GrzXvrAde2EuJUcKgxyMVF+Te+jG97aSJz5l8n5VnlSbBlfiMZ86KDX7Mn+z/Mx7BOf7CqPsgIGm
Ryn0SuEQFj4kC5kaPQLVgYXpc5iVaY/tfkp7SIZXy5O2nkmmST0o0RPRkRZiHT7jRvrqDRp7c1Sr
nmPRmdIdyWEgrZ/B635eMD4mf0mXupmQUqnprjcKHCRZG7ydEShigHLGb0w5C+PnKSBXpKygDQuu
SYLeiUbknl/uasT6r7AGes5+uFd+vhHawx4idCPxfc143/BK5ONXI2xsIQpo5yClK73qR03w7Nil
lstElmiHqwqR75tKCJUfbT4Bg5p1cw6hgfnAVi0cHNTz3D6VawujaV1meqYkBbxUMxEi+4ua1Mf/
THSv6ckkR5za8lFPNXbxXS8WG9mNxAv7YaEnA8JBxSgLdLy0zJoHByJrSTHEdXVDdfd2vrkcOhm1
i1vcgZ6bLedzrNwSm0/hjUzacFIFglJcH7XRzqLRD4YxBm4ERWeoKLMQDcC6GwqjOlrDOezRMbE+
tRNvForNRzF11JJoiufpuBfuK5pnGziNCFR8s8GNd8/GhtujJjWYtIpCcFUXQ2derk1IFJAMvbvl
Jj/VhXmvorkDasTR/rn6lcsXI7oKVGRF2lEjonY6/nReknNgV3H3/q6flT1to6f1AsmSX9Cajtqe
VlCbLSDCo99Ljy7Wq8UhyKf448hgKhdgrU9hO4XSl7xxM9HIvxYggYOdkTKyyZ/u3pLN8yRF8dmM
BjvHhdRLw95qFpH69S4U5dlm5DiE7+xFizWxEoXqfS2WgHqRz6fCuVIs8zDXEKhYC2iY009Dc3qR
R445u7s2HYoGt6uY+m+DZsfcy6UwY2msMrcpzxPfiV2aMIs3V1fThIGpKpR/hSeSPLb8i9YvAVMW
UJdnoFfskRVbHrYJ1/pW0w41bohwXjIJsY67Ww9Ue/3afhaWZ6xGhBIPCU265aUXQiP9mBNGO1RK
FhQqjo5jj4zjiKEGqzOFHJjM1IpGNQOBywY4dS0j45i70GDYDVUhR407OPpXVUx5XhNQ39GFRPf6
BUsjyPk3okfs6DodW1niVstnfwMLRE+eOXORCM7vHMhxVWnfASENN95Wr4hvQa/f+eFIUHUVgVMj
KvKOD5S2XzopMaQQU6ovBt+zkV4UHsDtUPRx2bwuEUawzBxANMsS+ORHKWv69O5NfZViF6F+LcNk
n9gpj92CHQsMaSx6otHYc3lDF7AoWzAtBHqEwB2k7Qx/1nHStXIVaJbetTG0Y5X/hzdFk0VXnghl
1/RBEhT6L0xAqamI8s4py5vZqncDwKdtwtpFeZVC0HqnSPXgKba9IoXFkR0jMRPEDTy67rdaWNZh
Q8FTJH5TxriWQeTDUa4+tcwpua/veVGaVrbYyedDFi+D3428f3nX3UvEYFO9YcY0gkwgkSWn3zdk
sbLcMAJ3fdGRxt4dsncud0SqIWjqewwCGDXZsOV5bJoo/gKMBnp9PKV6QW7WNeVZmuyMO3FK8qt4
azlX9EdFUB8m21zLv3dzKDxOYBJ4qzbh8VBIwDjLhRPQG/5xqsFctjRxH1EJQSaLuj2LDUQ9oUTG
MJQBbblpsuL0yU6OZ/pHyQwa08Qn5mSk9IEwsSbbZ0NW3NfKSGbZeSdJrnvtlR/FTh1S0G9vYP8V
QSM+TXrieB3soCRumDSx+Q7MKUXt9zkDPHb/j1gKCXgzeLkHZIDjMNecFqEGCOfP5xhvslfGmPlO
eInvVbmOZ7xzLdGxxskTpkhFhDwnx9pBuuoIsr8mJnIfoCKbQYqkX35QRS/Impzyf/PZgeQUyASp
he2o+vxTwUGM9ZZu7s0275gX3lrAfrapuh3FNnKvwwTUSQVtr4+hRGHHJ7XuWJHZ78S/XISB8nmT
Or6RbUqjDAazajQg5yZ/uVFvC1XJ9+vDG9Pj5Dv17nMqRQVbdf9tdGVbs+FvG1CnAqhAKeOpGV8C
GNaao8eJZm/0dfg29KaEKA1MOAs0k17ICkmEqKTDhxK411bq+yvA6UKoioocFW8zwhBq/bgONJtz
aUMArOfwoO8Mf5Xbxj7AZPVtBZc37l80ch9aWGzEjMMWiyyXfMZFNRQpmNmerV/c0ePsydLe6J+Z
BFvtXprlDe+wTR2pf66aHpgvDHo6h+/dXGDhLEudMVW13HXdK+vh+hBsy1FTvvO/MRgAayPLSobs
9j7vhXA2/hWzc3Adf6TlY2CJZsX6Hdr32L4OYx136wKAA/cTec+NJth4YWajDONdCHNaXILRrZVN
kdqmJe4S3OJeMN9cNvz+2In5fSnha1Gm6JrfLySVjTBJOCSGU5OYyZZ9v10PmHTnfQxbzk87IPYr
hAXSHa0saCkf1FhgziRzd/dMUYoELSt+smqFfqWHL4yKECGrfVOIdD5hYApesxBpaIOpChl54wnl
oP4wvp/EMKHBWYPNGTz4u5bEIATY/os6f0R7jwmsS3zaqMnYIPb0fKvU5VT3Yp1s3fpNRdGzwMWa
3qwLrxMo2gwM53kfjewl9ZRjvQAX4cX4k99yjHyYdgi7WqTErn8nCXTL6uuBrIIjspjbbfDmCUQD
z4XqqXkO/f+IhcHDb60h85xPQzS+VGf9YxE/nJSAYao8r3p+NUGOXqANrVXxpzXXuXkHFgDIKBaj
b5wfayVz/qMO5UbX/CHvZsb8N3vBj+U95G+1fb9ojhEV/bi207sbCmmlR5Pr7BIBCDIbFA4ymE0d
qb8rltazJ5VToiFDa873mHont4U8UymBCGReDmZYjqMwKXdXvezgYl7r9rAK1uHRi6ft5xXKf/kA
IXTBdChSywDrVKZQy313UFSHdAISLAOa+PpEyIXnTPHltN4TpA1G2uIb7VN00gPsZXsMKZyp+p21
Gf3xy/etxHbTZMx154e1VqBYyEGlDfTyu5yj6bsEAiky37FA03epsMem5VkAiiaJpyxoh9hs5Khd
I0qCeeskBXA8XvxSl0dF80fZGRZ9qeeLArtvvj67PeUBjxzDCEqRtDamP5P6zN9bYI+uVov9JDmn
TNSCylQZ8RYn8XZnIKlUcwmYKPTVDs3s5+3NFA0a372NfjrKZc5Ddx2Wnp5cg0BzPPNsjCciOc1/
gRq9WO2s9lOoHvwDCxXlWcrEatc+Er8140JS6sNn3nFQ7YiGH7iK8E/EDxxp+JTjzF6Rnp5H0uEp
DUTYZ+CnR1WvlW/HiCI0QlEoGM9YtFQDK3I1DvNB/YLbJWmJvzid4Mz5A5HDYQmi6yx0ImZKYufo
w447WAFhMUBt//cBtlESX/4spaU4tBTyLSsglFcb8TiFSsKh3ynKmrTAzLwquYiwS8Mv/qOR6I11
nn1Lqt5MM08ECDdPLi798p0RysYbsx4Jnd0qL4Hgj1vXe7zZ25JH3Qu816swUDqwoEmBJ1hzSZge
YiZOr/1CAv+k/w3P82ZDQKANFQovDelDLCB1addPP85yT0kpuPr30Yc19BURgKl4a8ke61agafxA
c+311Zz3Ppj5qBVp+p1Zo61L4yIjp+2yi8RR9KYPTgsdTDaW7kXL6V8kLxyqsS+KdzgUC+WaqntC
/v7+hBAD1k0zzW3MxUKhnUXFR/8wtFVFPj5vnmcGobzsnV3Ewz76XnaHnzfI1nM/iXyBXDGzzV55
K3t6zCWu90ij4H5Jxo/vjmDxnwykwdW4JLWelVl8EjeiWR9uE+rPVoOvD0/pSDio9fiNafdhQI3x
bD9/B5JNWxRRS5BLPeqQb6p9ph23cv7Tv8cVJQ9XlQyOGSbJ726HlZYTiF3my0lk2SqVGh8lgVxO
9ub9vVcsecaRWHHr6eSW+reYRiReilYUNXgdEcmemPuZRCEF3mMrapghKggkEzozhIANA0a4Pxri
dyTWxxzXx12Jj/hvLvyYcYYoKEtdVjetlwBCmSiKpelcLDsgwS4lBt+7hvFjHO0SKykn0oW7djUL
xJtMEhug3RtLA8IAzZBE9POiTCq7UhNmcF0z1EPk+/vmbuYpsMIsMOhgGVAc8rpq0OPbGJun3FO2
BgS4Hh72HrCaTaYT1irbW/gWEV8YPgLYn/3iJ6xxMWhVeE8hJhxFRthMHNvnhlTEvhjFpkellRPB
n7kVZeMk/Nl6mBXhwVXfywv+As9RXPBWFIZgL/7ttXbAc1z6N+WplFm+lv1Rv/6mA2Y1Ag95v40y
c9IVMa82Qsh4s3vyQ8i7symwslOYyfOQGGsF646AYqJT6cHTrD0x+1WPrUIp6OqrFwxVg0YC+lkd
fq8yTwuGfMCHVZZiONHBCdWCSAIUWcwcnfV1dF0yFNZk8VtL6/nrNk1EQ4Dh1zc1Pm6DgfZhdagq
Od6N6aAyobzaRh2pU3jJclrIqz7WtafYaG86e95J5vZSn/Uv9q50MQhc8HLYtLZTX1QgCd6QZopR
NpTRP4ZEjHggFResNzJXjnvFKH+AOYnBO3pWsXmRJsvlXTW2Bx3sqwHstF5cU0XYX55VTkMaVJ/h
0mw99gXUFS5YHjBR32PglH3ZrD1ECaJ12eAln+m/Fa8qcYMwsO84+iKk6Ual/6mbANqJOS7XUfib
0XR7Kpqqgv3C98cUq7R/BqVahnYAOBUAAqwlPdNvkf9SrLU5kAc5Zc9rOLgQtFBuH70b6fZbOqCw
CawAHnq899j57C5xgRoHyEt8qTnh56xCJXV70LmqVjBBJnqaUOL5PXPDDMJq/gcYIbgNz7FvnxE8
acsoxp80tyN8gj1LusteIDMWOTVr2bxs1wGWOvRgW2QopDnTaZqLv7cIZ13T9bTEjPg1EyT2JHcw
9oSXwRthOKNoeJJ5mFMjagbDWtKPzsZljB2cS9WD5Ghay3Me9aYuRKuq/YJ5AVUvYLbdfXSLdXAd
3WwYC6/0F+zR5DlLzqHaDXoTDfcIcYfsh6Fh3HN8jKy0Rws+V8NL+meo0lJVTzC9qW9SRJ5ZGra9
5jrJakRrwl5pzBfVvR5rP+dLP11QCQNi0IYQWF3P/kil7n74q83eXDWc/9+HSHQ0d59VgQoAdCWU
nXrhKhOf09KJ8h2Ux2OhRwtUu6Zp9sOp9sJabtgv6U4pFJNOqWCy4DwuTjUqxOvTzbnVrp9LD0HZ
4BlblwWR/C2X6c8p6tECDccygrUDcGs6o1zRZkKbIAYrA4DgX2sj24Fp12zNgCZr0Co3pZswejIM
UnRpbCDE7HKKby/H7LBrS5Nqvd+u0Lp1FTDTr28SAbuXTo5URx13oFqNz4y2bkMCbkPA/85odYKb
4/tf/gV2h24RsPiBvso9Q5qAiprwe9ww3B7B4O3TZi+dNCABy3H/7kk3E3UV1j6peIv/FtCbWipJ
FSUNEtlsBCi5kwik6zHaDaMR67Oa3hH7KHPq4wxEEVCa0SbRNXl9FyI+WuTZL2EPFk7inIUNiytN
PbppVm0rS9L6XY2gd/E1R4wn6jwYyYcUUEZOM27/7AzYj+muXNzlXnQEDKaVSsDOHQjpGGaIHXpl
tI/jxrogxj779qwxjkg0iu9gmninooFRtoyI0EXAAd70KmZCp265tiRGf31bvc7Lu7jvVJT9iJKm
0bSsbMJ1hKSzygR2NM2TQelj5DxH+7yR0PMW7ptBO2GctPRZURJAHKqylMuRrM3MVJa6jlmlkbTv
nNIxI22g7Z1TNNNREeC5BxBU/Z4Btl9wI9o5AfL5rbnXVjK8/a8COZf5RiQYBCewvU13IlPM4Puq
UkcN5K3nS+twRcrqASATCzlQQwdPqaF5w9YMaNl2ao1bSJDOGy8Y6AVFNrSlw8UHtsUBxfEu5vi3
PCZ6pvn5T8B5bARz8E03C0lbYQgj0eyG5qe8z88t+fB5bjebOrT1WmDdrvk92eBmCSl0i95tyJIm
PYnMZmGkrIg6bm7MGMrqzYUTeH73RiQePsC5rbu/q898SfaX7gC6QlD7B8HhUVD3Sr6pjxiVa5LR
wMMaYDrEnbZpE9s+n53TjfQBD4pyXWLN7+y5RroulYacwJCsztsSl16D/BuAjfUX5HfzZI7C53dt
VkVP2cNpq0p5p8mhv5fFJGcCVmr6CS/Fn2FLFFRXOaN3iyAiLKWO/yzqnokqmQPJXsyExtY6G5gY
/0sMjKsvXiuCo9q1uUPbe/rMA45uWdaHqkvwMC/V+MsyRwqCS2/DcQRBp+OJqBI+EmEPRav8fvhf
N94dlcSFSGFPOag1AW6obmpBWQWXj1HQ6eCGcexdKMR3gcNs8Inpzx486C+GBfmL62oEaFrmh+VK
xDt89/5hlfGRBZiLNo5c0ZjONQTg7zS9nuuyGwnOx+d5CNI9LhbdxRQgyrpkHZkxwAWcNV6AvcWr
Pp6eRbUKZRvLc46LPKLrrYrEb6zSaXkHMaGLkPBLg2zygIP2mmjuDsehWMcKgN2Co2/LVVZ5+nPd
XBSGnlnbjTZojJB7Ah1E5y98qtvAAagmdALefdSrw/JffpL7cz4+Ohm0hbxpUOvV4VCjYJppLMZk
4xz7+KvS2FopiZ97AYY4Kk/HVe0iMDdghmQULESCpZAZn99uumKhkcv4W160Yf1bOrD83b81kvfQ
7RUd3OeZaLMP4AnJnk7o+92/6QJ4wdc0ouOoDQilUHn5eEnf/CbjKKMkDg8A4trJx+ggG4G60Ul4
aqBaRh2HSGp8f1JKJqy3lHXBCfYBWc05hM+80QdjgHYqo+roz9LDFnJoDhEvzsWxN3K289aSN7A7
dzJna/Beou8RhLT2lehwaIfdOvbY+PD/4dHbVQGNwT6N4GP75b4cjhDWHGlcDsuOKZOv2efQ96Ve
fl/EF00xxuZ9sTfipcwXQPMmGWLZjXbkT45MSvDEktLrnN8HzJsfmbqlKyt05yPh29H7gR/4nYJo
Rkl3YzjoN8c8tmrwVTs1SkHBwdphcezANObt0lCLVdP9DvMe76Az11kXKKbawLNSIxbEWFSh8LNl
V0MnAhAvv0lL1Spvjsth4BIGpvEMW0iifrUe2jKkEPY5gZuKK7S/iwVbf3sZvUBc1M5Z1stUuBmn
WfzwwBUMBifJFSzVhhfuVDViwfBlProR7SyafcPBES1M2g2srspsBGr0RocU7z1VvfHOZGKEQWQJ
wdZ6G8e8iIXkg9WcCr8hgZSRJrf3P4X2VCpsQ/XYzS0nE0T/2DAPUr3aXYJVUonYQldMzEhlol8O
ddsMKx7Q/TPpmKwQYRHW2E1E+/HdbN/XZ6oG7xhJmdUCfhK3kog8pnTlHwzBqtuHVm9jD8ERIWcn
eOYSgNP2tDyUs2RSRhlwwAOyn/LznQqOzf7dk+Xmi2cJgpItk6QQn3TSJuoHTF5ds19BXXU4BvOy
Q8G2nbYJy5USLR20r+gcYoL0gHygo3FX//bRLQlS0jgVWJ1FRG6GlCr1OZP5pOIDZU9EqmLagDiO
73uRGVwUm8SpihR2MQ4yZEy8kHsKjW5aE4m5TV2aQmmbrZLnVA4hXlF3b2t0HKpFiRbM13xhLvah
8IQFvVBX1pb5RDGgnva5s3PF7TEsS7Ozz8YfOUU5nOoG0YFOPwX6JVycfqX0ksK0SGapLhZmoGrf
rLdMGdENm+1B/vfx+SRqYkVT3598F5Po01ENwWmMRj3Ld2XHROdZe1/NgQYqV/peUlJBFXIM7ztb
9P4Ohv249RekxyFp8VEk95LjGB7kfloPu0dZPZUDVcIX+hVdF8dc5TX4Z5d1kolzEAPOZnbW9pAR
LBkPOcQwnngIChMxhwOOL5I7kpP19DLg1pwh3emozXT3ji3c+fVhrplbabF0qfmiEy6ByELeee+N
tulDRZB43RYahPBmW61RmDL8kS9jTsKOmMQaS3TGhL4HS1dlgoRbmvS2yyLQy+yjPkEMmfgzzNPv
Mtw+E17VmjXFQvSsUJrgzS2ZGvx0B/56MeN2QxUr7dv+id6xJF0A3oKRafsvDS358gAmefg/7LQ+
3mXEzD+arAQ/x8fKuwEX70+QPZi/K+IOxA/8JB4APMKq4gAhkXIJ0vwscWT4ToR5UdhzvQSIE7Yh
ynCRoTxkBvPYOf7JjLTNwqGo+XRlq8TGosZfqKqCl931pBUeS2lq/iDK/Thdzr2hWTMO0oGbTK2I
C71dhep5oDLtVjrZZ5L75X1mjuy+Cgjpy/xjd7qzUcrfXGfITtcRBp/DwNWOGeN3KsuB0U4FMt/2
ypxrZDPRSLMrAZYFf0eSkHRcbtrO2apyXsMbPvHH+mQWUFx3zDGb31WzcloFClafmyyESFYjQSeU
OXWlztpZO/NyE3Tknh8Gmarj5CVomlIE7FQYd2ubwp6SXKl3yOCZznessp2UqbeTbylPoPPyHHrY
0Piiw+Co0nKpyLovUeXzPclQjWfmUwFG1YppYi5D0Vdokfi9jQ3hswWmj48UgfyD03C8ye81exbM
6wzIS9+8ZTY9jJgP2D7NzmHxwKbNzcioy2NOBOYhWvjoyL1dCwcMXVinC0VYxLn+gWyIp0mlERtZ
cK9E5Wb8jHtkeBz1YufSvM5w+5dwESAa9I/KjgIL12jGKuDY09UDM3BPPMtjVZrQSIP+QAFmqOA7
k4kXmb20xlnOrh3CuuJCEspjsnoCf/wZQJZvL7922DcHrqivBGkUt0s793ofse9sfyIDTJk0ldZg
oWz4IWaOaze4O5rTyXX0SNH+3i9+4DHPcfWkIfYmrHS6apRPTE2pM/K+M5t32FPm3r2BoF8Sg7nS
Q9cWnEWaJW7fnFnVStHxktffV6li08oacZWZEj95/oGW2MkzMZJWlI8aoyFNzO+SGId/NSTLmRCP
1hZB/YbsnfhFAwas/3H/gud8SIyE6tBK8xeiy/3K80mpYLfJEr31doUU3lfx3k/RToZPE023QX4K
MKzWZWBTfggHz6lHtexE/fOPRykfkCaR15ZgxacYqqPyuADDs74rnnrp7k2DbTBhflNXNIXPbYWV
b8O1ODA9IOBv6FMwddaW3nQHv4gmRYwh1HDrgMcdQZcpBM7fVpLtPVa2cvT/GxGwIbw/yvjIVX1Q
Jm/352iuYrrQFr1SUiF5HtgwBJjNptbfqptwm3DjHuSZVmhCkhc0ZoVrh7MsalwxGjonH99x7jL3
irLlTy/F//c4TGofOqP+VZi++jzVaDy+0WB4Nxfmq1CrO5Pz81Gx3L5eSiPzhjVE9mfwoaHoJb4W
ht0sd8SrZk1od8Nr2Tk8eHpv9iCNvPEzm2cPRbRgaPj48Ko3Te6HtKsePmrXmdyqH217v/4mreKO
eKddDhMJwKuQud8xtVnkpQyiI3faV0f7jbYW3E9QYrpQM0OK/sZ7AcmifsGRW5rZfwnEv63m0qFd
rixVHSFcBXiWG8036gi03rH8nzFaar1g83lShpYzWVNUVy4YBJ0wlgPvXqreL7yQRIM3RlYs9/q1
OYIEvil2d++uev7VbJOYkivLTq/9vjL0USM9PDfVyfzGmTkUj/FkhOhSBtRsh2s/oZBqfz4t1IfY
JpJDr54cth8PzJWE1sqc8c2TQyVrwho1aXfXJ7ypBTbrbK/V1yf1kQc5AvC8FDVNi+K+Owm4qHfS
E9BbSlS8eBblCcaqkKyb91y1Loodjs6Qc1Pge8z/piyyTnF9C+U8vjA0XcNC6iLZWJGRkEuzphqW
mYt6nd7yZDdlPZL8M0MjYp23TsuBMwofhg+vu0QkWgVj3tFeHKNZiom5hZNsjO0A0TuQGfayeIyy
jSYtP47q2sRH5bzQmoShDDzNFIJsZXk28Cs/gP7/QPCa3uUA/HhgcDIU5B6dHxsV7EerxciWtmKO
EpPwZbmi5qL4YnALnrbdPTD8PBxJM5uXYXzibnls4pttJI7UZzAWQSDpJNxB1Eokq1ag2U+ySCmy
cpmOd+zGDtVBlRv4PFcUZA4/RD/pO1maZ3jZ3NU4kPZtR/c9vh5SKa5PETJdkZw7//wjIWufPi4u
+1Op7tyOEs3wB34hOgIFMwPq4qW9JVZXenbDvoIGTkl8xR8EAXTGI6FK68LZXnO2jqLH7EN8ep4G
Ahv+3BZu7grM6mXnPmtIWVifxK34Z9kxLy1vyQluy2IcRAxlgQHeCYZkCa8di1AEGuBO9M3wGgOJ
ZTubjmCwXb+QKS9+0brIitHbbOnQFI7YJ2sE9dVK1s1/phfQ/jTWmqYU5hqYHhJ4y9z5IgOt7Fqi
DnRLZPAbiD1kWi0mKajNXIWpzyNYeYN0eY/NiQ8fB0NGj3+72RuqPiPyTbNb4MvI/PwzfOq8qR4t
xAdiiHIkXJqodoGn2GwEmZ+9EuObVFKs8b1IVlxZW8jqX6JxvgUe6msm6XnjxxFj9ENhFLzZsu73
Er7Qreqouo76QgI/SaPaN+P6zzvikjKXq6C9nqVVygXz9EXYQed1d494d699xnHdzT04y644/VPV
GXH1cisiL5saceLMtKaqBuYYubgCGJGI1wgGDEDZIfiPafsWR3E8tQ0ENPAeO1Yka+YYOfRiaMDu
VTX2V5qZGky+010PkeJBmYHusD4v9U5kWlPvhBXmFBnHCEFTDTnwFxCONgffVHDHb9wUuRhpwUmH
+imz52DpXd66sTShs+7gzCkTtIvuFCvU6zFneOIHZyWogVJaH+Doya9qzoPj0ibmIPt2zqx9yGxD
gk/qBCJJ/TAuvvfTNne2/g5wa13Xby7kY5VzWjFS6xKVkYQvBTogpmCTyxn3Fkd0lRpLNcIErOEq
UK8F7wZp7OjxgtDl7bQKcxtpCu88UapQEK/U86g7pqtu9urcn7DCLcBIt6AkEK+Y9BtWuZvPxl/u
OHsE7Mpn0VN6raTI85/oq+PBda4s85oFn9NsbXNahQbEEuk6R1wGnbPO9y5d4pG8eFiLaIF7yYyh
VK75doha0aKM2Dj+9HHZwxaG8iw2kVVsaV/PlZnuuV068yxpJkAW+asJSlIrkncnXozXoPtoh/OC
3bcMV5i5FokUj6zPV46chHlIFQeY4WF3BBoyZcGxGrI58zn/QHf9Hw6CrhFxAa0KOxtN4lFxgGQK
jZ+hxw/HcoR7Xnp4jl+jNw3euEZwu1wMDfpSjzhuMOehDBFQ2Xsky+k/eX3l/MCpIHCXT9H8T/dk
X1qt+wORawMNpGZ9GydVE83sY8jXus7OXEwhWukp0RE4jESMKbt8VnFyZGV6Z+IF1WeFSmTicpo0
gcprCHEXE7XDrJ4QY3ilJ9pcKYV70VwvTsIcCqaOwsXKY1jk5IwhQ+KBHLV2UMUyY2aBWbi+XMQL
2Kcq9PMhjh5AcWXhTRergb5Ail4+NIs8Ayy23cYqaSswk+3vMyPU0lNUaINzb7q5fweeFpbmM3qf
EGd58bYsM5CPDXTdXB0GB5cc2r0KQNKS/BxXqB9y2sni1JZ3DRodBMAEOFfeCXmroB9yGzqToTKh
RjTLVx9PgYIBht129TA44Ci9EaeC7alvhJ4Uqxcy8wRDRKfllFtslpl13m7UppYVPgZ6aLVrDN2h
MidQ8BOSNAYGjonD/Qlqcwej96M82pjLwUP+ZoE62fZV3HQmWlDcb3zpGWagVYPYH/6MqXpz58aJ
sGDlgzahy7lE3r0Y5JLmujhYOivvrB2NF+ZO7L7blljnKrOs6lEVPYtsXpC0bf84Nq/xr2qcZZcz
JikBtx0gImwRtjTst3INZj6anEUfH/j1LzgWU+0N51ardnRciXC9prwWjGKxS2xJrS/IgeSpgNXy
KZlQSPSw9YCEaspLB+j2BftSFwXJzpS9Td9VEX7zGcVX9toEe2eleevE9d5DBu+4jxicRn+U/ZUg
D3qFDBS0VfmWBS+sYcRcoOCQM+xLVpvE7iuMg7fe5pO7vKYFyFVRjNRIcLaLXuXoqzPE7lhw+XWF
9SYGPwL2RdRt/Cb70AD/H9S3cvXOwhcd3rYlp98gg6yfRFqCBKwvAqUzEUyX4fms6Wlybl3oLMtE
OJxZA6zMNjVha+o5btOA7u1ckEsVfsn3vhDRBfCRwvqbuqXCVfWapMdT4IDxpsfi0SMqh5nKvtHQ
nOxOU8MukQ2PpBPLbIRcc4N1g9UkDUjj7WMlkERPa51eIJmjCUgLM8qLaH144hJubFzZUXt1aoaB
hX7ZWecXDinJgEP2pmvjCDe0zfSRfgeLiMJAgJG4S222vmvkFgawGdSfT93fBFwpyG3OJs1qzfJf
IAv8tJs7eT2i64mODYIz2D1Rb3wFzvsmd5TDA2N7HHIrF6rwYWH8R6J4nF8EDJXp0XUISB+WEkNr
CHBrFJT9QWyPZI9cVyUMQ3SzXI3cZlySju35BbtCkg8k+RIMONgTEjAF3Lk3dOrCOokTVKzxdsb5
dGwuK/XQLTcD2AkvTgrHh1ZaIwgGrTZRuAPRvNDuZwI80MilDO3U5XmUIGSRGGRyJqdDauNiV0+Q
tgHmOExUIOSQ9L4tuoPRf/f3sJppi3uw+DzkH0mD2J5aVVdtbLAnVDsIUtnbZKu4X2Sp4FT/tKQD
Vd5UVKy4hdJau2LpE98f5V/iRNyPs4+Ar946/AGnHMMswxLzU+uREh7fr/QJpZ2i5Y5Ti6vH1EYF
mEyBbFU5EALgDoMbKXqfzOZsXP70Xg/YwqVH6Zqf3hEZcBAW6Iu91IZGwA9afqqhTJRuTu+14T9x
52y4Ukr8Dl4QEm5yTkbL2hjuVcnHkyy8Ga2LU8BJ2m1zGj3FXudUFVjt2whdl25iLfjj7rQH7UcL
HFNVvPEtwTe2EP63+Nvc6iWhF/Ajif8wmT42xAGQ+WXf+D7qxHbnvwcoRdMi63wETmBcS5rKMfR0
jnMX1XvkM+iUHn0QngxgINV4tIjZbNAd4MOnefuDuRahRtHYWcNUBxIxja+3CKA69aHVdnXVwhWJ
WxmmU6WuAhOvGgKNv7v6azOl2wkT6p/0bbW9lmTwRI8jJyPFhhUzo+PtCdZIqIXcAG+0zZc3dyHC
5lVlxkDJbOdjRzAblI5n21YJFz1h98k1JCUBpW871ACHPBqh16b56an29S6Mxv8l+/RbOZwMM0pB
Xv2ciIr510tjBMemm0bx8IVXsWc1EKTjFN4U25VGP7WUhTg7imTpVewWE09rfoXrvUaM4oUsjMVO
XosjPm88f4sFxgZkbFqKumZ7gi4Xqzpr1alApRS4+ikBA8FDdm3I8uXtbu1W2qoS7QRlviQ08WGx
RPq3MhEK2y8pFAryxf72fpO3/7mCeQRXfCSmOjH3JonfYEq68WkgN5hEtimtto2vuw0+NETtFptZ
dT6nINK1VYNhxDhgyfqiTTzxNrPHI/kz/PSJ/I4EOsyz2tPUw/eLyE8gTxV1MI1hSZW+4/YM+Ow5
/RRFhA7b4XmTxI8ps2MKeooen4vuiK9xhPAcAZVOzK0uUTDdkefV+0LHHIt386ZG8yaKaSWoyQWa
HwaRLF468MeskDbJ2jiE0rMtPw22OduXN3hwGpkos975ioAKOk2+Pl5kJ9Bxk9pJ6uWYmBmN777n
s/WZ1T11ANGkgFoMCjiXp1ic3N9l7Un8EVhRCkUOPpyk5foG4HW3iNSgi+CeMjg+X8ecvydqiSYH
Uyda83ZrfCj8NkrLDP2zle9WpTQRgkzOMQmOLR2a61pRUzf2YcQ+ItpQJO0Ptpm7pwUDUhv9iZc2
JX/j9pfHSC31R6nagcTs8hb000DcHDiFjOSMoc3yB3dYHBsEb4KoBr05Bf//ICqqsc89P2tr2pLI
oDdZ31ghCGOaM14UD8tJwquilrrRkBLFaapzzR+g3tAu18yCd3UBmB3VpOecxk1CaEuDIZuKUunW
ojDSvmcUBELTaYy1CVUjrN5MsvWzY0ALayklVT4Dz2YLiC3SCFQ7V4L3E/YiwBHRTIBNrP99Goob
/yQeZ2SdLD3vaymbfr2cHoFBEcpNqxA8Q+Ud4wXnNuQGv9Mof6dKH9LY1Qw5FTUZIwxXvg5ZPHKW
u0bJNAIcFbUM2iSVDeBoeBP5HlwfLIjVXSTVMRoB/DkeE87B+T0aogs0YKMM6eZ6z0N+Rpl1sMeF
AThv5E6MkVEU+gL8zYIZp3iZgZU4NBZ5GKe1sfJF0IkRoarFcXupKpw4T3cULK/MiIa+se/N7lF+
GljpjS/646uA0BAnuPqxwsOFsMK0wqP4oTKGpFeCbIyV5aqPEqhbd3jVQhEySJR2rJfXsmCOEbWb
u9r4MnsE/g6TsbyXrxWLuKO6CrGcB5xSqNRt28K8jvymm4K2dVUKYD0Ak2+ZYY3FWEYrpDh2P8qj
F69fOzocfIt0y85z08aznFTh2+jL1l+gU9/3RagUzesnE5Hk1U1FgoJS7j19DWxw7V2ifpopxZa5
4Ve37qyCov+4nuch+zB0ZqOZ/pENHYb0UFeHUdmJPk9Oz9qlS3nCFUK1kTL5bgLuTeZZFlLl4ikm
6++cbEDqAhhnFaCTP7r503ku9pxkwWtkvSbzQLsia1ctJKR0kQOC/aLmk3z/wJFpS0CCfhJmaD2j
0Q5Mv9UW2BZ1NU26F1+fyQJLtChptXtExmyp6M1oHQcmJjDKVlbj6HXk5cG/f0R0uj/ecRNWxL0q
aH/gJe8EWPgYloAq79FJqJ69385v5g9D2KyaGZpFV5KyrZ2Qb2jzGqPJB4pNHtPoS6uqdIx+RBl2
jB2vGxPEYMHvNSD04vZcZx/zesfksa1LM/udd5tQ1bfLb3Q246NRLPCnR/N2Ug0ENFte8KIH3LnU
pGT+2nYCluJfRoH12jcQKKmUz1O6zWw+jCI+b47KUsjuwINoJwSVRW/osDhmhlN+CfTqz5a0q2rf
83yBZYdZzVAARVBVnl9497L7F1W+ST84WAyVPAf6cv9HIS1i28k4YEXOirQgGBItKiQK0IALz89Q
oBfs8kblijykFvKsVl6qjCfQQlnydtFRUoDAVSMNLTdq01B9myqZe5BbU7nGvKEZ1DNuD8qi/W/Y
6TSBVnJZa9oLfhnHd9zA/4RkTHuooxJP6336Wg3uDgzGpulqk2U8l/ECYwxgsj7dkrw7z+6rfBxR
O3A5+HOAH5GMxB6qaKVpIhvjH7aG9zhbKNISw4OY0bK1Kq0KrInCtffTcLaGBf6Qoj7W5VggtLtU
rDQzRtfsmT85fV+VV9snbq5KwP4ws8XVI20Dvg0Rb4mhMojOz10qXGPhan9iBV7qoY/st5g7of4R
U7gHFA2wDiFJthWwAmC2AcShD07Qf7aVLkTGKskqBim/MAZ3OkAvxtrvG3vfC92W/r2i+kxXl16k
e9gCvoZA0KIS9go8cIGCYcOK570mFnsuZy9cFyiFu78+BcxFyCpkcaT1YCousr45vL3ZUJ2AV679
IdDbyS81lOas7CxUbIdQ38agFLqeIaEh6Pn9OEdRvFk+tCasWKAlJpaM9Og0JuWAowzg83OXDmi6
3c/sEWdNMF8LpVF1RQtVT7pYXxqMahgrJvhj0IN8mYPRxopGJQtmOOuLzXu+9j1h89hbO8FclaeS
89wztT8WUV24t9C5VnywIBFtQp+MFzlX3o8SooduAoqzYI5kgSOWLwYqLPYYnUpXLRZRttAoWFjk
Y48PPVuY90fo/7Y/k2rAeCRfk0ZNOUdmYZdQW7C2P+RuGpRPWvDc9QtshTbtXdw70ObhGwQrVLog
0SgmLwa7PaH52Hm6cRBTAa9/c8/++r0ns5VTX30Z/YQn0v9wEssVtav6h12DRGVkDDD0nS6zd3Pr
PR94DpubliSsxnq80ZUGn7LTtnhEU+R8pG76as/cW9S80JtaxIrPmrTpIZfzJ17gv2N499nmwabf
fBbXMeZH5lyScItlMiCk6Pxh5z+SgkVfJVgokXFmhGfrvjJW/RYmDXgQM58PXqwPbUCWmVzLkIJS
M2g50RTCWvt06XO+oe+m+ba3+RWTvEDd6FeQuqLOUPGjIzQCR/MthCVjkIz+tESljuRBBMyrDthQ
+OhB7T6ft8+YOAujhcIyZPMCdHOhZp7QVllQn2e8zi8byd0rP5p4GOLIe2ALmA98GzAKjDa6jQI9
6PamnpDg4hfelzc4fa/K9yMAjQbFyxpmtTkpnRCCjqRyhR7p1ZEO+RSk3D5G5u2Ai6xqmPp6wYle
bXhtO1HPcW/O4w2M+D8Vugo3/6guw2txi+2gKwjTF3293YZWfuOjqm62TtvDWJ23kg7HdO8yvG8S
uVWnLg0rP0Eu3NGD2dYtrVLKtwvJcL4erC3gQshMKSn3S5WxCeuz8/ripnvDo4jlIibRb+/uWiKY
XlTnQFRYS6JA3GhPs3NRauNsESrbB4n0JoNNe/u5pOQrRk6MwZPQFoPvLHN+URRmFxyfGi99gwy7
o41LrRSG9WO7X4Uc1QQHDqiV2L8VuU194SYufhOPPQRcdWseBzN7vVoiE37Xx+LtgpUi1G6Q1ZE4
KMJICKGptFnts5TiS2HukqexrJqDCIncdp6eMERU5zXj9jthfAQs4wOSO55VFhwcdB8D3doNkyoZ
BNCxbbryYkqP609XbEXFaQh/1nYhgFlJgaVc0ErPQLcOvhCwv5kDxR5Dsgp8087WuL0QuW+KsxtF
4bqiow3s5/T+NM/nubZr0iQZ/p6HJRVZgpOIGg4XUBdzlOdHEh/KGD78qZnir7+gM+vNcIfxkqhK
GnXDFJiNa/ncd5cRRrJffb5STJdv/LMVnqtdvsN4J30nJp7YJo5CNCGT+f6Orwiq61/q6ojbeDTR
DQ0ouN/s6lW7i9WV8e3LQ+XklwGy8Z3IG20uGSirR1Fv9Xzu6yuN4NlsBxhkIZakSnQlx5pj5fUg
qQSF/PX9tToQFovxvspf81v8P1dgLHxJvYpO8VcKiFtyfTYTJ7dHPVki9WAt2sQ8A9m+VpSFgn7N
P3p+uYRF1m9eh0vGZXDowG1CSHoG4IYG7citUiS3lh3e/pZercwAh+cLpQrF33kvWksyOjaXLpdu
r9ekzODfMo+pY2FKJCmoufTRSeVQx27oIu22qohM1SKV4kgV4bPp0GpmU+OOagsWtEW15EGu8ImE
sSBZC1iJgKQ3RAqQ9fHXiSVpH1udngsc5mu164gTLzrKJ+Z8Hu2+ODp8ye+aBoQ/qMYKLbqGxCgs
R7otHeNdCx8EXg3ZNFsLRLJgd0QZMr2yVDr5dfv5DvRhvGDem/bk9KdDH5ixwOpeHvR//NfInwUb
KVZAHyFb5Ot+iRNAa5eoyaUvdKGyslyi61OyU9UB9p2hOnP/5E/hOtPqlMdjWQmJ0YZtATpMeyWC
Q5le20kRgF/ogyVrUygogsLDaru8//2FZ3LvpgPq9aaPdOqfZN95rWrUkya0uBErfU/p9Fo4mQI0
6bmm0U9XU0OzoyUidE8NwJrqRUCvp1bBg02jinsY0g7VFemSNemvQKENn+dQtvY76bD4Yf40i87o
5UWIYfMHnh+lRxtzUWfRakgKNyVpymfffVRSKKsNn/TbuuBn+AIj4IMgJD/Eh6EPW3kaAnzUg1nA
cfos35bfdcy66Jt4rYCNfm2amqixBIHz1Om5QJxhiBd1+eU203R65wR7eFQWJGfzA+dHfo+RHORk
oRcaW8C27G30g+4aUUPOConRz0gLvyQbpa3rV96RDTr3gUBSCHCqoR4w75GgsAmxJ0bcxa5aaEXH
byrlcgJ+hcTe+A93iZzBwCUNtZLNkcUQm8OOqyjOyBkNJevevHskBDTedJl9fpunp5RIb5fmBlcw
6/M4IsJUCb23Qsg+g/39E5rOhIZ/Pp3FnIQbT7e5X5aT+4q96YrpC9hkCNZuySASTqjkCdB/zdrq
yHnbxE2EDOrMRBBHfVv5hPr7wzK8GxjXnwwbk51MHkWyclt9rdG1c9hkH4N7reM3AguNVN7a4FzK
7q22VNfbsWgWO5WZe+bLqPToJhsjHruC4L7rMrrRPxWLrbnA3pQZcPPTYCXFF+W8lrowMn5ZA25e
s9eE7e0Iqouwr55SSuEUb/ttyS6DCT2VJngGQfp+G02GslwwLTXYQIRKs6EtTntA7Olvu7uRRY7A
d132MwltUJpFmMp9guPTI/+11zkpGzedAS3HT5d+xhiEZho3oupdNkFhZpIMv2LY1tWqBJLj5Jmt
1jgY008u1/qO1bIKmj1iWHTSgvjftTuj1/Jzp3lK2ybW54GwdG/nQpCtcNMjLQwtMfn4ORgikxtf
gUmJU8Q/bTezEHf+6xGNlM3oaCoXO2dfV9Hb/EUr8T3kjdVlg/NnywKCs8snsGNGKVoUNA1+F7vD
caH9fcJzKo1UdXxSUBQ9E7ggotPRKQx7uc8JwjNVrFOCONbePDDwwhdhxC/bLokPY0mO1aW5aKCU
eQqlAZMhm2IIgNurai7DbXyqdlTvktFnwy9wuDG8bp5R6RYehC0X9UG/jstXH+feX4Q1ODdXtWAS
DJMKV7D8Mx7XP1qBV20knlKf3kTknBhg8MSvYadQ9mU6QNKZPyfUtrbIgFjaB9mo2BeFBtdOQUaq
gVdlpsSfaeWG1+vuehMb+bj2/hrHz8GBbpQ1Y59rO+9M+ABeWM6AK9gEIoGLTbennyU66wB/yD3T
AaevRm+xIGgvLGiS7dMcEHgdqWg3RP78npgrHVA6LleadspahE8rowUIHl4+6pPt0FMjP2hhojZP
b6p0kqLydpjs0cy/nqvzlQCrZBBu+rEyVSzfMtMV391Xw7ri9tlCUuhmH3gfCizrUAZfkSIPCig4
nrrPt8G/LQGxCuWrgOLzQk/AoGwrl3pm3t44kMqnBhOieCjK1h5VS6KjJJ++8kb53o3/SGGsQ4Xd
uIxl+Z76mbYCMUU31R84wq3Ii8BeX9yRhfpayKPQIb5Fiz7/Xp74NHunbqE3CnOP9jeAZ0fM5QBr
kZ4G1j1HeBPOvmpWu7R0HripJ/vonomXGYtZk+13ObUStx3cLckgExoQsFtoeKz7sHm2Wraj7yps
w70PlWspfZ3JW8PI2u46OR2REpHeWzW9rzmADrmEg0EJCGqt30NfzX97tBj48JJ94jinn0CyNCbX
B62rrDqHp4KeX8nIiE+YICbGeT4cKiunI8HnGZQeTXVLINV/tIVCO93ZGFbrihER0YY/7Sge4eK+
HfMWa33O91dAIJwm7mFt8Bc5eqb6N4sFEbFKupCjtAbEqKLW25fKX/d1VHep35NaKMK9N//FmwdR
b+Dw7X1rYxy64x/zSMkaWMiRg2WQDpM5dAyCb/5pAFuqWJNLPqnxhiijBJg7LlxEwrxIuguOL1TT
ERzRbfleGEEnBblIhpCL62e7DqWcNQ8evwB3IbEgk1eRsmKbDUpLcYeZfYGuYxmVxYaDrtvt2c7B
1GmGCZ5WBQRmVBCklq3P5LAW0Hypq4aKsi0fK0S2PeiVCSMnigh/VtxPxQ+raFr2gdSMy/qxFztK
JT6e/MxxPIthbvLo/Km6KJ+ODeCjAM2srEc8ilUGy5aIg0PSEttUo6t65Lm6DIu/HWstltEjjdRp
o3JzJFXOSC0G3ZB8HT+o+JwY95OvgPZON6/PZiMObbC1VDnVQq1Ncg5zU7qglhFnPZ3kLTolBBkO
Z8N9dQWwyW7uQu1pIV9OyElcF5hj0yEpOpqC8f0afrHKR0VXxgnRoB/yqeC8hn9ur3grdOtcJVxF
iL3zJqykUO6wx+vWMjOdkjwu3wVoYFoX2UHrOx6JNN2X9JIMmTAdY0CAZZ4AJ5mDgEUQxQ/86KNV
7jSxPak9vxws93z4UJKGooMofnQTHuzfofgQ163dymNw0QzCwVjZapyXE3+P8lOUGCSJ4N/edh4N
OkPcQp97P1bAR6kgm5/GVBEDJTkMTsZNhmFLtU9vkB2l830OpK1yVC3B/LLg3o78Tab0uz3fr09q
iqw9NDraVnPeL8NU/Zn9Z6ytZzX3EvEdXukkrKmDjERj0nW7LfJ6RMUjV3SRDwfe+nwNsGW4RloX
NmuaTNAJ3IjT0cO2Cnj59PRjOCfmk9YQ+BN31WsRwLCR7mbpDZQ7o11aayow4JWNDgKnqeZqWYUw
/VClqHw0ajIDGlzBqei4fCCvVe94pJY3BUzLgRrl++H+m60t5MwlIsudany5s9tHvDtkP5GUuj7m
vMSAtzLXX3GfvGsiCRrU7sF/MwdZIs+/9Ay+PIRq/XKWgp+ELFmu4VWZbfvktvzpYs0rz7Y42ZJ9
6eEMncLK3GLiSDxhz01fCrd8/gRTlFJiPW9UdTDYklPg1pCGbl8rsJRe9pM2+qmNu2e7XZ6Aa0zv
qHjo4ZJjjtatl6hyrmkY1Ty3ALue9UoIr3avoBkuIq5UNfS6A4qI7Rz7TiNNWl0qfhq3N6Cxpiy2
g5QZgyQkByGVRBXi7lHFDJwu57Q4oqt4YUYukkMuD2X3iuW32Q/ygmJN8wPLbHm0Mklbqyrbp9NP
VsUlAm1HtbpcFDh9fcUgyTR6XajlyPe0F8itB816eUiXvVfU7elDw8Kf357hsLVd5TRWspkLk8vp
fHfG+jYqWpIUGfgAdNL+trm4kJWXkFaPV03uEXcLLYyKklgb4VjmusKG1XV5TAwiH/t/8ic8rHUQ
aD1pgGj7hQDW7KEuwWdXCNsK1yMt2HYOF8xBNbWUKRSdYa4w2+ARNakG97JNi/2F3klu3CXEA8SN
8kMKZ7PtlbnkWN7PuhtQEMX1lgimI5fkg9pnHFTAECt4oWDxrRI53vWiACQivznkYbymGmidWEc1
/ENHNbGxAVDrRDCioIf442buSSmEd7D4Whws/fNH+zt25+bDwTteOOLnLMXNCdq48mvQJdTvWEPw
daMQo5kTHkRZMFVbx5+b5CM9RxyVL30DC2KGcamq0zvltllWRJ9So/tem8k9jnpKpSdiXbyDHyog
Q+K2Mz2jFRS5VlUNXYScEBAxKKF1u/jT7OPNeTWxSsmhk35E1rzfq5nn3N4FHiF8N5dd58h6UYES
aE7GRFdQnKPvyO1Fl8cyw5GFPGSN2ZL44ovKIv4XUvvJD40XTBwKV4rJA0jrwIw1t+Vd0c85P34l
xJyadj1P79WeJ3bIFybJCmblFPdMjPobnfVaubHVE85UMegVBtEz6pttBtUyQWOQAaCXa5vYbXn1
V10bdL/bMY854v6JJp4f4VdaouxwUOnasIBl4d9FfFk3gXdaZSdxA8n+6ZCWK9RkvRUT7JYz6SH5
3Bhg0oBByCmXwva71bB12DYkH+CTgFTGhLb+wj3wUWvjm1sZaz5fO9Wm16F//0Wg2n2mL8xgk6U0
VZFjK8SfVrnfWBQRc5xSbG5M7ccxPhm9RrSPD97ZEON8fJnZq/S34R7sq9lFqU7E+dlV7t40iidg
m4KVLUx3RCNE1c0IPKY2nKI86SxAFN/1cHaavOEccKy5O+AEwCmvqphHMXCtR1+pbuRGYwG8mDWz
z8ZtWS7lOo7DBiAUn+pLK5uY2oCu253BpIyVsu9aq28Dt4AwJlUe8/hfxeRcnh+nLCxIBsf7zXBP
ZBeGGMogfhRd7VfwqRTvhCuCaRrvPqBKSDm8mIVSFbrLXGhRcv/A5Dd2MtgMBXOm8cTyHqp0Fuig
WWy8T6w4YRUWZSziLwHY/+0GyQ+5BYI7NMxB+81iAXSn/KQc6OEVjJq3WCEXVANw6fSENSMbbeXI
lxAmyQvYYwoLyh8xT9FUMnUpB3r2+pDVq9thGyK8qIMTk2zZc6pqdXaVpJsfxQimgVHQSmqaEeQK
zKhhkdEEx52umJ/DXx2Osz0abA+FQJzY7vfWywilTjcDEUsL2jf+1jFt88970RBcFyJdYnHsquUr
MZRhaV+wUf/dFHDzEEOXIYJDOtqzVCfIeGth7ZNPOkcTjKIxpVX4GPceinI2Me8ORznySn7d/czb
RocFUNGdKB7Ry4aopReSc32yG4ZpjoEskCFP1pzO6t6fScgvDkxXpiIgKkGh2eSJ8RpQjI2Qr3Iw
ZQhNLwE8A3HlDS65v6jR+6/a9IjQ+nVy3xw8sJrj1FtSDLVHuZrrI37yV9UUYFVo8ZxgyvE2g7jc
15BhGZn4WuXXiiKEdtNjnPTOivCFY5S6ep81PewUnBwU+nAz51OjrEn9eJjMi5ZNVQgZsngkxb80
vagpCliu90oOXE7/N2CJwf44GzMRJoH+G1ombcDrPUlD5T5h7ehUDbaH78jldrMEypE612G3a5Gd
/CjXJX1XxBsusSaRLtLxkqXY3LknVjkfuCfqtnQNOmhDehHfRLn2itKXjkYxrQBRBtAhzWBBOvtD
I5KLhsxlQ43H8CSXcgukpUuYhCM7wzwa9ibIFTA2KVlITZSePYtz2A5Hmdm2WcMlBaf1uW1sPrX7
aVORoc9ERRCtlGjgkAhz4W0aMyGaK04ojBGqxzZotMTUePRRHWA1BufE4p6y7jo6iRBMVPk2Bp6O
Kuurec8HVre4GA7J3f5lGDdmxEw0CcQt+fkRMR7ZjZtSo5SgRFxlTbg+46K5182qnl2nk8Xhjxfk
iT51t8b0WSBZeI9UodfQiuINB+Zu6aDwhbgqmAUUvTCNVKdbFmojQ+es7luzMJxgFju1wMZ+Hv6B
gv3blJipRiOY594Fy5lZIBs/R4MkrUxxn1ykNotCSMRHo+xFIZ4tpYz9we2WAuL6Xb+oHumI5oDR
9aALAEAQOPJRMdvKeL6HQ+HX27D6naQcFnJOjzuDcdOPZYi/vgv+dq1lbjvqNcffJChnylbE7q30
+VIy4jfeS3LYwBd1IuJgJGQKKuV+uLXQuScx4apLSLNvD+/hKso8R7ucVyptyNHwemZd8dZUEcfD
aIh0SDOTOiR5o43B2unhrDZruUkB2qaATup5oexqtKMsgYvU/oG6xAcgyAed4mFS/DO4SSOwCk0y
dzQFCJ421PaE4pBe2PKEzYiD3+OlB1np40WqhhSIJkehsp8GDo1y2BuHdk5R2fUrRlFffM+A7avx
MDO2CMmBVz7zlbNNSwdMI5hi8isr8NK6YEnyGQExlwqOmrbWoHbpQDlsT23KOKlPE6Lum/VAcOKc
h9dSPKaC6wGZhPn0Fj7FZkJS3QdT/RRbUt0C5sjUb8Ki5mTF8JmOws8crk3vfY6Ybi9rJFaS+evJ
o6jRLVfkwYxZIW9yPfm+gtbkhAOT6WSGn7fhD3cyVEfCRK6tJDDWLV49CBkre/4JAmIqPzwU14Q8
j9Pa1K+3CM2wVvfBcafx3MNhdAlqdEZ4ky5pvrkCmbvZumrte2/me315tVYuBbL0xUq/URX+t+sD
NNRw8SqZkNdwZ0Hhtc14Iks769+RyYg1Ly5D99nEUG5iRBE4pRhNO+Y+QAL1JN/KqOTwmDRBz1JW
Ni09EifTcAT0t8N/D0ndPhXU/WNoyILCS0P973h6jtWa1t6kWizGKXIc8UzPa5lt7Ksn4jCZwdic
U4V97OZFsX/YP22MO7iZJSyWpjjTGUr9XXRZ1EpYUjVMLniV/IAVhyxA3nzN0Lzrzs8fsaxNJkDO
rQ2Rcaq2W9G3r3zHOLqwNdchIicoxPGJPiGm90lECJIGRDtv1BdOu/HrZDfIbBQiqoJbvDB17voE
YfFzTAweFdyRNvUSs7eP+NuJ+6owj0O1dBk28t4cGKa5hVEXqSFlugxwLhhoVefXZFMLR9LDBBgH
l5cf0UKwF6HIBSqX7LZoC9xsFMRO+tBcixJcxOVXFnsxyy6uAGN/vnbwOO5D8zSUqnHp7ztKx0Kr
QeJDjhutrTkFUlrwzZhKjBrv/Jcp3p7HqlflUFDsUGj2/JvL4bWVULRVNhe+ByBBDj1fgA5XMb4S
EwhuRS8Iz42hrcVV+xOh8YAyGFZMxxfbNRM40LZu8LhIV8PQGr6SOMrS3R253L6Ei0GMCypaL7hj
/gGRzpViYltVlwBwRO1+iNL9V0R3tfpXjbYQKWcRjvuDXcwQDZH4NoHXSQFUjTzX3A0LqJLilUhE
1qU/OtYG5+zdhKNUvI3FM77wi0pckMipsfWHtdiwqxCE7Scc67y+Ultl3axqGIYyelp7q3DsNbjU
ezQCIYpWGNwiUcNX/Xk+/1stDd8J+hyN07Z/OWZCCCujaFlk5UNbCAEt0VbazI5FiFIVWwN4XIMT
ssB15ZXOD4JLITTXAfTfpSxJvpr9mt1Jxm94LfJ5F7MFjbzgmISWYRXacuRAERn2/88b5CQbIuRR
ZNqvjrizWS3yPYLow3+d5XHLq8S3ZbJ+mXqgGVf97KQYXxD8BXRkkTym/bFhmz+KQgqDWqPq5cJh
d5uPDLGqRC//jaXozkYUwUcLLPb5uOQFRX61UxvH2V7qEdyUqbRHzX7FqXGa2g8pZYO83KEWfd4s
b1Ia1ydfYm8x7ByE1VrERrqO9pbKnzgtTDXnrecankfbiaCqWC+ulTn+S2o+UDNFAMl6OXEY8Gb2
m3qmvzJiXnUau3yjAvjZ88XbhLZXi/24H7sPVVa2/vwTtEQ9WINL6jkKlOJtq9MS4oiu6UMD/Rh8
kmDnT0fZcvntm8A35PsoFApPL1uln40G6kFVYyE0DXbYzNJNFeuJJoTI2QCD95G5OqCfKfZ3dRdf
QFzg1Eh0vPQwnPNeNtH40lql9coJGhSoVMvfG8NSNIkQuwvTho+9Wm5ZNjrlcgtcJRtktSguI/+0
zSfeaVEO0vA4vxySnF6nk7GRmyNq67eAf3u77+z++0GocC5LXCtfteRAKV158bTIIX7a+qrmNrkc
O4RmOKEJIzYJvxDbIHqhYp8e2Qqy/XLEpt6X8n4JyN6qHMLaveZrPvA0++wqlqS7rODPpXQxU0oG
0Enag05NyY5auqW1yqoUViq+QVJHWeVPt+SyQzsAp65981XksP5W6pu1MTW49E+0bDly1Bxtenmz
eREHYFH9C/rmfkvytnpoh66mEeiyOViU09VgQgwQCbfdAIC73XO3TA+hTfhZKhc1KcEh892SFLgt
oYGrdaCSthsI+a7RgXBFWqe1jw+WoaTA3jFR6jXGTKiYi4aYlKT/AhBonLuR27YAbLoBdqvz0vCd
kMf+gpP9/2RJOAT3NrnJ94Pobd7S7hPgy1OAyPyOFrLeu3/1k5hqCfWYtzB43L8ExE7Qy2ZztzNB
2KPnzc9JPZ7If+IExRBL1Xl6W/OS8ZiZDube9GA9+OI0OOGsFLNt+RShXQsfXjcR9oUdA7siW81q
yZrPF8AHSf7bFVADHPb3e+2LYv3kDulykRy4auesOugtknXIKKEdimrGfk/fms0GboULoXWElo6U
RZ5dsyatGNzHxPSqBNfn1Ws77WHCfBNxNc8fi/9oyBdkOzadvdVuKEJJwMmPsgGK0noew/I07I/9
sc2NFMxYd6ri1w8UAosdJuSf+rLGwywWmTWxUos1AceO/q9fIq5pJDAl7YedEOdFFqXQM8Odld55
6PbGJ3ZBSD/zjZgo/x0+ArY4jRR2NgFrptePwu5+FEXyyMDiwnmZyFNONSxl9V+73FMGIBZGMGCP
TNXuvgQmBEOXYoZLyQRxWMtNVkr+9WjDrYYWI5nyaMyTrmxpqdyqhIk8Ohdxqb1ucG9V+rbP1w98
iPM31P1vTSX9iabYcLlK7tUPcXHRyUOQD+uwomnak+W59U3LutHhNulf1W2VbYV9dpvcO4Y3G7Pi
ocwr+YUa/orJ/xCWMCt5c5dBRldvYE8iMH1rtPwnzwgUjH5p/ldPTg9i97XVCFdW1CJTj7byOEKd
YxHTp85B4tUWh9TEsUf5d+kigMimbLKa9XZ3H8k+P18Iahz+Np1Km7yWm6WZ1sBUEBxoaWRu529R
TCljpo6msf2S8Owmynmf/4o/INWTZBPd7tbLp+c+b5Dg4HBYlOShilOnsZ6VQsyLXej54cy3oWX/
cHn5hObjqQOOaYoPpiu/V3cw+hzZxrQsmNQ11dBOYXVlS6ZNr4KUoX+60Aa9Bf3rgSH3VjizMLQi
3MsN5SSq63y07NTwu2SXmJuj5hidEWHQiI5XtzHVLKdsYRxXBW7VgvHHTW6WtauImKk7pxpM/KEG
moaNzD/IJ2KWaz2ZFvy/mlCW7s+aOWyKgm4MFBivt+Zaoe4vnGSWFnwzjGsjMx0LXbkjyJgM7Kvm
mSffukMcSSxOooqZF9iF98a9rp+0hP9mBJwRrSzSugbE4cV/d8hZAuOO4Rkt9YGv/Zdjv8G+J+2H
7oSmX+A+ceq/Qw7WCHYq1BRBJLJkvk4bKVwPcKnNtoXDTFG5yRbdlhEQw/Vlqs+AR/6xcDsIjUW+
q861Qc+H1aK6HLvwtyhSGBkLMkKjeU53jHbbzx5XzKPk//Uoy8GLQEG4bN5A4lTpsmFBj422v3rk
+hRPFRqXVq9EQO2S25/h4YZyKr3lHLyBAU3ZDmYE+hygJcddva18MPd9oiwRyy9fu4eBnxTzQM53
Ov3HxJM3Cx7Kn9tM0ou9YUkk/A9OuscxA2Z+ltSj8VsTQU22RsROAScbWXriUXzdLJnI8JHfHDjR
pAf8M0RMH8vMsNGASHsJorl2mIaiPpjMEuGyZ5WR0CHlBizSbKaanzI/WD8cf2cMCCVOFbFla8Y4
QIpjsknjo7ZY6SdF/9wbeGrQCViNPPIwbO7YgROlpj92LpbjLd9jlBAY/dpiEWVER4/2yv5DOGUL
cAOAxetXLG95jvJpxLSacjMrVjxIwjT+TLtoq7uZHl4u6wkQJSlYa8rM6L1oDVHkE+HuyxU3txmE
JMG4yOJ4HravAsGI17iIhEROY+CKF+K2OhPz62BGXrkjxq/f2z6M+kATCIub1IQy7a96o/Sy9/TD
KL4IsEaDXjcFLpfigYRbQ4CRPne6WNlUCOfNCuuE682LrZf6nGyStczTtxlDVpk/spd7rF2fYdSP
j0DI8CLPPl1xsRNh4gqPZDPhFGWUG7lRYWm5dCc1KFM6BP35qhm75RjFa0YLvuMDRxA4sWmRNoET
sSz3Ce7+xWtGRuaBAdCwg8e5OcOx83aVbBVI2l98WFw1MQLylkrmxwRmzTdAfczWug3jhZCYEC+n
elFCSGsmw1eHuoRGOVSVRGrBdfB8ey5UFsgxjiFYQ96CiS6BP04mFBwvL5arxcwvq4m1ZY1Lm+6o
M7T6gg+lXvPZ1YVkPBHmXUtBuqOgSZejodfjqO8dhwcruH8HfwPthoJSRxpEoBFPfkQHYxIGFHHB
cW8edlBR/rIR96w7iOuxskDkMUWxODQJFujYE6lEOaTbrR6UqGpZPsKnbwncwRPVK1dcK+DA4L2O
F7r+u149TKLjZ+zqg+GYaKQGvqkuZCnppREIJ26BYAhg4IEfH5nC08MGkuFKEgWP8wDg4/ygAQeG
KUTx6GELagWGmz38xaW3qrcs6HveewqWQncGz00SZzrDuR3k4jpx5BHbXZc6nBBLqC5qHJ/lPodO
9AN39SHjQLv49ewTWfyxYj8NY4e5qVX8sWPioZEwq3NZuzZ34wc1LeNWxMgOrh3mwRBy75PDZ26h
wwoDAYC0jpnqxXTTL8NgQr7RXTmCEpJToHMt7huwY+yIH4Oblu//jY4po7BPSCINSStsnI4WTvyc
4zLuAVwlH3OFt8FJD5F2pg+/mt9hJZa1y1bPsfuI9E+M/tkTu6w0XlwfEgEnn/g/6HVvS/vBFPiX
3EQvlV25krL9rwOMdHYASx8MqZZdLwanT2kz+CI5je7dABKEWDBTk2GPaT1+rZJPygN4IMUu+K/C
GK595fayuK3JqMeUOn2GB2aamMyqyoZ+e8gdIU2Nqp1zMbQIwiREwHdUuS/1rk0LYNwO4Uih6J/z
W6QWxnzlOINYjTAUKvd7xS30TuLKlG3LqQzoiVFXmdaPd51qbquxx1K2mE++0MUGIbnsBypsMzZ0
mLugL/hCti55WyxHH7P2EIP7kyOeXsSmb9nV7lP9TIVc937/2CwOe6LZaRj1o1+jF6XcBWWpCosP
0z+SG3GkT+yFlzkU03rxb4HjzpuU8vOu9Rekr4JFNIQrZHoE8MOnISZ5hLW6wBi31v1wWQWWh5SM
OgHPkUvM+brTH3orL1gE/7RngDYZLhtw26qEDDBN5kTkMqkyYGoXKvO1Q/9V1P09vyx0dPiDHyfp
KJyjLYvW1b/Zwlnt/sRkKan2ZvaYQ6K9Sqmu6JDNEReUwwlWiu/SHqPLx9Yqu/rUr4m3V1pRLPVp
8O8QOKUxiIkNDt6PdPx6GViM0UBX9SRNaxAKggONv++9i+mKTj8NJap5AqlKu7NM/HvnMBOmy9bv
xzlrxztrlboeLWvWY5Aks0AnPrwK1n7SDuxb3JnoB9TMDklTau6KxFT2hcdkVpJJ1C2Hb2Rg52Yr
UrIOU87ifaNd4JY4B8y0rReRbhslvlqTw26wAkBCANO7Hjx+MAdZIphjHtZ1e6zZYhGag+GQUU/V
yPQORde9DWjIAc2uK1UfpCg5j5Gs2s95GnnYTAMo0p/1J3+p/PyF5luBsytdJMw9ThWc7zgXT18U
vKe6Fr54BsC0qwquPlQ5aWPRr+zgNg+TW8bFj9DUceFtDlupERPY3YpjK6MgBe4ZXxt6C4ftVbKD
Zb5l0EuMHlH8Dppa+PIPTKLJuiOtHVdygYbxYZj07hoLjz4LrcK7+5y0/AfAxxaYvo1poDfKJU+U
WLe49CPGYd0GojYllLiUU8O6mFN8H3gplkKtsyC6beBzAlejQyeyOhB3PfFwpxmz92Oh2PYiBL3I
1pAXLTWpZZRT3FlV3EhzYmiJLrjln0xp5/bFPpQRctNNErSb6UxH+n5Qk1vQRR7++Rik4/+5bjZG
Z/SzkGp/w9/sOa3rCmW4DtZA++ZyszliLOndkKzl8lkx1YtqzYb/YAzsWDgDySYNl/l0luF7jxmF
bpnyJZGLECtzQFYK9f/EjnS8nggAIPyAExtScfd4uMHCgzMJFgf6obVyPh1+ToPsGwP4SM6sCl0U
pWFHKRSHqeNOqWpczqVTDsMJZ4K9IUqOzhdutVoYSGuIRZ4OgHquvJVBsxP11NjR7V/UTgWLJnfm
utrEJTuyUiYNtFO5wsiY0YA21oEsSaQq+hzmuPsUIT1fKzlXEovBf5e+JiW5PAlfMz+UrfyfNVMW
zZNbEXSnZp2bS6ayz/rpsM64EnyZvgRSrpfITG2GSpP87svNW2L4TbSAEf7ug0/m2+cee0SzZwIB
2FtsqSb59xLZMyTvIQOSaCqpgJ0U7alrLWcm8t/AdR7r/6BaDaXXhh0iuJhijEyz0rZaKV5T3la8
iR2fQJ7uDrZsW5c5bE7owbrCoQxzJjwtoIePiLl/fLuAt1QbRqDV2lIdSs9mZmRBC7oi5L5t4kl/
InkTRR6YxsxqFAgQdokKYmeasHLWRK/3ofcmTaPDLpDMxqu0HWzVkLxzdvRpdXnBvTA0i7XApfzT
WD1jMZxb8QqELad2kx2eoLkx+f8d5WXShSrYIPklacC+Vq7zbiPrnTY1Dw6d53GnGjrespCY3vyx
RSkc4GuE/0YFStBEfjZxrh08kCET21+tyMJfc+rY/AkTonL8IZw5/Cd1yQghh1LwphrbT6BMCNTK
gOVrXk9uAlYEPYVxLHXJiYvR8LBJ3Zx1l9UDmdjzJSXdm3vmOn9TkLy2FhBeiyZJfx2sguWQ3B0x
3T7rdNsiw+cbnf7atEp/mmrpptexyzDYZ65MXuyxhvdPR2aQXLjRv2GKykxJ1PwHODpz5UztvIip
MBHZw/e36/YfhAcO159+Vw3fgy1JWBGt8JnV6Fqu08mjAvHYnMKbm9NIPE1+RF+ElGOFOc6oNX7c
13y74ZNZmVc37FC1bzga0C+UI96spunPr5XBOyXWifktCrg8hR/9jWmtRsO8aw7SBoStelga5nku
lyqlDDKWe154hcBtSDS7sWvJAJx6kkgqC70knAhScWOuUCo4uzzKwUkBIeuFaVaddmTSFRWLgFF6
+G3Aut4pUbPPLfvOlPKNMlvlWTgM+fC5MADWlF8qS1YD5//BZIqWcSD/+ywmS7gbzjgGLsmmgA96
RD7hPlXeoKwuHGOlF3153TBPhE8UVSSMulrrEPqvfkdVN+G6fN6CSX90lg7UyXyVyewgBi2OjmTs
1+NVXqGoy/a3Xh3wMnBHg6amAYrDe7OruomzInRZOTARn9Aa+8pm2bNy6omazkqV8D5KNv5zP+QE
mgftMpfBPoD2ysgAUeMpmNMS3CY513rymq561h5eiII0GteW57iABM6jWqO7T9EiM3ZBhWY/GU2f
ezQ35fhZVtC8IJY6r6eUhFREqkp2acRxCsIwyicjfITIO5dUJuVKo4uXfjONIWe5ZySICuxlXmI/
cOiXczUTK51tz8O+SXYZu4+WvzQI4gRtOq1VHLqYWS8vxSAKPCxcxaLhy9X69ZJ/I+iCfvnuvDpQ
M5IpXmq0HQLWAWvoQ+B1MAQWAHOSJy8PjbQHmVEJ+RVFVFq2Rfn85KcG603YgCosU3okIM/bh8c7
wUBnljlRyaV+h3UD2G4+fzxd/XYxjW0UP3H38Ch/SFLNSOIgeZpNYqj/5qfIlZdoTwN8zw3Ajwf/
iMdtREeqvNV4jD3n35fGqthY5F9uhaAWUhDMKcKaSUHIz3EiQPZS/cGGVyOxPqW2hCDPXiE6lQ38
BojL7eLE9GMhvVR/ETu5L+1ZBQ+hlKZOksKd5jt6HG6GnNWzf5le1vy8Y96yzrM5Gi4QNkacBaG6
QqCUyyKXe9+cZOP05VKn2EKLUGIplrIEDUqLsi+uEeNcwygRMOSH3LG6nX75MOyjk179mwlrJCdN
gkbHWVKSJW/I23caZiMpUmOUcAiXQ10CR8RuGxzvLwqGhiXxSrCYJQiNQYod6BSvwd+TXUcBrxGd
Ul91CJMyRh/7P58i3bRnGVMnCNJEAg/8XyR8Skr7UZRidLYhP8h/lXnbi6Wbp26JPhbE8jg3tVlF
nTSH9TMADJGQuWyccz721vRgNjspj7YAs83CN0s7uBaXT3prZj2auHZfl6D5o5tFRjpZUZGsWP61
X4iRuDUX+vU5RRCrWfk1vi201XpMb8xkf0baksshtcsCHgmZuxx0jAU/ZURWjseFLAU67m1CoUhc
CiMEZjU3sjbgdo/YeEqBK8iDLcuzYp5w4hj+GQnyx0DNwqYeDuuLRQvbeiuaCfgqeUz/TgFdJKwx
WbCokCu0EMuYuZxsOKN3qoqjg3WBu3citusfjNOXEOuu3okysokoeFCIa9/OmhmHjoxwtKxlHkkN
ZWTbRfygXnMCMUXLNF2rKTw1I78rUniMxKrY8QB80uRfd7+kS6pLSjMxb5hCDZ/stPpIHAA3YSwA
aVDHrSnwEDmK2SD4f9zM0SJOpLv6NumB0SlOfnYKpJ8JjyoLHdmG4IVqhzQcAdgOXWe5eQnC2jAi
8PeSHu6HoLRBXjPBXNFriEAerQ/tGmqNZsqUPG3RjPWp3FaYgm9UlfLE3YCumq0+TNCoX3SukaUS
xVVbasJXCKBN4iATUf5M0jrKoVdMHM9ZTItySzlLQeHLxCd+ZO/uEDpaF5/Q4Oh3V4z/EhdbsdBG
BUWrPDpRiXt7M2k24mYk6J74hGYceTKsq5YKp3DU4AVmb4SKTyK3Q1tHWH8vW9amehjkYzAAEM9R
/7JiYAehk06nWQy2rafqozOWT1dA/jOi1iX1tZiExGD4QJmpnFE4gYkw37NWf24E7BbIlUFKeyIG
DuO+sV+l548PJunWf9j9yqxj+loC1BufLtvN9Y2yRLjg2XTlyhxY22pG7lulwTrDmFq4/Lti4/Hw
8DQsnD3MNngpXDheo+aXdW7xqS9pDsgMlSW27ZCLMsaqrTgBnY3FEJqHH7Akt93UXz/qSMxjpfPQ
bQtZ447OQEfbyRDoPw9CK1IQo+C3tJ0bwQ/YMjzFhrTlO5Ug1VI1iX+a/CccXOPkMEEWZSSFAe9D
B4deDRnDE2qNshQog9znPzIrJyyPqTrFMHQdyR3ZUwrd2OGAoPQ/QBOifFHrOFfsY/FXwE/dHbXW
fRHTMIm5iY/Uvcx1+URPBwjld6RUTpu1N1CS3JCeBQUeSTjj7np0Jcurx1iVXvJK2aNcyo8jg+hM
anjP9oCvpaSEhOwnzz6RRS31tcfRa0d58qoknuHlRRNWIMd2Ef/4pH2DxXU4YeTpTFzr1ts2nZpV
X84O/DcpmumxkSDXu/3LXlKu5E1/U4uZdY+dmhLS2GY6XaFCk9mK4hOCuWjbSlnqn1gUGxdeDaeU
MsUMaRBgQJZeBMGiRf2PDegvBOF+dQwsj3ZPPYoRpIKhXYTXSijibjnQZysES0oVaSUXLfNNRblE
v9GMapBAuK73cepOu55RJg15+j9trltYz6l9pOVF0EUdaMa+PkvtclLXTsrZDm+5UaExibGnKwa7
XgAWd1tVQ0pcKVb8Eh2jjyAEO5EymyoJGFUVcgoeQutff8pO2Ohs4nFe5QPXmaY4wSl5rHXPNta7
pumXKDm02ngSwB8YmmHMjjM2eYS0FNKLVsoI0NciNeMg4go6E/MkhoybCF6TSi9UQvZ1fOzHOWRw
GRApusPTva+FBgQslP8TmShIPRORuUE80dj9YUfBER4sdafGAxO2o2ue2GIJr0Pj3FcoGcnzue+T
GoPK63Xw5/R+hwXuaiXmW/eixfy5tuTb5BhZj6aNm0BSYn+mw9bz0VUxI0g5ri5cOxtuHPidkgiJ
LM6NxJLffHNhlTHb0MOqAV/Bl7BrO68FM4q5Tf0XLdADea4kGZZh/2L0qBkFkO8whsBWnOM7JYaW
nBfTg97WD+qZy+iDUgBzXHziF/7M1h0mWquykf1PyI0Q7yZ2VFBIT9gYwWYX9rthvs+acq+bb/E/
Pm4GWTd/HExN/wIU3dHDKiGKEwTQRBL/gVH7qAonUGBosZV659D/N/2kTh4D6a4tqW63zndwpaQz
uYni+pdrgDg565sZDLyQricWgvqfpbBixG8xP2cO0BclexhZMVNvmtaSp4QZmDRNpejwwRA4PVo4
jIzQrVEskqszJjk63InLsPPVCjObvNQ6RvTGy5oyvxNOSO+1Txj7WExTFpJUTwqLmWiIbDQqbAx6
XUKBRq2lJBljX4l7tkDMI5Zaf20d/0poKX91/5B9Fh24EncSU5XoGUU9iWOAKe3KJ549xfceeP8k
gpwH5l2hzL90mgMhz+SEjs2PTuKpXxV/z0RUHdV6SmNcPw12c3xTeFAozAT1xyKziy6k/ZXvaqYV
XGqt7tR5+prDRTj1coG+xbfR+wJI5EopMhJ0Z+k+9tkzeNZPaGV2olXGxG0ko3NbXAm0t2B2NpZi
yaQOd+N6XMga7cLuxxZYjA2MUCuf4DayvJz5IoK5PU4Azv9jLUzJuTAGRWDp1iJ0XEva722XXp4m
dDAns2XNJAcJZUF8426k0+d/MqDY/ZPx2G7ZY2uF1a62eUKiaaezTUzNajn06St8qZWRfCD57HxP
AdpSJTr+jLOxaQhhBOLpEdWct5y2xRw8UAvc3ELsTpARmdPGWUcipe9ehTj9MS0r4FfBp2ZQwa4t
LZMDE6yL4zhDj4P9GN7tPhUUYod322q0v15lpwyP5IWoGEU7cNHxbS4zb3dYPLP+sIFFy+bB+llw
hCPvRdOoQjjRHWeXvF5fMfxNT9yfGLYXuFKyTKkqXrWehYnArc6gXZ1nq3BkT3zAh9w/ZFGqS+sF
tc9kbpBgO2M5DL9Ssd8BEYLtfmtBY7SuNqW9+Io9r1EcDVkW+sHQG02wPeZx39fKI3/Mbw6GfdXE
CQ2KiVtZ5pSW86fw9Z1PWO/DG5AD242rm8rKNM0kvG1IPrR4mZe/G3muEUfYN0BI9WKZDKbyq75A
o/PLkycU1nAYzwpNiqNkCGaoqv+tGOg4G6qqXHHaqjMUs2+318edlrZtjZm3bCPR84mx2mk231Bn
XyVWOzu3bUL+mKo1yk1H/h//QeJo3diQX5osbPaN6Ub30/v2F6eXP1oc9/jctDLw7MCcn/q8TMVf
4FL7/aMqCKqpqx63N267U4MNynvgBJ5u8AA0muCEWrRlfhJybx7gshjt5dW2+UQ90CDmw1q5ukPE
006/Kg2vlKA0UDDhktif6xwSI28Cn9boIP1qYFMRdfwAcjN4oYZP6DQbjQfEMQn6nsO94srL8dT1
77d+9QAOlYsdcTady2XV5pLTyOND+LYKAeou2EWiZl2saJH76ytNhcNb3iyNPwnskFAQ4Na9vcLa
UK9M08EdPG5jW77ZY5bzgRWCPXZYnEAM0BqFzXHmSvTkpXe56Ysh0maK5Vinyz8Gn1IkORR0T9+J
WY2HMAAe+2yx5xNJXqGXwIfZbvaMb6wnBVSEl2K5zapiwlZPdPKYxa1Y5ZTl7Pz2E8SHT27o/DGB
SpFzbhBsAQ/xQIys3QJOA1m+lB6q35jUDSCORlRBtdofEgr6DWwp29nfu/HhUxM7nOpOfM5oaBF5
1F2/yLzxFVtq2s+kxi8XFRLnmpyv7XeXkkfKW9uERx+TH2fCkycWP+M7CJwIiCRxiZoCX+aN0ccG
O6AfMj+ZvQHDnNTOZuCq8v2IZEp1KGWXVZtMTSW91zvY7kbaOu5O5HDj4n6YNxLra+LgjsodnRXW
mPuDazKQwzaIq8HHxhmLzfRkZJfIWVZeANfh0Lb31CNcunIBvs3/A9MbMBAVtT1FiQ5anOMHlAjE
Lcyn/133Ar4XuKS6P9P3+LsD2zIKgopeTR7veyjxoljekSpgLY+Nj8gT1HRakWaby3V3GnkGU3/i
BqV3wy8LWad08etq39p89WVlbH7oXI/owve8pHmTHMWcJIguf1ygsn4JGxhNSPU1Ldh4TN3Q7NXQ
HDzQ/Yg0BuSC4IQHCO6WkovqTP0d9lhEMXpD6Yn0v2AWkVNzuhpAK2N34R3/6tBaXvUT8txca7dc
DRgjW9OF5ooNYhq+kiNKsLBVNqGuplxm5fDVfYQ1HsBAnOZLBwkMIacFSmAyDb2zoQRBULU+LH1D
WIKRXcMc24yR6HpOm/EYaakrh12Hjm2ozkINAfbFJ9G3JYi9lLpp+w8NdpiBcpks0Qfi2xoj2uIg
t9uU5H4OEqWIwaoh4xDvgjUPjQF78hV6n6zoAeZfO5ihU01YtIQiBy8sjnm9Iz7rhl3kXn1e1JGz
QhlECzTI8wdqA3SGhhVDB05KVjiSPJfw2hXIVdERsvhQH4XLKggOjbIGGO/Q2mR0ZpSnUyvOTuG8
LHJAaxz8H4zabdI0yyYhnjv4e00P/BuAin1mVviCI1RfS1dRmVMr9f3fzsYGBly7/OofeeLlt9Uc
19CpP68m6dWKRZwXdCCaS/YqsTaBaABmdcukYvP9YAYi5C583BHP/ZLiYDEHz63KqH402nztUq3o
dyqR1nDwx/w4qVpomUaIfmIyCwbk6nGMzXUKY2VMxDHV5iJeHnQvynEIak702YGef+WwVHJwHzhE
+PJ8jkA3a52t9W2TXmMRV105wPqr241L8rVzoO+wvrctQSuQfdDEFCM76rE7ruELnwLEfCoXCFTL
GIuvsGe2Zs8Rz4JiPAB8mTFVjCG8WGVQLlkZZXOVRWwRfSe42CfA9fzIMuxEVJyfUBxhi4SPk7l5
arWtMt7NecJfFRy3WkOZ+6wp2isr9LnSfCDCjQ48F2XT2wg3w+vU4NG6eKX0+da+3i2o6iFO18jg
jTU0BXaCI57T2kgVJMfFNi1sF0M6IrGBejZU3DyrOEHlraT0zlpdsdKEBKgDeYpKUkA+oB6L19li
FFbOcZGWKzDMRDzht1DSluGQFf/e/d9klp+sP2/pZCT5mEvZ70a2diNikPpmNMtgBPViFNY9meWi
ZaLdY1+kVgwpLg19uaavIrQdEMy6qVfOY5H7azU61+xPb2dn3l8DbmravrHANR329R7Ep7a4gKWe
CUa5vuLpqLmrN95Dt9jVgR+RtXRaS1IdIZhaQvaO58tKhhVIfB936rYqcLvhycOsuWMzl/EJv+Sy
mrq9/tWxSfr4hY8v2wb6dpQYUUBOTx1AhcaAfXbxOrxChxdskKocOOxd5/JcA+nyhj31BFtTszuk
J9NkFUG2LN+ROOH0Z6RAJ5pGBb0jkz5vEcjG6SSw7qC9RTpl51CsVUEbL4SVkvvFKmtvMz2snBch
ws5eZDVLbKxcP3qGHAWw3GJy3rFsK9K79LjBZOh8DfMDum+GwFps+vQO/n2ilgwa8CQOhMOEYMre
C3Cb4aiMOEsNESQA73rpWRfiwbVtTiEZqh97zBkBnERdBQiQ2nUr41aGMnqC9pmC+eDxj4Q77Twx
4RyL4lsnE4SxBeC8QwLbdtB64stUAlerEWQXBrjNKwMsIihrUyg0QtkZguAGbJBk0rNWc/ode1Gt
k6nPUPEWpcb6+TCBjRMa0r938fkAnUP4wh/FppPxhWlbsBPpbyBkuYKzrpwkk5qPwZhUI8RyZM1d
Q9W2/q9J1/lDeSH/CLOyNhb6I9xtaoqao08J8tb2AffGbjpDpokjtjlVsELw1jIJGZZibbfOw2s3
4s69JKawPwcVtIWvXtbdt57yaQkNZNb1qcxZSBVj3z79y8NpRVqoBl7QFaSKnZ8OgbZVlQjhCesw
/QiLq3dopXfMoWOnMSjLksMjNGzJmKLhuKauskitSC2/D8WJ9ghe1ugfjOzNUzP7nA8tmT/iNRTn
JNWBwb9sZil8dTCo2kdfCe7d0XK6TFBTrT7r3IQXue8ShsqcH0I8RNq77ce1y8s8/mg2s/9xGHV6
dKGKP9fSoqSW2VbkbivAzZ5yISE543yB45IznRk993l5CVQEzWXGbAER1K7b3fLBuVF6irKQHtpq
a5FIiEgZnHOxoRBFUcavXKR+Onhkf6asiXMd4Obedh9E5Vzr/Gpx1Cj0eMPgi891aS8jiivwv9bq
O43Nhqm+UXBdnEPPoOdFrK0GRFYOaekPjfcPitqC3QtQg38woTCum4wcZBCk77TturWdujGvACm8
jcNckmpeN5q6iokW5JgehtbEoETPpppMbgJriS7158mk8Z+VelbBKbSmxKW7lBjdqUkKy9N9tZxw
/9UfnmMCLO1ziWq35CWNsD9tAjiZ6xaF4hAnB/eBGkLgweDPqBpa9A1AXaI3xCn7GsDMiqXvizKO
SnmUWDCDirn5u7Wq5+iETHmtZgdCbX5SPUsYHYpTu0p5ltk58bzSqAtr+bIa9sFzSUIZmqqNVN5M
HN91WXbpaFEhL81jO6Apb4aaLthwDVirVmC0mly7dRd1ReIlvkqQ7L22CH/SrjSu79VaMf6OEfid
ZBzl9I8gRA6LdmSGAQ9SdlG6L4vZ9VME6t+lcaUZjRxCPpidsJ33M58wUelr09VunGwGZdU652dJ
pxz/oZpQvH7n9z01HK0oUzejfHOvaKnYo4XSw8yZHxrRN6HOGGHS4xpCDHxRQMncMWvnE7pEWyTi
DcJ3ksjyDZMnUviGkTnHKqc5X63JRO9UbssND0KbPatB2aoK0ZcIr+t9+0RHQPqckH7by7eb6XoM
a9Q8qmGtcmmZnX3dkUixSwLutQga7bU8s8SOQhpii0hjIuNuLX21uX2dKj5u0+3vOk2XD3myFZha
tzNVhm8L1HVEguFYLttZWbWSxW2gfEbP1+Zz9rxjLOcGyQo+beNxK63NGKJFXAdNI+vrQ0cNxPCo
D5EWi1oLzyMYpuSqbwa8noTPACDCH8JFe+07lgcoyiMG2OaoFhFnH/ZjKQhsG9qpJdMEyNzSr4fp
KwfojcjnuCKAyqql+D9x4SkplS+6arNFWOc9m7KEkZH3BiNJPG05LE//QeioPmSIt9sV0Ob41Zt5
FulqNTjfWcJTfq6bxNCqyhOgHXUqdf/4jkqv7XceIQYT9gb/aTZROUr9eT+aQPTCmekVLbeJxWsx
5uq9BFMroiw7FSiMqyII5wf5oj0HtwvZu98WelNc6vWZcQj39h36/5kLchBxMpaXcZed+NA5Y7Dn
nhG/Vn0160srF4Xo1hztW5QrFazulBdMI8cWNAKN5EE69ILpuI33uYeREPfts5j+lnoeoVi4G7WN
ij/eV6ST8vIg8wzAaagm+v/1lQjAQsEjge5AHSwPQbgqqip3vGSUaB5pkL4Zm2GedWj0+/QrYoCf
WFf8/76oE5EDE2zpfKrTwlbSzKegjU8Kz/wg12GVDLevCu0/V/0HEF1HazZwhliSYFkBUALzQ/Dw
DvU7yjzvmys+ws5aORqcq/Y6r8n0D4/GYSxVYg25zShGSzO1pMW9/zhCeQZit7VSZI+CsTEX9ehh
bi5SB8fpLB/vF8Yd22TcsDC25tuMo7EDytk/5bLD8fYedM8RQkyUYbtrdUTHKRRubbqIfVENwQjY
mJHaacL/d9vdGn0vXLlSHkb8JjozkcI8RY0KYC55Co4mIHe7itK6tTbrOAt4Ie/jbA7xX9RnHk1j
BjWhCYE2D2Wk2t+6ovp2TIU+ZEyVqwomwXnsDND9YMuCbYTdVzxBc8szI0LxzXTS8KVNY3aHGgC+
s/kSyx1WFNaApZ0ubQ0KKczVuvSjufsgQvg5Bkb/Ra7JXnPpnfnT/DRM6hNGc/TkNSa8QTo6WGP8
MMCrCFVaZBX+s12CuRIS3gQcFxCqgo+mTVVqsSxQ73yq96s06adBjiDL+nre0HssHmWMNd9TcLfi
YNtrPL1UKijf6PhMofW6C1VMjmcvOPYrCB32F33oJris1E05xS9GJYUE+xbyo8/ccYr/fBN3WYzt
wHVT2IywxDnEcrimiiwABykdUmoqGQpKJc7Vl/kOXtFrZQD4pEBBDWxkksgoGurvolR0yZ9PtJM+
fdOa8uzwNx+O0dBv0rN6ANqDtL6zsAlliy15mtZG+9z+ciQWJX47WEyKgI4L7n4cZswUz7dn8FmY
cNmrWyWGjF+t3Ri+pbXUNrIM99GBXHGh6HL1Oy4y5rECdRHUmht9budI/rnL3HouqmYkfqJPHebB
p8PKT+bMwIk7jfuxDw/KG5DdHMAM4UwO4Wd7l8nYLghY0ic/ixIGWbPysPxB84aERgBBBrLz6I/d
Ba+wjrQkJbz2vLcJlOhA9pGzzx4yjlFXWBNcN8LVIbJAl6xUJDq3asbjYzagCzhbgiEk7d5gjLxN
k8HC4OpavD9QTWxdeX05XJDEynNXqGevatNktiLecPXuceR5NMZ0Td69H2bzK8+SJUrk5pyvEFLY
STYPYj7nEIu2+JgWhzQBywHGGUsT3/5QyYFvRuhGKsoIpcvVDZCskSAK0PRqdgVoqPAXIdzwMUos
r02gr3lvhoWXkNoYT8mA1OXPXohaphzB2F/DePuOEj2DP1LNFCzC1EStgct0BXq/Pe8x9YpIAOw0
6tuJRvEPNI52EY64GVFGf/X90jGjAjbUFvsFFqdMfvGNK1Az4eibAgYxs4UzPKTkwDD4MkYQpJ/O
3N5DOR82Ilv4AJN12iMPbAE32QvqJCrYLkuG3R+vrfzMZLoA7FQONh9YkEQ+DFuvRssh+eyhNGf5
dBPjAXswsS3xmtV0rLCnWdqMVfkuXQ/oEhyReQyYDUFEMeZeg8yhCpC3T79zt0PewpNbXecmqfpM
rQ1Xs7WkOlGzJ7jvyuGDU1USLCQreRWwlij11/DrRkOLuNajFJONA17/y5edT9JpwfGGk+bADcyv
SCQ74ejZHwfnUjUiitz/0ZqrWXRDfVad9IthEBwemPZ5RifBYCE9U1ZAdVF0zbl64gRxT9XFIgKi
4+xI9oIoAa+CP/wJ/tyoTMPvdUviigMvw5eWKuU5Kim4JRmQeTYuJ5UeEhHZaAlQBRTOL33kPR+4
r0PnEnYanAeXPtcOEx1E/VBI5r4HiQSzTX1cWFbYv19Sum78uHIesXZ3S0c+RBh8wo5H/HU2SJY1
yR7XvrvKUPNjxBHgsIiO2MFloV4rxX21iBFlSKyW77gChxYjry05N0LLh7iMzXhnRAjoV6kxZGoQ
n/zXQLtuUEKKPBsBoh7sDBrITZEvLnhUoEO/tpmkagkI8zEqHb4perKm14c7BBmPUihVqVvqrm1K
IMT/ujJthRpP0MirXvguQoEtvkjwESIci6WRcykahQZLstkdLF0sgx5uT+xO1tK5y+nOYaByigwJ
HKk3x9J0ie61nH5uaBFjcIRCc6w7Atv9BhqoVayYV85yGwAnYsFqwCY2neYGQDPi/40wfVcpJpuo
FLpYdoEuVb6KEi4Q/rISlWueGqC/vsemPiWR1fguiuLF1RGqaeRSdFB+hYam8AbNzHNw16Q4/wk2
LAuO9oDbsl8Jrqdsuv3QvPmmaKG/d/3+KdnmfGwNu+RAUz0syCmJOzhhKvGzu+s5jf74ro9MKIvz
eKD5r/z+vtxrjeXYBFaYg9gZjpGSD0cMsVTVj5EXNXEzsvsF0ZhAIXY4R8zPdQausc/v3rB6ka7t
NoVdWOCUCVnY/D4yY2idX8kdV3wqTYU4t15slKlELmkH2+vr26gcdMytBUi2+Cx3Hk+82Ji929v9
VciHr2veMUd5QYpGYLCez2S7/8Aj91Xr2IUdHF0gkwyjtg6mj3eVjqt40Uh1h/xpradKQEFKMjJg
EdPRpxHIHOux+tRrSzhF/zC6lQoRad4UemU4gXs83IKw+9eGLerrmJSMbCjrasmoHV2XhbvxuboC
yLD4erCQzFd33jbBn/sJL/F3dd9Pebs6BKoq3MdrLhKxTCoDHJnENMq/qbS+30fX6ilFy4J1cgUe
pH9eC8ozSy9QCOxYG1mdk4ZTp6bbSAAYMIflOqL6xoI55jWOwpShNapeDtq/0oD5RYeraSC998HQ
jf9mxu+2nXYB8c2DvCm6Xfs+w9RpZj4YnvdS0+YRCmktgjD0XoYiqg0nvqimqKZJ8Oe4mPLm/R4x
RwT3duZLALhGgJ2FEYy+iqQzSv83QXIwV8YGLaeHkvRE4vhB1YGLh6XJM37laYeE8HZdM7aN9syk
3kRPNliNOAvmmsvzk1cJdPt3e0vZ6zqpZOI+gG+7zJNy3skW8B5wRwndxTAB1HroofI0tvT+muQK
Mm+wk0e/KkVYHYKJVpLlY1KS7lnykZqd1t4zfo8U4pLlh/37JP0dNVis5T/CQTvQZ9ZJnCH3hpBQ
opZIV884GJXdBzIZNKJXVZdziuPQJy1CnV+r75AVEgMxtaWykde1aHgGphuhxOIkKOJNDxLd/v6/
UThWgKluloiCbTGj2K+n56O396niIzNR/QW/PFk5DRknJ0Qz1b+IlY41n4mgy6xG56UkzshsSTlp
iRAj8cBUTgyb/YPVnBIwQB+FzeSuOzdSvuVgBNvPP6+8kSGDZ3rPO79bdxSrrQIX61IzJfHeP3HF
DZO+9u6zJHbsBjXaM6GHPZxu2ZmzyE+khTPLKztU8u9x3NntZlL8khGXTmA39RleR2ak4HDTX006
SgtPb4LO3vuh6FeRCA78ZGrt5Thp2QsQ6T0gtJ9cd9RkWGhflfOBdmeENysvSGNkv2a7DMH4fFeh
DG2ce57PKuEhFuK+Lb2UaYRVkHzQPLBJA627Ivj68W6xSG70ErHskECBZA71kp+xker174qlzOa1
93ZMVB+HbhxD9JdyuBJwzhVQ94bFg2WcPhSehpSv5oYCRqUgNuAE4NEzVG1DLQKtm1fozDL1tOT6
T//7sAHXABoimp2AuXAPXfGS++5fSK/6MXFTM6UjyBCJcnxzpQ4qvsHMMrKNOGwX50WY9KmpeNk6
qjTp0TDC57m0VKH+FEZQYUIyJW9TS8gCLgAKRvS1BZFgR7mze2cRoPrpM8XlYeLIbo+w3lDdfQlr
HNjMVyxwVUrIfNUn6QT0hFuQeXoH3ekQihM/Yo5AfTEb7vVz59A8j4Q5x4oDPC76amlfAIYl1F3G
SZw/w3TMKL1zYTfEfwFmzIj9zSkWq6ceYsouSVKMUROY+bFwebZVR+MRwDpdsfpNOj3kB4TK3m8v
BYkCIWg4Egt6PmmJqzrVZ0hjTjLq/nM4LnJa4uIu9YvLuDnIltsp3fD69tute6gloN6MovGoIZ1s
iaMbtiWi1/loa89gQ1G1EbAs3VRFfEHO+I/TXw/FxmvRKjX9QQEH+TdrlLatkJSWKO8aZflX9uMv
KntWdW/y5ivy4wNArj8J1w7BCakn2Ee0UqKm9oZXTV/737ebzrMyGYXqL3ak9213Qk1bW1Mzjink
/uTC7qC1Vgiqm5jRYopV4VWbXgk9NnJ69MnglY/WhH5mEI6WZQvtugfb3RleIBm4wSX3aUI8qgmk
Vm0aoW6M+tkMAl2jOAP4ND7tgoDXFoMQYluPfQXRS8G6qHZUGBjnYcRodY9wgqYFM9UP4BYUCQ1G
8HnghRyUHJ2zpQ19EIeEzOM7uqH/aRu4ryniuRpHOLr7TbMJnMA2QzA9la7n611tCkiJqg/M3gj0
TXdVs66K+MSFgiJ0gU2EFxmOmCkykH/+yJ0NXHQ2ovDslQF702XksEORvNf4/PUe6Goe6ksrSBfI
knV7n8lHDXmzWS7hn2G/5vmcmjeUXZwCZfZCKyHbTzg7QRR4sruEIa4aIHDldpTqZs6I0+Tx79/r
JTNEros6I2Um5LJ3XVm7VcTSdHX9XIbwjtR5wiZIttUQqf+ESMMwKf6id9DFpANaHrMcxv9GKkhJ
PJ3QVeBjBFszg+TfR8OVw7ZassvoQvPLDuhriNQ7fcebulZOGcb8ijFX0LeELwz39ti//TWL4rau
r5rb5L3IMxgXcuOVuHKiRZ7e1c1+YoD9PCMDOREJK3ZF+O8MDbyM8zb0GifE+6pqu93cqvpvaT6z
UgqSf89kPizUdRH6N+275+uvi3OgTDzOkf2qqeVt/twwqrO41B5KnH2Y5YeENM+Fkdi4ZQslJnFM
PdnAf2fKjJRNed4hlDIyiSnvgEWZJxKRkfymJbvq0QB1DPFxIvOzuA6dWiLoXCwZMGLYLoSUxCvk
Q5cmWyMO6U5bh4lR1PPVQFlTP1vlgKzX6/lsY8X3gmGiCSD5XKDkkMThduVcGYHwr9In0y9a/0PP
ZVDZe6TWb24kgnYlr08fqwsjB7Pv7eiuVxErCsyAf7XLatdzyMExF2YSZTAz5D3xnw9Q4ijHnS4Z
rrPZ85X4j9Ls3vEDiA2Jm4rm6lZ0+wCPrdqABIM+qrEhD0FMEM+Tn4Q1GYIo8VqipW3qsWKhBpyZ
T1E8efsRRxCGC0QcdArloffuMOV7b1aEoG65XdYNDBVcTO9wKI+dgkqQjRcRRqk4qC9IImLGTVGu
AItzLHoVse4k9Zd/5rs73fJgVBQNZtTF6szqNkreB49ChxIGgfU31Ko20HjZj4ItruoZ2ygMcUR3
kr5iGSTVdoQg6rwj6h+UbhFfJDrXitqzQLkt29ZtdA/7OjO4eeWaz+/N92GJol0/M7ReSNLkf0H6
RY0sSFVl8vqaZNyUWGGr4Cv8RtWZaRIh7rKTdJTfa2lWoTGa9xnODmjdyukYpiuMF/QlH+XPp+1n
65cLz6S/lhrkjYF9YS4HF+hFzUSjSQnXGlmnLQu1yqRVp+DbTB4Eqpw44WrEh4gs2yvfw04lfNOZ
WeFRLN7m/1OHtOI1FXl3AjfAs1eBcSM6SM83BcMEmyHnqHOzpgGA9au0wChDhTIuLktrJWB5niKO
0RKmPe962WaBLBZz/Be8Y0YLFy2Xl8ndSMhQOGkCOmKIcVcwpFDGTyCMKDcPbNdK+UlVQOiOfu5a
wEccyb9vXxvFFyEnt2afkriRv+rVeSLCckmdK9OT9jbZzoWDVp0ospWq9WxIEt1ZCAmtvAZgmjPB
9mf+q1uX/qoyyASCwY15Zgah0k1UISwzkC0mlqxt3RYsyiqG/GVsS1aeszDSL/ICylNOc3uzz1Jg
9BYLwReiKRc/SEVm0J2zpjxQtOslusgoLwjHZswDFgi/VsSCXTygQMNh6P3H8uPZvCB91AiHHoEW
2Ap5Qvzbva6S4FCIQ+aOkDbngF9CSrLzBV7TLQIg+4falnOQmBpwr4fzeUoOlQ4bpQzn8YLQbR5N
Z05CT1tOP8KAF8nAIFbykMoGh5uWbF9Bf9vAFwB5g3x4iDrL11nZfapolZK2SxjzCdoudLJfsg21
wrX0HKZxy1jo7kWY8anhuK9rUF4YiUH5Cpj+/hzAhZrTKIQwFb4hyvDX3lpo33Uu1yU5J58b0jA0
AG1lxXX5l06KLXo3Vhy+6evjTtIuJv07QXgHFwWqDl4Zef+7clLTJXRHAD0ZfhQpQwYojoBvCEgv
KF6N950TYbn2zZ/87qrGlpFjVq4hME18UmJYb0nlg5THhKUo4ag0vtBfQa4WYbYS4KMPYGVCFGS/
vSrzMTjdfNREyB20EgQcJ4gO8L+zdKsGmvTh+OKFGTKcxCzVMN2IFdILYc6fu6inLSvQFg26GIxw
XrKSPRe/j+ipQAqvWiEQLSokymwDRl1RUTokcpjU9ekrJnmGsISYxQ71bHq2z8WaU0589eurlAdT
dvAKooReR7FzglaiJVB/0micwwXeDWxY9yqcRwuYuE7MuoazhKvloBW/JCsv/NcNcPUYs3mlMCDD
FxYnA+GzPQfP1/6pipgZREIqem1kdV7MVIA5zeSFGrXd+fBvwY922jH3DOTQvxAoeLEAG4asz6ff
7ONJh2CJyChJSiBRB0tTvgpfaVCSPgNaHprJlbtoNkA1O9spLTZ7WxSs6zpVwz4OxUhFolPff/pO
jfzoDpAEqFxmjkpvk1voYw7K2iKTvESOefheLp53Sx4N7VVQ5CbAiL/D/Awhd4yBJKO+Z7pu2jw4
NyvtQTvEcbz4EZ5AYN+itX4bCjJLrlgyfuenAyygl4lHD2P8ifQDpU2qnN0ihrN7sjtx4MzwJ63V
+qHHdwc9gsrGp0sLBXMgXdwXOAOmbo/t2xoecY3bcbk4zVAxrsie/m/CuERLwQ99VgB8nXQQ8N70
8ZX5W2+BdttRtKN9R2WaUX+5hjcHv6l2fItrvkz9SseusvOxDJz+H5ybsVoGUc8q+6p5dJG0Gc5A
PLDRZHTMkT0M6Bmf9WpnJs6ja83ifA1v1t1kQtmwF3vjk5ZQZLLwX9ppWcy8h4VVnJ3pCM9zFtIb
tA3vclZhlYDKSk3N/erzP4aS7tOaYLVkI06EpaFzNoA1qy9+fv+dioqXZpHfUXYv+GXDB7Qp9uZL
B289H15d6nTEoD24IpFX0N3d/0Y8mQ0FcVlN5xSxqwsuiWA+QKaHd+6CHOv7DKLLxoOVk43x8yc+
VVm2zpm8z/Ix1GvEY9P/dcggyMbBrZSoStXLODAqXkG7ZZQ/1qtPLwmzeKlreCOz/n2Y7ZjHFETA
smDuqZKRVvCVRZOIkKLP9mVnclBXNUrkU8VQdYxhdI0sQYqa02XMO9BguOyW72RtJTWD+Cylplp3
ERKCOdZgsP9sczl4yUs9DIu8bRdNLfBO9VwPFxRJ+qWoddjSraxMMBZJdFxFahQOYyr1Vk3OHAIl
HEQUdVgixw8jTj6vEdW6oa0CaO1mMbEl4YiNPFW+pqDXEWba9NQ2v0nmomFieLRKfb+hYFjo4htK
EpHrU549dc3rxeZVlt6pEl/ViiO8Wpc+cfiLjO4BgbT8yJJTEPuV2WAOBkXCNLzrpMx0xhiLgTS1
GlAAAv0hy5poH0AGtugRcgu+NcUdsRV/Eplw5x/kc6HUMTEvy9dzM5WoIwDFA+EVZChpDwtpxnKc
QOXx79GeS627BUOgp6zeqReYuxpO4G4jfgJTKJBeGW3m0Kd5MiJYVz2eTpxICF6XmNXcNfdjGxZZ
pLS2XTcHXBI4UZXDJE0OThFgjSiX44OEIuZYJ0l9Wd1hy9yB7ZioWtP6U/bGMQwQX7Wrspj5apMB
+GbBIQA4Wet3TSV3oKS98FvmBcBYCdpNTaDJbIWqjTBh46Yb2yG3+IdEk2JQL3fCLa2840RQSIH5
kV59L3cexqRx08s3ZXP9FaUmKOeIo5OWPsuFZX9FsVRfSO+/XKkM+DQxO2kqrjIGoT/Mn/AXbdYl
eKw4K8sOJKYYhQe1mTnWdtkR0qtAgdaUKFnCblJSVImecG+xKdL7w/7wBC6ww8mYjIM6CXDvLlmq
qF9mMjVyWI9bPLLPD6MD0QB6Rr0FTwyntBEAxJ7gaNP8YpPlSx2B4bCyCmF/0Z+myjfVMmeWXRDH
dEOwvOeTn75KwVU7GpDmE52UvcJZoRIeZNqETIeH4IXRKZ7fecjpZTL5255ns8COHaIYiQqkYYbO
y5jL2b+Fwsh4uv+hxV/iHzGddFbp7HVmiYSS6nXLV0zwdq6RS5CMXEUDZDKAGL5OuGeYUWmhlG4N
V5Wamo/gp2R76QMh/DeShNsDydcbrl9eQSIevt/y+fjpYDYDBChCpKhueGuSJCu5sYjQBekjjZzN
mBdxj+Z9/zMOeiWQ5loRsixpGqmKQJu6jV2XQaQ8UaEDFCZFI5iYT2ozXlX4pAqL33bLUKz5W4AZ
hwydmYcNZb/joOgiIhKtvXY5UJBgYUvrgQ3nXkqRr8vIARniUd8XMhrZWX6b6zMVNP5I/TPYzhif
43Jwk3ECLqDTdaB+I8iFxe5YiYWHolOVk8k9cPUwtf7NoOJfGkI7+N3X/I/fVdwfqsf4xItes81a
mpxEl1d9xWkv4WcVUNsqwba77qXo4fdjAyB/pU3uZD617ErAe2vz545ybNDXQgYBLJdMLGzEnPqS
P7SyienDeH6CFCz6ImnLxj8lbejbdOT7m02WZffTyj8DFSYeGieIr22gelAbX1BCBqHqiYnQ5btY
LCkB5N77hJtJWfXNFu2raooWZFR+0zNuZEsdQxrIhxiAexwZMcP4Z46o1DnJHNGJOlEkELPq6G/R
2dFR6iwpJRiOk/SElWn8E4K19ZwtVP03ZTXFGPvS5L/ZVIf0ArsNECtsCXMm+f4ZpBGw9yKxrRQy
V0DOkmQMCBvLLz4+Q3N8zJp7qL+rcilq4pEr38fIafmzKtjY/LSPZZwEz+JUqAbgizpYn2p5GUeZ
IguUEMYp8+6YZeOcCd/1YPPx5ePyt33vJgVYtKFOgSrBKomJ7bP61lwTyKRbGY/41Iz0SYAXTguQ
b/phMbemtTkQbFJ/EYTysLg7jvrTMsIOGphkp3G/hmEKU0Ft3bVP3zEZ+0cpWphqO7fn4izTQ9lO
ViNH/tpvic6Bh8f8g1dkAn5ld9mwA/fn5TPxwNP4imoLoggb5asV5J9NfCj1AQz50tF7GpO9F/4b
O/iOgzb3Z2nMfCI8hFZsP11hwCX+I50GX3rwTJjAo3iQPnDZBsBLx/yr2n9UMlep3WyUGbViU8Fr
voWsux0x8BJSgfY0gyC0rCugr87wQvufAZCEB6WffMDzRlbG7eIJZwL4l4pPTLDCfBKoUqpvimHQ
qricmVW6aynVM4OQLLsqxSGv74tChbKjnhEALlHkQsqLRWbMBm839Gv5yq6gT0/e1XiYe7YLDFf8
b0KDnLi3P69M//md2POw7zXKYu68m/ENddbEQ1EuxIyY+2TUMZHiS30ps6dQdz96X3DHnuF/1HHW
Hqo9CiskDkznRkK9ZiIb0208zk1WzCjjFy2rDUijz5RHqUrFXykPuQUf2uJ/0p7VKREgQZKx9gFS
NCq8cC+1soga7yu3DDySm6NPnd27PFf8BklVhDby9yRedOdcB7c3IKrorLvOt1rC6GTonFmWw94C
rtoBKCNU0N5tNk1DJmDltVh0+bUYSAq53W23XuiqFftugDsdpt3R67ofVTlYSEczFMgmfchcC7Ft
fpsM2FZGcl3XTfdoFwwWDFm8I/DJJzfLCCyhTE/0qw3Nrqq56OqMcy8Fm2V+F4hC6l2O3IO8DU0A
lynw4nXYca3ewmfZ2v1FwMtZnbKuTKTeVXCRtGGKPR7D6329exUvJLCR6ARXL5zFwjj1P7+gbB7S
bFDyH14JLYJMf1/RGfVl8jGJBGqnn0U6prlL2c/T05rFBPvM4VONaMb2cLltXHwJdKBcZY6bvgyJ
EW2Cl640XiAicU+YkABvffuqzI8nl0dbx5MX/p+tj3ztr6kC7OZfrJNc7OxO2o1LH5lrExhr6kSW
sKEOUss/gKvHf80/mhya6qrDSL4WgLb7vKuEdWLptORbRlJlA451NTOlK+aZibYrfjJTTQ+QRJUC
t5ZdbGX93XbkjPuMwQiXrzLwW4x0ju/emFQf7A/rDLYNKvT1NRzzagYaOBNNYnNpLXqaAK64adMZ
CU175fwHokR1F9tHAI33wr96n3tviOyOsMbNfdBoNk5EO1PTQC0mReVY7VHZPM5dw5rPzCDjD8IN
cBFVUrsCOWG8MAK+s/5prc8gKVbQ+fN+gzD+HMWE39VXUcvRungUv52x05JxbVmk2duVcGgl/PpV
O2P6y70QgEn1/tR9gHidW1Shh1Cn0IXj2K9seCHCA1PH2bSX6USTlvOpmIVjHew7XhXZfsFlM+ns
Vkth0WoD932vegcwxVxrfMXuyy+ckdp8mbd6DaQcd7ioLGRKZD83RLIz/aDFsW4oZST/xquu4Aa9
Q5oPRVJdAEOVCiPE90JSNM0VeQ5UoucSMmx+wnsGbdnYCSOypO8KAjZZLbXbQg+jGc1BSJLaKLpf
miXF0LFfNrBdd9l4YolcHa6bjwsJuj2kcQ5Nl5Dxng4qw542jaegpy8CxLP0jP/FJyq6qR4Ybcw5
+vU6gUSjHdbLXw+MoSA0SgegIskCGOr9CqbGDhNE5fFeOpRYyLgWL+Y33r1Nm3oW2aipW5ukRgL7
8G6p/YVOW6HxIlsEeqnfQE2QET9wLa2q7QWulp+m3BUCRY+Co+sziWjHaLPKRexMdy5Ysvc89rsb
hgEpPu0KZIh7MAveQf7D4jk6q+PY3duAxCFojvB2iPdqY+xg0lnPmnvzby0z7aECj0tzqMGUL6rc
OpLr/VnyU8L1252RnP8ipk5lBr9VOka+EodF3ItFCrn6N97xbzAXLqT/IApXa2/af0tPJpe9bP5U
MOVNW3z0SG/2Rljj3tYIpS++kaRd2QWC2DnGlpT3mv0jtQVr59Wc2SKlMmEtZ1d2eLmHmjYCfZ4L
Z4YbIGioyiEs81c6Ju/jJVc8ZYQQiPeImCDW23XAKgGa1RXvyegZ8mGg02sFPUBRIHzMbUzIlhWa
R6qdRQjR0wpGbqov/EE8tglXp0yBQSREQio5YIPcMJD99NSrm09viYx5eRpYQysFs4IZkQ2vLgIL
sVcKQ+K6AQIUZaB9AX76cHd8cCyXFLyW0YR9Z3k7KC22lP8OLAbAjf8NIOCRExDuauMy2Qeji5hw
u47g2Nwqk2gi1rWkJMO9hbtinj7Y+a7twnlkKh79A2RVRGIlz4KoibmYdjQYOdCkrTEoKzXgroCd
f2H+KpmEYfkPzwC2oevGSmjk0EJluvkYe1K6j3UyLXs9zh3xerhcslEvuwefo3J92CKSa0ckWqUy
xP2RpLSZo1sRIh9r+iV96Pu3wrruLBYu7OYsL7C8539MHTuMPO7ZO1YT4stQm4K1UlTcgvXWnsUk
/cjIndpsINNooBhwfPTgbyZC+/Ggnz6dfMDw4WFhV8jyTvMCh4fnIq6ubQJie9+Av8qX+awJypxg
wemZ3koIdFCc4zLbJp7hUT9u6oYIGvfj6nMD65h5p/8aii7pSJbfWBL3W4z6lLzp9+UQYlCvwDJg
sNW9q7CHpgiEuxhTcqz+1v052vNb1EC0aizWlOds6Qik3kRE9hEnC7kJya/ITDmFpHpoLaGMlNQR
v6WBxUoljeqYrR/a9zmLyiJQ2DgJQtHheYyLevbSw6KvhH0sx/SQpqP5B8jwPQALHnrxA9Q+scxR
USPPuLciVYBTibrn+ptDLYbGfip41lG5fy2SCkcSVxXDbdvvBAskAmYfwU5PaZcryXJWdWFHU2wi
WCk7aOJgByHodLNg/ky+GjDNeJJpHe+MNKf/SYKFNaPZcqubTl+ivCoCdjj78QPcRvD101WnW785
alEkBbq/84x+qwxKmtB6BiRXxFqN5FnQmfD4c/FdtgX5C0sTx+qDD0wDp0yhVacUIGgHaLtDAzro
bbP+QNa6FeeAHu1E8yHQb+xTOFIGf1M6AleFRlYsEHPHWsHJdrW3RJtSWc5n8Yndc3YRBhC35Ect
pnxutL/e3UMIcKX3nYjWbqUZQrWJ7uptIk1i3TfW5SDieFhGo4fity8lzpr1ZrNKdiQ3PE2QZ+VE
UkOPX4joccQbbumNWoNWFTAmdY18mXAznXH9vWf2xKpuEu1X05YoMJ186c1j8oCs0YUp7g2XJzn9
QNhdPIsvDzsZiHJF/unfcJJmPHNyHfHVkXclKzkrilJTIsFLjNs0ljFUFncMYhBRCm6C+NeEa4Hn
e6I3uvz8OwmnK2Uo7ooLxIuAZwUprt9ukhIdHLpzdkZJooZCiWDOMckZrTmyuigQk2xiljTpR3Od
QqyuSA2ts1skpUaEwCJ2G6CnPzvEXFtzE1wsYySBeS0/rxGbqnFxBe+Go5iPHA9g3FlTyEcuY4Ik
5EuqofF1gxtdFINlPMiWU0UtidKv4J9SQcZ8Gi/iARb82alRPRWJYbM83HDXY6Yx9imsdGgP9SZ7
E5iZeu//eFynyXqTZPxgFCFNw6Wd4z8vPyXMKLKtpRnAPELRniu1esVvOG0CnQnqnC+vtq7FKCED
C1YEowVNFkHAclGbKvMVN34w+X44Ebk9zkDiezjMkLGuHgJE1cVyb/+503HaGbI0U0oAUjKUWTPx
2ZDrgAq4WkZD8AftUKAF51WG8dp9ylzD/wAHuuXiwpQ7dC3BSa68Pg3gVkvl3wIhzLp1sszytP/w
nsqJSkzm6DOrOSLyuK+1KyD2E36uxdiRKFZlgrXbFitqZHrJ2MnYMiWweFGFRHePvep+Heg7Tjp5
jvHRCHSGySyT2um8mksHoDUeyM3hu/8p2XkTCpsz7qi7N3hxpFUcgG4GgoG9CyU4WUAm3OHOzGNv
lNEmJjoFthRTKmxorGS0P/VyZD3+T5U4JMrWv7++u4fV+4PO4PY4lZrFCaF3AuhvEtO86wF33PBW
b42ZV8WUyMi+l3oRcyFdrpiSdlZTUDgKSTa+s3yrFC19JjrYbq+i8Pbxag3cfQLUCwCuDDPbIF23
WAMrjZxh8bWG32uE53QvVPN14xXrro38qr6eMWqOpk/jG0zVEkN0mJhGvm0ltdnelfXxHxyOlI8h
djT9Mmb536qbqPL9Iig0HIC1r2bNxaraLI/VdgH3wy723nNL0wAlaod+YfpcsJwf40qBTmPv4JCC
on8lqq+vbS12ctcmihbHTit+6Sz+WqTeVpF/XRlF8tQoF6oehznzI2UwEgBBuIctG/ZcEJWcm9zf
sxIDzwFKyFBG86HieW/jEsRCILpd2En0+CqrvKoxSvOmERa7z7HT40atj9/oJIsLQiclaKcuDFPT
OvbXqNktRJZMaIe7qyqcKCspRFDdzH3sYcFwLWTRniiSEUMfka5RUV8ss8UH2U44ngiFjKKNTsuG
dDNjkHpGv6G8EOZRb8FllhD1Evq72TOiUOvLIuHzUJf0bQfJLuHpvC2GswQjjg5lph3D5d3xOhj2
TmQdH+/OX80fE6JSLMlRwToaD635H7YvDeD2zatztCS9x8ODAjtcuQeYdZ5jesb3u41hA1r9ulrr
8vcvFIHU3xUQZFqZ/pbfDhAIVIw0JJrbhH6rAjEm7w4936a89BCRRAFjtqemSY3snmHplkkxpS5O
aa9plY09Rfnv2uZOovC1wnBS9tvY/P5BPNjkvcBdP+Z2cbigjyNGBD/cjr8/ycGT/MPtDZXkotWK
k39usjflE4kjdL8Bnl1Vep6/X1SaO79tF5Q2EULp3LU+nreI/YRc1M+lu0bY6yyoAwg6JkaU4mnj
/nNIaOX0UUu6lWc5kkxpv5E59q7DAIYlJKe0Lu+wQwX8FWIXVe/vWfikwd1e/c/spzMkzQouVa34
6teZvMEwMbJqwGjQbQVWgzSJ6tvl5IG9zR1yXUkUBTXtW6TOtpzC4Iz5zMHxyXOZlwOghleZ2bzO
gTNFpXOxe9YU7JngVEgzU86lH9tuh5D8ObfSt1EicFjgzrOId8Gri6G1Px9n2vYZaw+liqZO8DlB
YF+pau83bPPSwvvmU9zzhEOqt2sD9xZ2WEDI9aKWmtOwuo1aH6Ak/bECTzEalWAN+wqUfp0v+jEJ
GFNJ5bTkbyUTvcls+e+JYaeceob8sNKoUIrkgml49k9vP8RYPjk8daETy4unOyPuBr8IZBhuIS1/
7Yhxn8EIk1KgKcCR5pbjZUE1A/C0P0CLO6sCA1gLK5sPp8rqT05peHWgtIIF41/8/j7LVzuX/4pD
HbaNmJn8E2wdlckv5R0P/rqXTAlMDW2k9QBQwu73jgiew2ejReR7Oo2zhIL5HWNVpHxoNtq56L6z
193Ta/P5cBpp3z/BvxCYP5Urt06g3c2aHm0xrbLb7uhPn9jmWq4JEwrM7lOJl9dikdKntFXVYDpw
okppbXUFdyDc80j+2sTdNbCuxQe/VGQ4vdMWf583VazCQnsyssJESIMG5IFx2hPi1qXhHdiBFPZj
RrCC8ZX16mX0TGn9gRXt5NA/JMGHh/kPQimcdGcA4DCdwi18JLSe2nCKHEvHTleErN6s3jHOYvtX
zoNmGGBPHHnni2xsuz/Yj6iOAvvlQUQrE4HjYJipsh8QZ/vfRPubMWW/H7cPXx9+kBIfJLliiURb
D0AnvxAOSZO6OVc1KVrjy+bVWJd9U8RuczdYHRXiIbSi0t/wjvW4LDJUihrfSngH1xRIgT8gXlwC
5udLpq5JFbnkCILrm6jfCmhDcF36lxjd/ZqSu7GicLHljq7+HRh73obIqCFjaJ0REoCWI+NNHEFu
wqIm/Zs4CFoK0ObCoctyHFuOj07+5q0vEwnPUT3ZuMk5GFq/vWTHZEyJJEzlUGKte8X3y+5RRU+v
jEY25yGULpf9zHfc0kunn//ZGag8Rvf0HEbz/8nDvBlN7j3bA2QD6KRNHkPegoU3wTdYnC636S3J
8bS06SouWlTB6BMpjBkRr6bnubkrf0OP9eLQ+YthaSXUrq7ZIGwn7eyiM0602SvCXPRwiTGD3UxW
/j2EbDDOk8X0Ra1pY2yFDhsQhZ0svjAZFbC465NauAUC+VcwjWEzjQqmW8ME78yob7VJ4bXUbN5u
7dF6XsV83I5sRMdL3eMoKlampRNtHYTSX0jdTc5C8aGgX7rqyAJroDAPTD5KCW0IHd63ljdPZCnj
Bzc1Fa4E2NMyXayjqNyVTgw94mFcj8h0Fgi2LMFhkHL0j6VsLbKxLXapE+wpKNKl60dEm+Uw/EOl
hlqVfUammkdpKUIArxJAmbFEasSFAsGJGFizM5/ywLXArDk5+yVTdGgLHOiFXyiyN5CiIlmZS7r5
rMp5cmy6Fguk6NpNQPHDwqUh5TSWPFKvj1CitAHfGl9olABU+r5UV/ri/Oyeuzmsh2VPC7VM4zNj
JH0fcB6X2HJ2s7sw6kIB/iNYODD4qkjTdt/tELjsjL/5Zdnc7iOhuBfRg/1KOmqLkQH6G+38qe+c
BWAKC5PrE0ShyGKc1eWc6o9aHd3Ext0togQ7you3jC34fGdGRzD4RhNvS3jnvnnM01hE+9CUGG+o
YZJQQFI5chhgxD5hob9u3PdsmSV+kUoBThZfV/2lUsT7gWD4y6+7K0qzB7n4AjHN9XuJ70WVasmc
GhOznZYPWdD9Lk8g+96QmZ1z/BvGrBPNteFYFIhObnTdTNHVgMQOiGB4SGX8EaSVNGywrr58P0pF
GTup0DzPDAIYmO4NYOzUC9OdAtFqrKA5uGIssGrHaMN1DmIJvDcYtysT1XDHUgm5wmxl6p/mD/8f
A4BBicjfzomPbF24lWcfpcWfutdfrzwmEfC24VgwsPpWKD/g3OES5p96CrCWRq22tCo0u1L9iP8q
Lp/tcmj8tCKJFD6aWX+uWRuhvy/yWrgKWw8nbjL+e9GChS+oOUby+eZbg7ThdUZbz541y5kg4BaM
RSYNbFns/mBzQvQ96v4SBDafsNs2SS4q2qLn1ai2YdahLZafGiWNBeKmwm/Nh4A0A+MRJth4Nf/R
4pqdyCtWWHGiEZnhuonB289JST2+MBVV7qqg03mE3ymZXDuA1We5X7RqEghylUVrgUuyRpoXDZtm
UJHATR3WV961YG7EQSnreJhZqkW9zaPgk4a+slDSspLZvX25jq4ASNEoolqRfz75ZDets9Y7twLf
rt1AmEso+FQfh3tZHXisd7B7q51dAo+VuXaXs1jBVQFlgLvTIfMbdLMFmtz+MHATKywcPq7myZoA
yySYrnVLolcfFOuVxqKU1l7NUDVn57qMGPTlpPhGfMqp5idVZWD7HtQ1ycLA5CdyvDZPNcdSNb/f
9mKIkVfpX3nvya0L/KE5ItQs+6ZQMEnOZ0sWHfaeRFxrFfZXOlDn7WyRN0l7Hvj6sVHWDmUe5vLg
WvdhGJmeRmYPD2NyBEcXv4XV6DzkClP2zoy2r8DFZIyKrAyPDqviTlfyGQn7I9nzADPGBVOw7cKz
z564p7d7OsmmN2MWJOK1rd9KCLYYCemCO6bJjz8mAYybOca6oE8Gnkpi1BoWi1V8jgBuXXb5rIl5
mDVfl42nyd0zmuN2YEavZAZI10n9psjgujdGLj9TJM+nE+q7bvsvL+2tegDf8nsyIgbZe15ShKCC
MwCSQC51mLJ/TCb9QpR5GMmaGjlEMIf2JSIXaIdbPzLfX0pCzHJVY8yBQlmpvnCwPx5DUQJzFUqn
wUnHsaAQKPDsOpgvZPc3pSaM8/ayqVEyqDUADRVWXyOAEGhpECVrRzhXExjsKUy7RqQ6zk54srCG
4/PdGCIIzSXMBW8hsyUaj32BwscmpPkMiiaO69AlnXE+yfaOCEYnla+PbE4PDxYQ7SjeJZOMmyaX
JULa9BV1W2obOG5aCij6bE3evuhVIlk7t96iGq97NJrQEvmIndWRAyDadlwdTD7SIC8gLG0tykuZ
WqHwiRruHqz3ni3QKd9awTyXVyVzanK7SoqK3CUUbxroZeBACqfBGj+LAEQgqdc5V6/HOw+D6izV
9BdGPgRRi9h4M1Kl++qvekW2W5oMgqCdzGk0S0NWp+hHB7nyrt+p3OCziFZk37tV1c8+0usRnQ3C
EV+ORzAOiPox3GhADd7fkQQxKZN064bkFLl/7n4BHi6whhJ1U/V8oIp2ewD/8H1eeSVi3AbYhCoS
aHTuxmQ/iLahNTWUw6WdLB1/GBDCiFX/gbhwXANdLeZgII4960EQcw2baR8t6nVlRmVuxPrCI65o
lBspX5jhCqJhON9Gcsp46+W9EZAUUVVYCfvJfd+oi1kSl5oVaIb6ss036DE2cNhMfwKj1BIXPnOr
+zcRqkVZ1Yt9CbmIdPQzw/9jONgxNaF9EbiHjOWuET2XkQ7Z+iR1K5FCM0YnHlmXi3BjpFse6DQw
lwSBJ89xLSoM8htMIGS0BKkk7XrjySoRjxR+FZxQj1JQHrTslL4fGUmLoiH2bSAasTuEAt7SpZTn
eVoQZqxKcLSLXK5+atTQ0BQM60A8v0k5anAgj5LPd2sUT7fxcWWBSU3V1bDzfwUexKVpyAjdcfBB
iMILerECRhZnmAWv4VfJtJ3BY76l+zyFLvhmLqGkCnt/iAv+F4EgUld6MfKkFv2+oIfi6jTX4LmR
O8dX9siMgLrjqUIxAl8cYz7UyRrppmE0job0fosWwRrEiDxVUwNZSQhBt1kCHQ8BXeE4P5qxZtzx
mBCbYvsbW0Nq1HK0aH+4+PoUWGTlTMqWzpZciXVXzgUW4HLUaq6D9gQyVg6X1DEWvWQgdy1rWrPD
/igT4FxRLayX3GSza8SuHq0D8OAdY5YhFswGgjoDnYIoOw9WyhZucRpeppi1ELxGa/vZSsuGBCE9
9iWPlT6UZDYN+rQQI7WoHCRhGGkHPZawrsiosx1H2Cm0bjdVWN+ntfd1mu9O5SpxUM0ID+2ZvrRi
oI+mAgXOJCsZKNU9pQ5vlub8OfEk0jTBA2/xwwWxKZgCGI4ObzGjqVU4OtO6doMtuMHae+143ZoB
iAKVsajc3tEZXud2/Wt324ZkA32rf51hpqE2vX9igQFjjxT8fffz7/kt0tHJUTjduZ+PJnZ15CCm
CCKmwjUHJKqfHgd/KlFE4FdZQpptYEtFFizFNTtocZ6G/EAHBZbwhFf0LuQZmbfGQCJYFR936M93
cAjW4S5Htf0bOVtVTLahjeWrSoRUO4mLUDzJRr5wSmrZ+GqdbrRkA2At6F4LtH13milRpMBJxpga
CLuOX+UfBXeK+sLVsMIsSIAFq4TxIuqzF8xfuulSbh/0CGuhneLCu4Z6pmB2umaLCJ+LkJeQYiZZ
PFN7YjjFiMN3Y2y6Vi9L3/UH0bFGQbPvinJ14FzJzglZvme631wTRTJM447gTHrAUpCVYFINP0TD
0MCkXp4RcsJYiazbmEE1dL8aFOrHf/JM7f2Zna0T6nr+ZTG9Ya9q0+28EcRuX58sI1d8UQU65Atv
IcEFGLz0g9ENtoDc1OiQ97aiYal5ZjOUuTpFeWW8OqozMrepCmX7oeCf5jcL6G4yQfemOUk+RLvR
NVJu4mh/GjENYX9VLcj/SvN6swOsaoKfuVf7GHhW8BfDAU2DzCZhqIrCWKfxaTb0Yl3c9O2R5F9L
IqvWrVevi3YQ5HkxpJpog0fmN4E8njQCG3rfdyyWkrP59hIkrUnUiwVNLaZwg6jJ8cyvRDorOu7f
KdXYYgrEcComrPCRig3hlj4gZMX6BiL2qEbFNjvZAYAVYJGRVGNt86BjKWPrivUOZOypXTClt3Rg
pHGoNxlPpGS8xYLpgCPU9tvm0rOT/hf090VWyS0uRFc3g3bO2gmmqUhtFxrcmBuIyRzF3MVsFzSz
AmyvHhGtKj4DyZ89wGzTp+CRyRXWHUvLKepu3whrfZqMIde0rICLefjeQazFEXRXkPdhgqE4mMwq
cmqgOEgYmKJduWWny56k7wESt94WMAbOWXM+4GWGclRvB1/IzfVND9QM9F2IMTuk05QjF+61HHb7
l5zvQ815+jemXv7CHn8sriGcKSxS0oOZmDJ+YbW869WahWVMjDKkjIGuAdV8YvFLEO7xjuikT3tX
CcPvr8lM9cSRmyF6bnd44yUFFJJbGC9PQKO/OxUEJMTj0Fk7DRWhAsmEvPXOnKeH5u3wPYjc3SKW
LNHAzja0E4QL7g/xUobj0mWw8NfYibe+9VqXAUSMVcHFNDyAHgpM3BVpiNypljDdiXVBxbUPRrIX
GZQi9typF/l95E4gKeg6dzOa8vq2OZnynzdBBL+bTn0lInqZ9auKgjlKoGhFCG5d3XAi/2uaaMVf
drsoD+FHlYOV+CS/gISTUjCm12dXGyIS8Y3uPZoOyFyyb7BrKmw7VT3IOMU4jb3uNPLQCkFjHyqH
T+Z2822IKaJTxfPx1+2ubZ+nN9bQtbnx4LuexaZ2Jv7uBJ24Be/LKoT7fvgycpWvnb4jInKkS8W/
1jxfWAwdJfRS8pM7zmNbbIn4GflYw5lWZKB2+EglsVWIzrP41E194xHamXXtaBGXswtqRfeU3+pB
JaKryghtMugIMryCCOSZH24ILbZc5bJPNtD/8mvOG2fiJM+UI85/6ZA2SmDatMrWxNen6NgQ+hoh
UmY6JlzUuT4OKM9KM082yJbMzQj5/boa5oiLYPTrXXpKtGQc5nnruZYVUc3XV+1OaklyTCAUbDhY
Kle99QOzXWKO4jXylLleaEornQZf6JeuiwOn7SHNcUkNbUrKF9XFjR5/ISFFszgPxvJr3H44deG0
HNTQvkIwWjPyl0TUbPlTnG6fYo1RF5m2L3br7CSxh9aV3HUCf1m86zDDn5gKbK+fClpp4BGmfSfQ
9IAD6qdMBzu5iwoTk8452Xboi3FBFfm5WwAWgLs/y1jHOBw9vL8TLjQsdSKzmpNSpwwC+w1UsA2Q
pfaGZlUbURtep/bfMewME2iUgLjJeMC3EAsXD5ZJnGFL6Df5F+A3gHc6TVIzy0p16Zfp7CphDYXS
U+qIp23JRK8wxlssiB3DtTWWL0cMdE6bJXqRr/bjv/uuy6FFXTxNCUlszOWlp488IuY9PjLCAKqX
56I4ztbFipGoX5y++PuwbiaBmaOdPPE32TzCYazrALiI94EJBuaerk7p0kuO6vXH8iKHqnsdkBo5
cimj8HK79hWXR+9ap05xb2xX9pjapHNWY0MSX77FP0N72aAJj0bXXK57oaDp4ksLo2jYX/Af/cI6
QHmoiF8cPZlpz0zY2Q1PPYRpfhGX03kEDuUAh4uNSkAaT5mP3cjwt94QbAfCoKoVO3HlxgYVkZmp
0qLnNF1ayVWN/Fdmd7WPC0pMxcTbIij+fyEDA5pxmAntdm05BgoyRzFQk565Z4dw3otl8cW3uJEG
/I5E9HKe0+DRhB/2X7Od3OQSCuBu+YJr6DeXvPAHxq34v4BgK6qxU0bih/f/l3dL4yoHaFtme1xE
buktvsmAl9EhJqTOUpGSkg/X7Z27UsXsOZO1QkFzclF4Mq7CdLCtopO2PSsGbmp0AQ8zUM59GehZ
6yjasPXiosADZ6RMap3Y26PIDxr/E3Ovkf/7e6nkD1q73aii4Ck/WDRwJFsESQqbO/oJV62/0qOH
SmBzYLqCTzHGPLKdka6jh6Nw4zC77vnGpzL0qGO/NhgnUsm2xfeTEOtf0MUI9LqCW2A2SNO0l9h8
FwHL68mQ2dypjpXF0O1A5ZLHJ+xIT/H12q8rC0IqQ43TAmk17SSJ2QdSvEcuxs3GWe+4RfqkTqqK
8QPxSzMZ6I91u5AGC+xbMCPYafCsKEx7SRdJJXV/H0vTCBrOqzHu6ScCcgRUWAmYnKidNuBEhQrk
z58B4+UTKHlsMFHWdbHVwvATigomwDY5KVMy1kNDq4+0iGOb45G3lHpYWrV/+Sz5wPuuP/eAoQqf
oZapNFIGFYrAUhxnTkxJL8/Zc+fVlU47aSt1mNnIlh6GWQe6khZQNjGWM5wmGMU4keqD5wNi3FUa
VTG3vRFpamABzmgzHAPcIVLjbCv57CXNIQCaQcnHNSYgNBKinM8JRLiwOWwG2Tw9NM0zhV6G/wuw
pgKwsCue0jCj5hXMsskOTafeaX3XwFv0dhYA8gdRqf1j/FauPuWo0yBQ9cuShVFtL/2FD84d2hGW
Eg18kl5haFwqMDBT5rO0r87IfTWkE/CCwqcJI/z0eEuhJiBvFh/7AbXZA+oaRbntowga+G8oRM8v
fUdE30qd/b7raCXvC6GhesyBY+xqkSXJGtE609J4BFNNFFo07MDMeVYds8HhMIkAVet1PMkUK28v
Jd0FSwvHpXQAsQF6OodUJPxBQ8+mPdVV2FiMmw+A5K1btm9Fxcs0E7oTwXlPKktBPpjKM6WdXV6E
N4KWsb/uOBpoO/7SzLU0m/L/i0XXMdlyLSKhA0+O94As5hhT+FB1Vq5oef5y3RIf9umR2A9dNyfo
EEEYpLSqYr3Qehb/+Qea+berVgC+MegniKnE11nDW/J+P0sipyvCeqrubvIXn4tqsquUu32cYIor
Y2dztxjABPPLGiAs6lAU02kDDv5zroutlF9LojQZ9cBfj+edEriGsqNXbtM3D0dm2nN3XyKLC+fA
NKix5hcZ4SbDntdnINPit7PFAVYgGJtFUNmtY+crYcrG0dz5K05dx5DE0KUMqZxoue82KCtwVKjV
WWKjWSMsQMXmhNMu0uBupDEytbfc4UFUGqCby2JIagkfJx/A03U4ASaewsnF5ImceSLVabP7xA9w
Y8I+IOKAwnARFQas5neWcXjopoeSY5wKMFOVvUZykKOXIDoyATLzeUtwZ0eoO3SDCarosaBGDdy1
lEqX3TrAeYpk9oWcVRICMvmQqSybiNmzUdyaKIYReqIBg6/ldivwUeeCp1zh3Ps1C2YHOxPWyPAk
ngYatuylgz7v2cSsJp7HCtvIWQM8kOPnpXj7/zgjOKXxtdq2lsLujJQ9pFwcI/Au7jKVCq2x2Xvl
yNimoyDMKPLwZ49OWflgVUDrGy59frXnIVZXfgTPeMyiQkPPbK4TsHxpFcB5zD89uH88TdkzQQn4
d/ZySpw2kuQqe9nhmtC4Qwm67S9X8jqZ90NdOIf6ZOegxJ/l+tXtfSJ4lIsp7WLOcEIUbtXtcUmZ
F1S1wd1wBXgPiZXvlsoqcU/dkVK8Yb3BcMiH0WONX/m59zfpQ0/Hdn7Uxha5MMQ+QMyWO5upq3Rb
c0Wiv7jEB6FvS1OtuDUoHosYSd7q3srbdK0XQXKlX0DYbgdzjkheo20t96NVcZhp671dUDaTUQmD
gjjJRetkCHL6bpN/QP+S0P822Un1cGDU4zepR1dGofpeYO7vtryMoH3AZCWmZTjwbmObFWoAQYXu
AEDbZZ3CQpzPszH3rOW0h+cKzAVoVqOlCzYp93Io1/OIKCz630ObwxTyVb50rkltC9MjfTFVJPnG
lsvM0PJwETRyx6gFegzL3CCYYAf8ttOdIuh2vtS9WEXvElQSyAJabgd3CDluugk12t24+bP+bdHo
UPm6YJtVQlpoOWt+LYeaSR/9RSmzfLw7/sikmRUgpDD+ttmJpkYHCnRjg8dlRCD83UduOWZzJXrq
3sHZPUrGTCKdJF1XOlaFAYC2P+EVlec0Bg1l69Suxniuj5++UJ+7ToCljLWoma+M4TZ7ZD5kdjwL
z/Dea4QY2QdYR34velM3V+PXFCr9zZRX9er2IGE89fZhK2u9f2OcxL0jAcipXuhmjhpAFLT9Md0d
qEGD778NQSblUbNAictiJYrWcIvVyRllSQvVkTnlyKstXlDyJujzNFzdIVsnjze5AXXeu1XqfvaB
w6JhIJeqx7BIToozJtPEvB90NVMNmROaZRP1mKF91v0ESxa2a6ksCfPRMPxTvYkiJgcR8cK9V3rl
GhYSfvq+ysOIsioBEAIJXyYEFGnjEQ+18s1SsQJEQhg5SJ0VJkRKUYuLUb+DAHcTgZ+evCcAvVTx
ImXIAEFvkmkjU/xCKcUckgKGYWYibI2pPfu5NGWEB79Pqx6bKYlimLHi1GjVcdvZfBeU88V8D6pc
HSrg33w26ZeRsX1W+RAgIxNEgmH7E4jjbWx/748C7XJDsPwEUK0K2YWcn2Rucx2Y34sldU1i7gdv
lc+F4D1R79PBRJlH+tyCu3o4vyZcHKUOEy7hi1RkRaKtLvfn3drXOHf1UsM+fb+7HIxN26JS+tQM
MYrcjJWbBGgBJYzuAKk0JMS+0COd/WG1AGUjCYy08qNs38WqFP8FGBIn1ziUFQhE1hvMSSRk+voV
7zynEWq2WNnEFLtfeCNpInMUuG2/rjktvarDjJ8caWjVvGkak7BVIjuzYOJV/X+pcIwiMy8QpPUs
RKLQjzeY2PEN2+8S+TdscSJzJgUYwrLlEtf2r2O1m3sOOfRV5DaA/utQZOIh89TIM/VYueCScWlT
2RwIh5yDvvAwMhVA+HGqmNl3DgAsAN3Mvwmn9qoLCn498M+otK47ER1p+OqH68P0NqgU4i5SaTXY
7XZD5oM3avQWGoA71J3BGdmakQDg0BBj3TB52j0upoq0vwl1qZhYco+c8V1T8xXuUo3kUbKu+znR
7V9ImqX+bpmWqPntmc2Iu2QfVEKMM/F6HUwcNZZ5gSDllwXMlr32VXW7G/V0y5vB4Q1kwJ/Tp0BR
KGyVU0ot1TBej4ThWEhVUZ0UJjpiXYYn/ZjqYMMCtl+9+Qdyc/tjvW9O3i0RRT5XLQ3plY/Ybl2Q
kew92ut+Pkdd3J5MKCGpApnnjYI85zCu42Ex6S+V/9ib/rKVJbIxVmVajXxjYyoZfCffQOC9buZK
Ygs5GQN0DvgFBLiSr+LqBvcP7ZCwV1OlSNCM/Z4BFaLGuwM3wRf9MA75TDB8kzZzcLelrIz5z4A/
L49QulwBmJZPkF2DBYmL3UdUT2M4ht45q4IdUHb3D//e6Vdcu8WNvjmXd4pj4KlbWvC4PymWVdmM
m5aVOVuPB/JjEO3I9QIEIlonkqabFe2xY2A2x1Tv3QDGP5zkdN84WxqWunmYymPv9HVAekccDh6q
oIN9YFijIM4/SdLSFxpjprCbaIgiyjxflAT8ZfM99p9fOYBFmEFQ/XR7DDBuXgP5fzsAhK/C3Fiv
kYKUmtdogWpf4gHBEetYLUuF6cdTSCQjEYnvVDVS1DAln+X34EPCtDclCreVOht1UiWhCZXPzwIc
0FAhbMvNDCctKucDIGGr8YRSQs9ArQrOk5wCSBprVI5rySJX5J46HQyX+rjO2WVt3I0ux0UASeVk
evILS5ZFkSqGxW0PAAZgXpexXbV4yWTeUPTCJbmdELGihDO5Bs6lzvhyKBz67QJNFHS3s0KnSdVP
LNkre5fUA0YUh55O63tgEigmaPE17bOmFSADB/jNrDHc84TPf22LlErlr40fjNsWVflAYKiWqTbv
Fo+vuWSI8DyU2fBgagkpjczwP/h7ZFvKpV3B91jp3ihnC8H8/wFIXdGX2zvPqgHfRCl7Vn1B4lFq
wU0AhYcD1RB4l6qyaJ1cjE8v+8uEao/vTHR6Kkf0Zw7OMQF3QMjxmnySxkgEZ0lOILl+WNnhVflC
flGfWPm4a422qLaOvngepIeQbzHwNGpvBK5TY7m33ecCVBU2OHjWX+LaW/DLwUhQyw9yaCuiG6KP
L6t6cGfWtDBUcuOJnNSit/xI5aIJcjnWTc5a2p/FNDzW45d6vOwo8Mol9vla42QdmDQFZGxC6uFc
HUryPNbc/y0ctyHTz2qilVTSCwmVWiUSfC8Z5u55H2Q5+ZTWi7OBnxUrYjPyc8rvjV5IhEH22KSF
bUodiynm3ERhPkCeRsLOCCs873Rtd2KgENPEf1Q2AYVQRvCyxUTJ+NRjWMh6B/Hig8wHNL+8qqcp
08yJJaE9M50dawEzpT48FzfD5sji2NMAP4SHs6BdLEDReAjYKM5YE9LigOj0V/hIGfuizE0fc745
8Y9+6WLxE99FGW4H/Qiz0nSoaUuj2uAb5kGhQWfAj81OZ1r3VpM0YXdAh1N/ySkBB9c/U/X7Cl4l
eLdw/pzIunkvkLHRNma+XPu3TpxSXkfeXN7MjX/X9PZR3ZlfNryaJHEZ0NCkIuaVDsmiGHhmynH0
glUYyV3TNF08qBPz37HmzKAfgd+UX0nmumGij5xmuwLq2FTH8L5XCZPHgvD37SqFZ3uT+ydxlMiS
8MJQ1jl4zrrvUYwH9fw3n/mvXPSq6aZ2vy+XNgmHWB1q5O+JWbse+EJsnF5PYJ71r2gFcsSaiwGl
tZ8b2pUw6mM04AdlUCFq1YIDBZAnZAW/94en0WkVmyfiVb9zK+68iCBJDuaUNZzJ0BJj2TLD7q3z
Ar8nBSzptU7wtpEESt9gxN80T2baUbDQ7vHX3PoDGHzoQbhTYfs8mUv2Qqtco3PGJpKMnexguR97
p/pj1+2FvQtql+0pTDJiv4hOX1QCiUyNA8A4rgWqzc4SEAuq9KeILlaRdCNPpeAKz5Ur9eNpJvL7
6eI3vVLvyLo0KVGTlRcWyMLePsLP0DnPkLOKeRp0sQ9w/23TW3HrtK5zXzGGP/4YsX7BYQIOiOw4
BAn0C6WcGjZ3YmhOtM6IdYyoDiOvyRcUgT3Bg9W4DGTySNcq0BRu2qbvbgxjXe1ff8a6K2LQsoWt
eg2IqpqC4dwOtYgpKcxN4A7FZKVVl3WkwSgkY8fs/N9qAyV3P5O3JZMQGWHQIvO+LBhb96s/lBSx
eBGxcqq2dx5cyK7hinQ0dpY/e/DtBZkp4nnJx8b0dEhLoC+T9pkjJ4kHf+1oMv4E2ex9Dma7w+us
PHOzOwzT+EUuHZiGymvFxERBhijr7SoloU30M2yHem3jwRR7S9+rxe1xi8RonyIkk3wN58TnmG+C
ODe/k0BZ6EYv39szb5cmHvEM5/d6Ww3L3sMN9PDjVqCS7c6f1VMtDD8TeW89Di4qr7cEMPbj+rf9
ioEYLeWo2V6B89/uH4f1vkpe27nyT3p8xj9jo6tUFHODGSQtltjsGW2YKOegKJKeBEMhLHLJVWGg
361ozDlAfak8ZISWyrJy00VXUV+3WiuP/bYAQZyGjpX1ic/bo3wSkwpF8wJlqc0/i1SGlDFlf2JH
RtZLbqRNL7c0HFN2D8jeR3z7OAhpWFYgrWrqaT5jMQvcV+dDrwzq/i38t20k50ryA9Bsf4aM6qTK
z4TLCgILMPCA0up9FqCUNqbNdfT+R10/aXuqtwDRkMG0iQ8W7BNOLw/pcOqTV1agZaYnCKitbtzG
JGBhIxvEIiT7vrFYMVROqB8hyxjeyYeIzmv6HnNwE5jMSzPN0BNLgxsqbASLdM6l5ARaCP9M7rKw
gf8RFWjovFwX7HKP24/wIcC8+DD6iXEXBy/KqHAn0foBAISgRkBTKlyegmtngGTGGqM0s4WA9A00
B1p83BWsuFrvYTLsbosWka0LVpYe2K6xp1uq3mQbfQCwGcseNyHLDb64S9nCv+8D1ISz5VBGWpf8
3W5QsRfTa94BZ+Q1RMxW6QDjsiS/B2Zg1UIqPAsU7M9CKjvNTaSBQrtPRQGu9V4g8UnAlOyMieRC
N+le+YnCgRLt7ijyy2vWoAHxlQ4KpN1SGMJOcSJRgGaoSs1fykROGQVQ5h1uA79/2tsBC0pyaOA2
RnszpGGM0kLB8LK08gJf1T1zcqyJZEmYV+JfAjeP5eFHjNIIILJUJ5nC617Zkn9MQii2kic+E6i0
4R/E55OE2bB0zdTb9RNSEgEZM7XksGNrH03OIcGsaqvt4xnxe6rMLUFLjOlgeRtjZi1i1poBXpFV
oyLEQgudZRf8AZuBo1zJdUjLrC91qveP9oH5//arKFJl6iLQlVUwZ1FfsmZvY8KpXA+bPCHEVqml
3Ylo6uBnn52yjwIhX/fY52T3tjeCITFwMf28KqAV3zCW6sYKFCQcoURv5NUYsqrEg2OkPOfRE1hQ
svTBZz/M1qhA/CqAzrOrh9EKc1z9ef0Q3j6ePixtf0R41iMWtspRIhvfNr917NQ1m/e5h3fvKutA
n7e/Po1q4rvdGAOA1iiSMzk8V7jCBtv5yISUuJx6PBg67pYN6TH54y+wHicXXRDlk2gQKeNvEjTr
IL1jPvzDUhqBZEnOPv48TqGVJ8AR3OfbmghKAz0TFGiEFrNXVFxHz5uVYTIWaUPcbFaxeaVbQ0X1
EONGr+MDjMPWSPuYcxE+bKVfRJSIvRzWHXVwZewC0grKLnvqw9SUBOicWoFiO3OoBVHaymQ5HN5R
j+MwIkdKKv5wEEBMo6CUx8LzGDu668yFTzqf5Qr0D/BsO0ugKzxWytWpnuqV+HeHlOkZvOCYvX6x
AO5QiHHFAUeAAdD3uDgEZkFaE+mXuGt1V3/iX8ZHDipwgkcQXfVgkXiZw0WcG3qPHr0pO9I9YhlS
9JErMdIckD/jHJO0toedkv5UgwE5BR2GGdqWmK2RGz5AGAHqTO+bk96tlhkP91rGYFZzDu5o/ax6
+giADB6sJTQMISV/6lBjsow0LkJ+8Lq3nbyhWVJIgGSltrIoTMGsR1+pUXFgCGch/0ItICRE91j4
oyKI6lSgKv0M2Z1SgIaefxAaPXfNZGuFM2iaZviKz0w3SSx+L/CdF3UlPfLzoFIAOBPoU1jcKxc+
mljny+mQ9YsU19PGhz5/kcV1zbzKmdS/uKdDKpgNXKrhX9g8vma9HXIkKXkjgzvIBXhmvfASr/RB
RouUBnd+WohM/O8ByIl9ZSiwpfOQ8ZdMoLC0OkzpQK0cC2QHWMxc9rF6q+9JwWlQMuT7NyGYx3V0
hveilVJtsM+MraJ7C3ZiCFFwGvsv0HDur+i8S0N7KUwsWRnVFk62doViP3c2pc69+kCdtOStfIxr
HNmG1nbvPxlMtIOCK6sJFM5fFfYGZpbivwrfizwowO+pKysbL0BKQKuUEoeXyyTgjQrdIekn8Itl
Xk25Lni1pY6BDsE2VkILkOI7C4dBeIyi3KS0YYrLlGfaBiqgw2EvUpRsPxndRGGwbrBKFYSDV5IR
ezUMfgiKx58J+dbfHUKCGKk43fyKS11abUIc1UOkbMHyg+d33FOavjBVtqaseZg+4MbHAmxv77tV
7OexLBUNah1darJXKUEaAVjmpwJN0VjBjSUsrJjYKs6Dvmtd0aQ2YCwPk8d4sz3HpnIC9VKsY7+2
F90ODnN65C/n7zDKc3HYEjsnxET1+b5Jl9LEPojHkBjOjU5UIou7JpPPh19pr/mZfYK0zIR+OHnu
zgQ2qPekUJ2m9+s2sDr89cX4koLzXMWa4o0t8PWzqkl6Ho/hfRoOlOI9469SyDpy6bXd75mxpSAA
SI/t0KpEaFQ4ajeHqAZAeBmDuKhROHW3eW399xH01zWACo9q+m7zWlLmcdjQrftkIBNYWZqs9WdM
EK/VZFTOVYmbeo1Uzvu6TqXYKUxL2kwMA/out4G1MkqDDvK2nJR8jeOY71jFxPJRqq56stogjDHa
9SqSt0nX/gr7/iGRJ+lwb5AB3/uSL6NnKX8HaDTUQpkihrNFD3B5Pbn48GbEt76mUXKR+5HXyWvP
hsRtB/k9mmgUoi7/5csJZUa1DE5xglHplPqulZLyYnhbGmWHXEkFLZKoA00ijdOfYMLSefJ8xmp9
2K7iEyRchPFGXc3/emk2vlZ2li4kwn5TpJ2PX6KTRLBtd7WxI1MvCgfwJ85ZFSH/EUYJiF9YMNnb
hRmuoJ5uktWLp/tYk/emsOILP86yE6NtpIFltD/cRfWspeGBA8LiyS0YZJjobilo6udViuKzQeRQ
BLKld9u+FR3TnDSRr/1iFQb+lqy5qBWeAcCaDzaSopN3Ylgl8PZwz/FUhUva7hOuNM39tI+iKYau
nj7GL1Un8FWo7EV+2WRPH6MuhjbkRdq7i8ePZXXbLduaW0DS5dL6cDN0+LQ19X/GGRbSytCbUZzP
Kf8pYEZiY/ibyuzb5Wvm/81TkBlRSahTUqd4rnCTSVnGRE2bYcIS3sT7foxrCJpjmJq21Xw2Zx8S
7yWckCYVrYZjcsbfK0GJkQNEtGFSUoadVLOdfiXut6L7rRNWmkzVBtKX3tcKUVWoKufZB5hxWmOY
8wzBKceyObyIVW84ZaVUl7WlA3JJSsqBlGduB8qkiwhE+jnQSgTZQMRfRMvnMG/SQHK/eUH0ev2H
iIr45mnvargWP53Ldj3wNmYIjKXAFbMd9rvWiZJAR2WB8iBHXZ/is/vzicTxQ5QtkkuhttjNHnx4
KQv/QJXfr6Hpe28O0c79yJ6OZFbcEuQ26/fJTOqNBzGxdQIfGaTEFxNTz/X6lE0BaaCcmPVX5es8
2qkMOTqwbjjJCtRqZbZZHud6+PvRvj+naevsct3EnuWh64Pl1zj0Uj8JUOJKq8MAEUneDb/IqkiL
a29thRJw/sPxSOHaeLgWCYTbDy/o+xE3/EVYJgvv18fVIHLMJcVxnAADc5VQH2C7X/7nuijdqp24
teUt2/ml+PeXcERkIOodfTHJ70bHjuFVKp7TaOqzPLHDrD0wKw+TT6oBNSoyEVEpzcW52t2EXHje
oAEwIv+7gjQkouQ6rX0aauJzktIZ1hAfkZLf0cfiyI10GtcfRi17lElhsKSD+HHb8AD/9ee08DnC
STRMLR8I7bzrhtqFZncocUSDG7MnSDFVFD4qkf9ALsR/eQA0BNx4+1sfKxD0cXSrnOMd7n2PCkaM
Urxo5nj8MBu+55ekHJ2McOB0Bs5qNPa/2Z9knhPT6RBRWid3yCcS573d7lk+FtTwFKvVhGHFrXO8
KdcKumQ1KW06VtNkhzrzOl+K7YfWoxSYjSsGMnvGSe4VVTnRTjFAxtF3Iwy6DyMgnWMLx5kTvhx1
fUQKRmtRtV4LTiruQMiHuVk2AUptF8HgEMIF2PakpvRmVA3QAqofJuc9MJuq4+KSc7pbQ8peylPo
vXfcQzXvPO8JNARO8XmgHGuJTINkL4D5rZ2zfOlD3FSEFPQUEpzPrQpG4zayiRtkuXmgHilHz3El
5Z9L6ujdVDPKJhTBog0CyOXnM7ZK9davrXI16u6iifoXpWBn255g+4IYWb/e3XQGMCopPMFETD24
IAhdssFqK3/mSx28nSBI+AzuiUJ4gid33FOHek1hEIRottYAu8LGUSRjmJy0KAYNPBflbTXfdgNc
JesekcozIQUcDcUwpZKSGVub98uBzIiqmbZm8TDAs6wSjIAF+T7hS36t3URzh7TviezZs7AJUwz1
B28AqBuSOGBEv650pKbLsckM0nhD6mZ41jbcpIq/P6MNXYH2J7EBaPUjci5kH++r1qCRuKKEl5DT
YRBZui1WJdhrcpJ9vnrjMlFm3D8tzo++mLDqwMPy0fJm2tE/YWpET+KLhp7Ah1fRmCmXFkpvLnBj
BGSZn6qsydCJ4l/cKKQSCv3cpD5J4je1QltXbLhyqUDSmtF/G+W41EmZx9zrpOD+a3YoPKCFk9Vl
9CUixDk4RBoIjVHRs7hseCthfBjvqjTBkwkPdHJyFTuZAlUCxo9yN+r/oDfH+hjzZK/838vJZvCd
pfzIVbZol+AQpqA4Cz/vI0OY7GzGIuKIJfIiLwwjOieHC9378L07RP8b4KcpRKlIuUe9b3OO3Xay
N9QiF0EV21c0tA9yqQglWj+yJ4S4OOA+ctVJg7CsDSOWHh6tdl4YafCLPfEyRN7iD5hEz8F2npEF
ylsPTwuSUnLHzgP9WxxSu+AVALUjYrA8Tyq2pf8VEh4u5D49tA4z0Pv/TA+5rwexNOEJ8cdHYLJf
kvvpGXYtCvCqfwGNB6Svdjwnd85Y5b2H3yKuTBswyBdq5fezsaOAbgXzIy4+GQns37NxFcjusNz7
fTIn0B5OTHb6oQKMsntOWMNkCFBKE/5k5sERCH5eB9T0n5qJFnfzaxUWV6S8HhBSK2RKUw3w5o+Y
PprzUNe9MT8R8Tl/Vm5VEKg0qLpWNUeFQkiBl7HL6D2/bT3hi2Ng6RxvI+GBjO4aYNQ4zRxVkxh5
2DsY3thlFfN4uPpz6pwHlpbMvZWnndDC4Gjs05kIiE+eT1xWPvCC7KuiXpWd93oxf0T23e+K0pER
t5mOl17/V4SIJN2ltJ7K33CfLAichbzhzLo9oY2jEcDOxe7XjLm799hMmW/8s4Axf52FNyHxtrEu
A00kIJOxDCsI65yiobLlhAmzQvvvt3g3OurBISD4GqeAkGL1TlatJHpMx7/INFIV9LAXxe4Wkj/l
GpPnHMd4rinZBZJqJiH3+M/a/mLzfeRXWI8+rrne4Re1LLP04fvYAWbu1NIjWkulxCSVEy/3VGgC
HatnSsTua2xq8kyY/B4Dbt+42B2GWoPsuysnvjkq8Ko/Gj8yNqp5f+bCdwYGt82NZrMZzm9DuA4U
hXg95Fpc/HMqBHuQ9iwCRnZ1kFUlQA7EwtaJH6gPlXyRlzyzvfsI4YxvKRAxhzFY5e4ISiTSI3gw
ebb7ffo3l1S0lCgXus/4af+3R/gf08rJnr1b9nZbpFDj3wPSTPuEKZtNA3SlNl0OvMqC2va6ows8
AMHPA/ObDk3ugx926CfKhCDLfNF4fvHpZIAbuoFADUuoogT5VIDj7gtTXPdvkMecgijET2l47ERO
lquOWE5unbDaxpSekd5opPBvoaLMgl1l1XIgEUlwk7K8TMDNdyFBAE4wPGREAxp8Tz5nTZw0lYfr
3Q93NAUOeg+zD1hqQqY7DFiutfs6eZjPFK25q67GwUqZAq3YpR+2u6V9lhjNUssqCz5RRtXjCmNj
5pjfpMTYIR+N1d9mz3slM31u7zDakboK+PZQfsohZxsvJ71wsalMjlhJ+FVZbhlJ6N9UIIA95ykz
F9GW9LBqd/tU6N92G9ipx0P2Ji7cAEPUzPtqcSiFA8HGKYz4pYBi4is504Pj+QEIFDeRR1Pv8X9K
1VpnK7mWfS56cQujD8MvB0aX2r1ui/qHmLpdQfq6Bvs3mXE2pp1YgVyyBZTL2aunsRrajNP8z7FJ
P0L4hQ3tn4n1ycfGig7RiWAg0Ot9zCLVpTy+2hlr4C9bOD+T7zNvOxhRZnyWyWbRSmxrw7pKa/nM
9X0bxuZLR4zbdnzWgFzB3RTUmYizlzX4H38HKwLxvZdsNmVIFNz9RkwQwGjS5+uzJB8IHpx5tgRv
KMXXeThdM/1YAZ5IP8sCYGbdoX7b9Aaqw+dsOHxwF9JXvrGYYMdiSwY95zAXpR+4XBwzYm6A0/KN
Mu8Wt+wCYAZ8T+ecAR751fOc1COhFdSuDTIIXnnDjX4qrywkV2T4L5IRZOBNAF+/CTgffoSVhQjn
G4VCkf5VJTYiTyDei85yQcS/LfS3LD8YIigoiiiCWAIW+WHTm9KF70q9cKC+nEpVb/Y+fgk0fXOy
Q0SvaCRGTrg4CEN9DM/PKZtzNrxR8JqXALJE4pUCZ1MOpCbBItxwPx69WNJOjnLZTI94JmjLOxcl
n+LWh9ZdrOlFj1pTMhvmAq5GqMVe/zvuPGC+/eTZxQCpsnOfGo86DibM9SJvMXSF6/Sdwseg7E3q
OGoHjpP+YSJLBf9iSs+/hBzbIJxQpX3eRmUapFxLFvgswHLg1rNMyZr2k948E5WPPpUVmYQ6E+aW
6NgrrqzhCoX0iIBZwJge7TUy07WdH4Taaa/uPqybnXyK0gPGZj/B2Hz4TMvSRu9NWSVoKEjlRzmO
MynpMIiIy6LLEACBHEVLGNw/CXvGN6AmF1LmyIZLx/0sKXdXwmBBIgRhZKB0EuXfEVGSYNgecOlN
6C6u9XEObT11Mi4IgtVQI5bJk4WlqYe1hL8yFmvETjDidUxGmPqDSJTky3uU1DEO9MteZJotXoGA
HwiT7bz2ME+EHZ8nBngds9oRTAz3+YncVOuGXhfJ/j4d8MsXAyVG0EZiKi+eaR0YH1ebJHMYwDh6
tUHa2FNSJ2Qy/Rao5aKbpCQEmkncztPnMK1Av7EoovLyr3qgn+kV3M0ju9Ig9sYc+A4Th4kuOJRp
an3lnab//lsSmpMCabHgqJhM2TGzcddmOiEOREB8pr3TCP8bFyH5B9pKM9c6V/K61JXVwWzVpWDV
wqQAY1Sb/sPH8b/VsfF8630sU7qoI2C26/Ir5DUjJBlY3cwWoAn3c3Nv2tKbTnN02FkpZrSUe0dg
EkASH4MzglXP7aSgCPOQxetoejMC7lMVRSFM3tXrw26O+7fiSAM/+zaqHqG1UnoraOo8ObDweMOS
BOzqWmLCDYgZIh2bHR/tEwAS7/668Z0Dkh5nUoEAQT98RSsIIUvs7abBUUPaBPrHPny+tqyHA8L/
OzQSM0HiFP/9NivYxb6I6arZRvIVkmE+9Vq79/aeaUe+a3nRmHjSamTzeHSUgzasiuhPokbA9g6f
Z2kzC204ST4QOoyiJXk4pyGh2OrQISvx8uAPBk7LIX20+vBfnBz2auD6HS7i27kx1Usl0oq+pMWF
6AUu/m6tmjLNBP0t44xQ2GhuT+aR2VJ+qGXuZbwfURBU+wJHtqbK0guDhlY1FmWf9nHgf6rdUIR4
mofTFGMY7ZvHS0KDhZgbYAqVbYF3B22mXi1mQRERl9VUKTLIBDFnbbxyjhP60bi9cuiNFoeoW72w
+0gbmBHNLutThM/cV0NRK3d3o6xJrgXiyrhnlwx9/BXuICZ9T1ZQyRMRpJK9oUbfVlnwdUPftoDH
BJm7oob63g2qbSfG9tPxDk0IP+x0KD09vEk7/3orqWO5P7DNe1klwR7h5ACgPp0fQnyIaY9TBFA2
nNmI7hw8ygxYg6oPQlNXoTNgVfqk9tw4SJ+tgb+i0+tKdV90sZweOWf1/wvrV3iz7dnbKcCQZgN+
LvSO4qmfUvaWDm06L4bPmPx1W+BX4VxG5oCK4YKriBKMDG4H5SOMWUjCL9BACR31I3If9MonuSfM
pW2JUJyzNvwKMj5Y6JlyjfVJmolkWWUI7sR4Rhfkxeg6swAplpB0vZTyqxyNuNUNIXxryWtxiZDD
a0ZZebSkCKJuJBdo+L/fDfPy4LF0zbe4Um5T9jUq1j4sfIP2JULLubFEL/ywFrLdFKTRULfn0XsS
+EoxaBsaZJ95Cg4jdMTyW3CJyvjjpvFHA85veOkPeNkF++msym9rGz52vAZwL19I3EBbpd8HHrkP
D5jXipF/lXDAHyhb6mraSrgtZ3DZR6EqAVx2jtiDafU4U63VyVOdTM0UjNzuwMoje3nPgta51glg
uJHJ+JyR1HsA56yO+e12wHlYGSkLNjQ5D7OtZMURMF2bvOIElbIHt/DcSevZ2DK8NsszFmHL3D8l
xU5nwvXzCKCN6CHlWFcFbrB9ujSPuLB5WPhtuqbQmotmMRnoB+ijTf0GqJz4fECEwzTI4gtgZtsu
w0kzxtcMVAJ26accqtk1avXTck0FSnJBRm4Cpi/GknkCEMVqzKo8jPOghVc3KfLkbSNo2l3lth8d
NKDGpJpyvjdY809j6LbcI8I0XIaeqQ1bRFfrKMyPRAmMNk7hx9keOymQwxGQ3ye4xwWJQAV6yoz6
leBqaZUqcD/PAyJNxBjZTWLcUdNazh4pz+t+4ZzuxV15pRFU3shng/lxkTTFZtBSML7zL+8RnhTs
IOKyo6jfhpzoWt05Zc/dX9UA6BBiks7VdGOGoO1KcOgbOfqalDCA25JVYqUHla9p7qyvTh9Fiksd
5KGrPcVMdairgAGMv7dxcCYVT/Yf1rXu0cTyeGbOVmP4KurLdKBjAESH5v+swxmrHGjqNYw5t7yM
cvrxdW4aiKaopv/IlNy4ESxlIqwl9yqo7LDejGmQ3OlrAc85YvUHBj2rkPCZjhXH79qy1a9EeYhy
iqdznxltuMWLoJl/zsXAD+EJNGA++hTeSP3bAAM9fdS8NTIOTGamhV5oCXi4w6yJNHDqxitH0KH8
TinYchL+XqMgzRT/wdsFiaJkgxtGQO77kkx8uhtCI8QFFHTRmwBgIH4keNObNDNEfohSNQZmw9za
3IFkg4Huo7qYsWGkM3OQODryLD+L+AOon5OpQJaClvQSW86UEMCggS4CZhBymGvpUMaBtHZ/hoLy
6pJTXPiGO6uQQWoFWyXZCaoSMUnsWPmCL03e00mYx14B1TcCgCKxInCls9rZmYxl8QSNZgcZTGg4
We0gSwTWaTEjR1L+uQeSuB/6ChZZV2SUoHB+ytUih4fVsm3q8X91v1tz1+ItxcOD9dKbfr/8y2kq
/suXaGC6BpPInoaPTnkq+4N+FSCLvhofJGV8U3ofT7R7TaFyEDSIK7S1Gimj8Nva2FoQM20sUjM8
KWaDpY+U9VtLdz6pHsxbBlPwF+R/HKsd5K1FXa7FntTSymEO3eckszEyq79s8WmVs7VeB0/ATJbU
XYznYst3+RUGDFQJ7wLn56eZ8hl/yzChZMWsaYKtgRBfkJs6h27dALQVTMkMbeJOIoegjDqiqTF0
x2Oc9VSG/mi3ehTfViKC1CxDynFYRnjoczN7UBJWfwGWtDIGBX/89QKnev0bVWYAkuPM6NTpN+vQ
We3E7mrKRI9H02NaUjLyIgx+eCOrvZQ+fSFXg+ExPMHh/fXw+5kpuz08Kai9iV+GM9B7k728l+Vk
gbh3NBaRcbkbkf5d+dOC8r1ZPI42kWrrLWv5fd1tikShPKXkROkC5JBXxr4nu6cUKvitrnn6O+In
AMrTff7bBv8RTZ5SRuzGIX2578juj5lQfRemrgwhfLyzM75fybxjmVHMri1JD4TXRt7qRNlERciH
+cLPWiL8dVhQwqnEcp4VRPzhCaMqmsXImn+ukhqlNt36LMhLoqN97Fd8mBIhuNePXG2AlZ+P7BSh
dBPpuyAZ63/dWjxh6OLJ5b6SXS9lJvNLIybnI+d0kYHI5WPteGQi66kGxbkTyZbPjMH40J1fDvTh
+noTtmuWX1xGc1DY5o2OFmwBuHtbDm0zhi9XWhVoRXgluYN1T7tBS4TXPalcOUI57psFpH6eoq1M
IRwIbypg8TuT+xzlLm8/6eR20sfQYGxdcxgLjoRjjP28/k/IpKMTYZVDttzx23g3FRyNBSKz8qtc
8JnJzEDz7qjU+iWcPSQFLwJV5KdSs481IXx8+6j930yKfzn5SYN5N4566HzAZpBfk6TvkX89oR3m
LdjETmeVekg9l47ipG08Yrbu49Ns/7BLL99fWLrxqf1gjqg2UWoLN21FsxSJrtuwzdOn3mLuY8Iw
WjS/CrTv31K1TmmNCBr6DETiqr5dAZPxGDBUPxie0l2aLO6D2UIZlArjNgLMvwj9VVxQHOIpD3N5
1e3AqX1hJMjpdg7emWuNGv4rfobDaapZtfYXXoHC5OifHwCX5bB3lz7dZr8gcCGaz3qW8BEqDyfS
EXqZYv/iQ67h3saYsEzKfhG6DejKo++zGe1xoWlDCdKYXiIzpOm1qevdH2JJw0OOX8opSz+QSkse
1z8wTs0scD/qpKgq2/Obfs+oQjxruWi9SEMjrJw+Uu/6xTE8u7/tasEyw8t6aahk3cRey4VdnHR+
wJc6Zfh/zt47AMtNqLCxMtz8RHt3XQ3K6Nc41g0qFPynSPFs1Gb8a0cMbWmOF6T/DkIdS3zAa7gh
QkYZ5x+efT8ZG/WuvGRyTHGhivBxJJscJiNk/hqN1Uw2qkRlghuogBrvQbaxlt/qOFiLcVVb4vQJ
LpcYyORIF0FL7yPPwCCAlEyCn66ggBO/ZQFOXRm3Pgf4JfURAXxK49dvzxEZnXY/hMkRUsSyKOc7
xDlPl91gFA1oZAZ5SgAwgpt9UNSHri1Qi8d35CeaPEM8X42W+Ql4Q6Vkt3E4fed8m3Xy1Aq/IEQa
BSsTmDmOmSwcoMH8miDHC7MOQnTs4VJh6RzMHQGA1o+M1KVTGIuTNaY5OvjcpgzHMmeltPDb8GoB
7tAHgypvwe7ZxeGDRNDX3sa65eIt1enrcAQ30O/qTsRM1SWRP17WALPfLT3RTPX9CMoEtpd8ISoI
JmIc+upD/ql7cZ9erwlEULGJF/so5O/7OHOUy7raQEFJJeVRk9V6l9nzSrTwtbKSuFgIKYybqCq4
SGitP0wm6axzFEHCtCafdSLujYOWEOoIari6HOUv88XykfSOBZTCTPdyLn0jZvl1D0Lp1OoVcoHh
YdTwZCfirbeZCcC6eff9uKo5/MhtLSztT2CzkOsU8HqYrnLwYPEMZP56kDe1IJNxC7Sxq3LegDp8
UswAr+GNOae4iyIrYOc+SDnjMRlddl0zYQQoH1PbLtnmt1eZnfqC5oU1Sjcaac1TBtVRnxV11fHw
nlBkBpzQR5g17kX2p13dpzgtvTki/ky1aa2fBriggDVVFiOTK9KhSRyvuLSPMJW7kbCeEaq+wuVi
/p/17kW6/A86MCESRACWjvPGAvwucJew+ny1CcEm7Xta9Ch9HRY5jIKvAR7Ca0rgsAqtrdWhXunY
cGXU4E9r93OFZTZd4MfQyGhOd+yZwXt/uCYa17ARXkc216iVz9x97pylKOUkxF0Yeekg0cU0mUFz
3JfCDBWhFcz6hNsUCVT9rksZtRQxp9XmAQV8I1uLFCWcTwsGA4qTI/07yamjFPfSIKwvmYD90GUx
YXPe6DUiafyTJ/iSS6Ws/Q8pT6EO3305Sc5Sw1p3njCY4bW/6jCimTxBfTxbOalBrSFufVgSZLM4
QSoVw1lHedhct1wHinuyFut2lMswW3KxFYd27vpywtLba3AJro8EgiCjN83xnbXvd0bxFy23gXWb
mBHLyd5f2+ZNJrt+kYpzo/iHH03gvSP02MNdGB5D1rzv+GJ2TXHpu3RRkXY6SKKpcBmrXo5YjSdk
RR3ZezR+bGBIrNUfTT/5QedbneX5rhGLLcxSNdt374v0fKxt51HfknHv0lWRjuYGPH9yPV63kf5I
Il47N0rIRqr4IKTbNPw0w9G2VwbphzsgoLWn66AZYMv+WgTfmAvFi7lTRP4QMOPcOTf1d27QH1BV
iRV5Qs8YR/EiyT/clmzLMBYeC2S+vYB/5HxJ6Fj2klILpWwM9Kgts+bCJOhYN56rwlTAW1+zGZ6n
KtKyn0X5UxCAhQ4IlZoy4qGqkchazgHweCRUqBjxSKpttqn2BnSRi16ROMIwWw/gZjw8627RRuuX
eLkmqAxoEF608QOwGi470XXP8BQm3ewroUtvvV7/Gw7jxsFynfLHC2uoPSG7vXBPryRLcwHKMFL0
Bz/YFRWnfU5S2t8BCMNii3uLbBETSCSoRK91JQ14/Ynkky8xoUL6ZNN0iCxORa/3bbsJ6CsrbSsR
93atcQDjX8vPeQVOmUhyxyPifnGan0tKOH9f7q2ugy7KZhC/u+r8iNs6XyqcSec7HHcbzRjPmKTD
59StIhw2cHDe3IyDBZo8+GLJUU7cozq+R4CZNBQ8Bb95RY3aDg/ruWhA1hlNTVIdkx9gCOya8j8I
VpvajX8Py1wbqP5blzS3lkubcxHuOWOdOJQMk3TIdtd/DzTKGUKWlTCb2lYbg0rJcYqoV/xcfOM7
1QDSpCd0BgPBimHfPvVRytj/5yK9jDgHggE/Hd0yYDKPWZHxMdLTSLRITSbWVMGBZuJSvmxanzJK
DMGAiS2znBv+1k5smX8HIYaQRREDr36YOdVAoxdFxqS72Driwq+aIW1xiAsmdCBCaNK8rkeqqznH
0xs6MRZ9KN5vghQDvhouMDWBhgG7ryKpw3JqDztU7i73E+7puT0g5RhLA2/CPywazGSCtgYEGJpO
TwhJr7mC9ROlzJX4NgS89VuhJO4cetsIdGvklb598RJHAxPCqXVdM5aIsFNP1AaiA0YwQ2W/20Xk
rn7XHqPcpyKBWJ50lXeBZCelrzDAzGq5C8h5YlXjP4OJXNrzCTrhabzQlSAVQCkC5mkhAymd3TVI
Y/ZX4oe2Fn08yZyRgD14zp/33Jr72L+J5mNJnZPeRJTxcBwSn7yKo/dxfRWgf5FH/lebFGjVdDED
xtaXVcUHE/4i90tU+sOx90SA6/1/nZYDcBimIgSG+j4QgqdIkrZJD4UD0W9BhtrOXBP5ySkvKGFe
/U2U+NzeSSV2VaQL2RoJ1yVQemxJRXEv7ejaypfAEurWfVBdIN/gfSItWTdWjQO1p1wHJXVFa9dh
Uh/9w/1fsFT8bPAq5JpfRa//ehluUJgqzUhEtx+pK6bXWhLVeJ/MBfaqeXfBmCEa5xI5DNNYaO0X
5ddkVV6Jbp9ErVkAKOzSJpH80KiAU96EP8Rl85EurPh6CaVOm8DkQfyah2WroPEAH5MRmojjkEEs
69w+rJAsdu/vghAtV/dADUMO+iD0Wamm/HZHIjYNNqnzh6sM2dbEs+5LQpFSrgpRqxYl9uzBfABY
81uuLFjcufaAv+PbQA2zL+qFHT6RQDiceMZB18CtDwJWeRCMYm1SuacLb+YhbK5PXu78mIegwsMH
/uug29hGsXtUWS6L091MZmuKllAI5yu0CfTEr63MwM55/ZW0zURfOBKGFPQ348U0ncUdrhSGtfHw
A9VqnmVwHBuY3ASwFUbkLwt/RFXsNgjbb3CHElwAs7dbflynMYVlyGrr4hKtr8NVAmmhFRIOGAGQ
D00pES9kFKbvxWqb8PgKKUDuHSY9aH6seML85E3hyCX2MbhVjF03Kx6qrnUyAzDknZZx/SMGzyTM
Ejut6xBl+K94gP/JtBfER0jeXrNLfYO3Tg4bcCE77cnq0pVu60NFluzSm33YYiNgySlwurQQ3RC2
gqSEeiCSQszMjEgJaL+AmeJSQQFSUfPbddT3cxXw1qkpHXZCJiR0Bl6j33FLiKjHgw8OgzpcCPtx
C/bMFjl5Ru2Im3F1Bn6jsaKMSIfOPyZFEQzpdnbjcDXVsGO2zjY2Lqc8IX2qCOlQxANOMfTHPMR2
gHl9ZQMfla4obX2xlJ8OWNS+hnJw/eTsov02N+fOmuNYxTcXaf6jAxXH8SZQsNsQDwqtcbqIUHNw
mKW8SfH2EEumKMgwInpGeN7vpkE+ZJ/3RLYiWOd4koIwI07fM/6OleD2tZl+wOtDotTUYHK3gXPc
WceyJ3vZvqdmr/t9Sg4+4ut6BAGwxYEPF+Q6G3fOGDczcDuloHlYpnr6s4K6KgFFxwDO4mtN9QiJ
c95NOwJ8AVfuFcE+x+czO5QuhYUrCoGJATrWGPWrVZY6I4ChtgI64YBF5XTIpZaCYs9nKkw9wWyK
P3C75Ao7eUo/vSN+1m+XyRYe350Pq0cl8Wn2QiAUMIwHDLV2XAlO/telgKEEbbI/oPP5bSqSu6Xf
XtzHY3FXcs4qABFIAGetAaes43mFOuF1eiFgXLOJaOc6fC1xGaEoNYBdL6JsU6grCiTX0zkfScQs
ZtKOFCy60jNpW/rok7KjLNoIdVITVsAMYjPGZkYAJUrHD4CfB9d7lO7avWiuvVg12XcceaiYl7fl
HsUauvW4CsQh+xsorDmheVUJwYWiek5CW/i15HHv2eVr0Xt84dMCeIkAyoTSRFh4IDltamvvUBqF
Mb/ABWhXhYnxw5pzDBWoUYbnOkAAuB45fDvagQzw/8ybtwDI5KBYFux1yNWUla+ZNSb18ye3k10m
lDvgUuL2Uux8Uk7DXPYTUZ07f9hDbkZL7ekbxkD77yl6seVJbMeBuA5wpghuWp+BqPQrONhmGyZl
R9DLqCSwbqGCWGBwNBaDjHIWi/PGoerpMrLtwgS51ntlN8LVqIJQMoydDpm67+yp6pa28X6+4Mea
PP0AiYMRyu5fj4kG4YuuiUjWGU0cTqL1b07XYoGqNoBm+3rZnQtQQGTt/6iKs5+bb4CQlz8j/3yf
BCVjv/GXstoPmEVISatYrFBEcEoYqiAZJNPisUqcJadCxluGpcef/3GHF40ciChEkQo4VApbz2c/
IAEDnGUUwYVObk9DHseC3pMG+fBQ5du27NHe0QFaaf/k9/ZKWgb+E9XmSliTQB1hDG+FN4cebqHp
4oUXf50UyIj3sConu9coE8YLMGl+ELhgQSGghIxibj0legEH5aERi/I/3x5xVI4YEXQF4sD/W4L3
UrEAdmk3oAqD7Et73MsGP4BW+Wmk9PItghu0OXPn+lmbUl6YOoRN2bn/FSnLYT4GlkuAl7hE+JzD
F+afcYXlu/iZIBKabHoBD0ORjUdD+3FofzECVBbBGf2QlBQtTabD81V/Trr1T+dQvBAyypRMusrr
V4QJ6ylZQ5QWNIa4ZsiDPeECogVlC+QLTEVRTeU41R8odoyDpzMc9To5NKjUOOiLYsjdEJhbQKdx
U17c8VP9dwvfcOFCVDexDiBZjcx5SoP0DdUYfjGbIn8YYfmja7vFrf3vtZswkOx6MQOA02k3ETWD
xcs+6wnedRVTP/cp4r/74vweGn60a3eA9NnISzvGtWVO5BYCh7BGc2Wc4QrWAs+aZtakXxzfI+Pt
cpZkuu6wUmfkOq9Yg06yLlQyLn4DEztnrm5Kd0cVmdrTlYj8SL8RKrZzVl2auCKhzQHdv8IG8u0W
49SzPZ67rz9SIG7awc0Xa/WKS4uvp65e5DRJmZAcQzsw3IgTbWPnNap4ZcAyZEz6QcR91I9gPlA0
KQHhHK+dOleCVx5puOZ+Ivg0NdX65e+vCiP6xdtA6zEPDuOJaZx6Bgc+R4aFlM0gkdpjzTROwvQI
0Do34xSWQGilURUrSvSjHi9P8BXKtJo1y1j2X9VBbr8zA/c9Z+Ao9ilz9vZvjMA/aw4+eVwElGH0
rnFSt4Wl84SRY2SauBy77WtzkLDLjoqYCFaz0fKtOMLmZroM8v5ApcoTWVKnFXYDLjQWaW3aI4Bj
Ry5aWNghKrKrW55wDxBaijONM12PQbMol+keCPcHFj8W1s2hO5DwsliAVNoowQcYogCUXa8IGWLN
PRCt1boPCnlzHSKtCTLG30I/yIWHjPNWDwctsOPio7hj7aSzM8O5G07PyBUPb7uDKhpFVzQFv0Ww
zaFZtkC6FvGejKklGrKuhEsZwUo6q22lTRqJZOVDzVUApBbc2vywJfhxlci4Ky6u4gw1gwEvwy2i
CBM/ScthqcaClnvWnwgOXBlgP8++lpG4ruZ9rTHgsUD0dZ/AuTOrLkXkmxK9asUvWGU+fSGsclq+
5wiTrZPT0EIe4/pyRvnU8aJrMoSAFQCQYIV2Kvlx+3a+8LNlX5OUQeu6u6XVkgfjWzE5OGpKGQWq
00uUak9lOUR84LPqCXjaJOhO4GRq5JPaUaJ9W+6zgUSx9HKfMRqjr9vJ0lmLBhGYL2VihPljp1Yr
EGlZOR3hNFwdlcsCPA/YjJMHzTI/su/WCbS/OC22x1SpmKKvb1etLmEbYj5NqL3+OCJm8pW0Z59O
JjZ17Vk3e58CuaIgHsvB+QGUkgZeo7/T3XtO6GL+PPp5txGtXUU2XyrGdu+MpyQsqBuz0zxl1Wi2
2JhHdNizKJWu4j+sMZdJ3xbqULifmfCek1ajDIuAh5pON7HM0yYLkcwG29b2PvEtzJvEpEy0UsPr
3YKZb0wCkU69uVSgMHjjDawa4pP8kXvG3N49bAS+gtxqMf/4oNSRb6ob2S3g1bAPSQoWvR3Z46EB
jqfnWVfOiXf1NDWaQanMN2+sW4LLUKp5ZLi03FEvlSroBwoAZ6WUkCmtdTmkfKw/9rNFcAoLclta
azSNQZpKVjDgyHrf+cYLrOZ7DTQuiououd8GPqb4iA2mZfyENqG2K8MiQeB3Y6cQoe+wld0ispHZ
QaAL1AKaQJvl6iCOSkJgsBQYL1tVZ/YkYp8iI4q/gVi3SS+L/QijI4Nkk9NQuxHjIUJJ4+8009ZA
IH6NgZu0zHqjfD0Vc1yWGRVzC4veK05e1VB1k9ij/MwdOYoWzib7/qDZpAgKI7lmM4l0q+u5BHbt
XsYG12FIEqc5Du4kIv0gj9ruUBbTRWyo3F2rnuQm/jKxoAMMxk5F+UIlpizBoRinz5ee/Zpwq9+O
t61VvMIppQqRddSGg/GT++aNg59UJvV+e+PYnCNFGS3FvsDhOivSe39ZXqrMSTXELA/nQSjIjxCL
+cZ/I+BT+dP5bs6oQjdjEke1IMNIHtjb6kcWo7reiQPQi0qnYVKJmXDZgTB3tyzpBtnoOn6yrPmy
LxEEe1TRsCZBwmjhRCRAmHMNtuoMPZJWU7tiv7/uvBtTMBVhGw5vZZxofilvhohlL8GDJ/9lhiJg
+UxBUkDfWOYQ0sWs9ScJzgPVfRL5uHFU+dVOcZjWfzXtJpLfaRw+05YjnkN763zJxiE4cOd8/giR
cvzDw/ESPq2dR0q6TyV3qScaz2xJUdthndkBN37qDzJsP97ZcOcasM/3vTsY45Elg6InGl9fj0FT
VSoTVkl0P+/yqw4LAyO+HZDaj8dzm+NfgWRxbXDOUcBYOA39rkRBSAw21v7ltE6fx8K8Uu7JtQ6D
z1dKC9FKqyxg5Cntb343bo6CQDg9HweFxWniz32fGbmT5v2FSWgrSDPdS6DEQwMo27E6a/o2JMLg
z4hzR6OGwdwlTKNClq2M4YhAKYsEBdcI4Mxpevx/r42+JmvqKlmNTRBFe0K2E679Rkxf8Vf0qgT6
dXAoWNQmiYy23Hecfn23ZJ4opz/iWY4PghdgzQTEvj+w/tacvvs0yo7sUBKTFMKzJJZx8dlmVmwk
JWIo+hou97dN9OF0p8GTpUMgmRlNRRaoXADBz9lMG9OeTn962orfv4b8jkqcXCN30B/qWUcw8Fxj
HYBrvhH4ANP67/wxd9kbPTNzLqycL464G8fAmg6XMUjy8Czbb8QZDeAZ2NAzZFqKCfeOGRcF45Jh
SawqeJhCuY+vCA06kgKlfFSNJx+jxHbBOq7T8CYiViZL7E4NZwoNPUTuPaBU1uy1gO3HSAAC2dvf
ZJoC25H+r/lm2/x+IhXzeXYA0oCCY9JLj7EGba0Astn8holVSJH1F3JXdBCa5G2Cyi7doqJeWuR0
8S/841ms+qgS8B1mmeOTflD19mkysYsyumYZnM8oolY/WiN08VSi+rCXabcoXSgow+L8z4Pfp4TN
LO7Oz74Ojp/elz0StftFhXRtlXnHCTMQu9hleIPATjeMW/wSEreQR+OCW2ICY94Fgd60zjjgMnND
jkjHYyaEiZvS2JeWoMrSTdA0sOKDt8YLEDY4G2Jx6gNbfF1in0Kwpmeviapozj8qDS5fxJxodv7A
cXbTDPDdBpUAGrC1UxY9ZSp66BI3qKx9gbAV/0cNCo4ixYZ8gNy7B4HJo9EOzBJWzVtOCNFYe08U
E3+Wee+V4Hdac8sjO5Uh47g2gI5icv9jrj4U0uBYSHkaa5g4fUCzPl+LXhy1Ym0Bgdlb+jNe2yHR
669krcAFcbqUVLXsXRP/4RgaIUtiZld55uePwrZJzD1ypCli9gj6G+dSErzDFcKMCd7qufqcICy0
K7La73gIBPZdlkaBcS6EvufS+IjxE6RlX3pumPChKL2ke1R1XsYzIOok1DqnL+JcRdaFVUhQG3gN
fiPfxwGsz7WnWPYuIMrVtiqKW04RpQeDiptd8HTfRVfpkmyizUzll8jMhR+Y4lMA0CaSFqy4ZEkz
AiPdtmhL40hDo50fSAquBoSf0WJQ5/Z/ISt4RmnMX5KsdtOKTl4UxagGPidB3MrsSsPvwDbUvQP+
9IXbl+0MZYACDkLpYAdKAwplvUA6zmYiIYrOJYXCSZjBpfsz8Iunc3jIccakq4XZ/ayocZWgWwSy
H0x1Kf63hWC2YnhnUQ7wneYgpjeuAI/JeHgREY9pIUYYuPGGO6tLYlPDF5b8V9bBKcJJoLsm2BCK
Y/hlltS+f6R0MgDpYHA4E/x12Xs4IhtmiVsOOUw0v7cMPAph9Re48+5dRecSRokOUAhEIqenRuST
Jd4HF3WWCQSnWWr3I24hi6E9MaUVpzirtTOXZ12n8y9LQuWU3JIS1tY+rmf/l+y7zp4NQpP1iYYa
9pPTo0iF6XT9epm5CsHT8CBtUcluSDT+qwq/AbadjZItcC3euWXsFLIvjyZa0WCtSdCpsohPoqcR
LyP+Hm9ugTHKhW8RKL3frJXbNqf9WFIrP7JM91n4DtJZOXDgXW3j+1K+dBY7IthbYxVxnDZqGvhY
CjolMKeYYBPYEEziSuNqGGWwETin5qH2VyEMWH094OWwUhYKS/5gGMx9S9s9ZHCT1tCKZMpKCv8c
fDGfmh4LHFehknKG29iVV870cbSlZaiY2PEBLo90jGItOUVMiKhmSCuv06SX3I4r9aQqjYSCIGN8
nkPWUcXEKx1RHrdMZZM3nTSeBM6oL9gl14kr9nDNjuMOoDjh+R6MgRhYam05mm9cCkVDHbK9Goki
AgULdrstiP2mKMP3+UbAVrs5w7tfkjaqVaBfEXa7EIEQDrp9eNknXX5hq33t6D26hjcgtKUgM4qK
q6/gFVDlo3mbX0pD3/9RsL8v14JpTcPXvgVgSgNxuZs6TuP4fj2ejbqm0oMuBK37UPO1yB0P0AqE
sS2PCO/9USybtl2gw2SkZwhOvEMuetP78harf9X4dW62/yPOAG5X60GTQ5UzqApA19NQIP5cqutg
wTm6JD+R22tACo2ifSnWV3xjPDHpnS25pDukU1uY/lzFDKBJHRVZjZhUQji5lcQhVqtIwJjMLckF
UuNf8JBGVYb17wvX5Y9KR5usHtFxDogz6D79ygLL8cw4xPrjSq0TDHjzxflHRrxMHt02gjwADOGa
NhQrcvTA+Yh89gcEG7zmN4LqzrkeAFwohRCJtgX670pigOLUWFdQwg56+2F99/qbSboX0+rgUPFG
CJPuMavRk5h6KekuEqqkhQaXTgZE1f5uzP+o3TvVDHXHZZJ+lBnkGasJ11W9KTkdgjuPnZBXdQnS
C6aeOJM/CdnimBmOL/B0z2ZOF+PDEjKk/03Q+fVNgI2l9AFHmS+NWmePfIzQ2Xs/C+qxfl+Ao6QF
jcFVquDcc2bTHb61zVKoKZJxkHUxOSDAF1A/79Fhji0Z86EkIcxzFohWqtdCxmZuTIO8ig1sb9/r
xh/G8cDcgAz5zOhaPNf+fTFChBLwoeM6TZHmPVi8WjvWmqVha/h0VEUtrLdr1dnRApbZb9y70y1R
1NUrIot943LVsdrR/4U0n/U6D7J/8fl4GYXVC9hEeaphnplNBl/LuCHxvFRCZNxl1ICVvacu0bSg
DbEdKrDzs2RXuYLtlI3/AIS3qEnlxbR3pbe5DhQOznvmcjk0gG/Oea/HdettiILne7TYj1iqgqfc
321jAzrN2kUKueGtNAzzPB+1ENjNYNmOJMGTHbXr7pv3v/b+48vDaIPcFcy7LYuVo5FeFu12qIIg
+bSxrubgOv63BlDZEjp6NHYjRpKRTwEmEMERw2wlPKc3rYn83tpEVB3seb4tl2pvp0bqASAoSKK5
DWJI4oHJecJSpWFSHpWIIXKo9BHGzHSXViirq3Fg5KGi1CxoXsOk+5JS1UY/GAdags/vvXp6p9/u
Q9rlbpLJcpN3AD/Z7DR9raTp/3kn0Qk1yog8DmOE2FKPMEwmLqR4C+TSTtA1yZ5KLP0oippUmRzv
ngKlyYIhP9BplJ8KuZssXE2dPgvV3xxhtcbhkmoy/zj6pTYO4uq85Jd9aJuuIm0m6qoUqSWmqnBE
kAaRmhlUM9omKTI38IppnDmlANiyzH4Us3FEnr+xNrCrpOa06BtDB6WYAaq2KPVwooN24iuaSAG+
mYs/RSVr+nRyFN/wejOXq8jyO0ceZWmCsjKb2e7aC8ZrhDHliWhKe5kjOCC48Gaq/HPeNpGMo44X
Ay4YJkQLWg5l2G5CGKrpNdWUaQTqEzZBwPWBLfhGKXFTJ6RnPLwdRaZAFzdapg1xhJBtTYCBeFr2
1otSnUvMKmzxUiAU6MaJ9Z9UZmY8Pyeg2Qu9N9YAqCBxi2hT21zd0Rr+FV4jRwFIHRARfh8mxYro
lP7/RHwOknuBtUfa+V44woccFagbyuPGvHl/WP9EXlJT5rCU8T7L/f0BRlDJDZiS/wgPr8hM3PWc
AcCj7PHz7D+jjXLp0R3N1myqIocSOnBlUf5pHzQ2WAlpabJzVJ2tjamMyUNx0su+oof0wSINwHbc
3hCV7ukTUMxowquHov2uWgYDuHqfVT5qJmePvhfXbp8ufWWit0ZG9RX4IA58/RvR0SfrQcjMY5d3
Yx+/UHlWCGqhzPT4CM4o4zjdd+CpG99FB5UwudWJQAjjD9UzmZ9YYaQzWtJOqeaXeOclUTQgMYUK
iwR/If1uoQDXJ9WJJFTDO36KHpNqfU9J5jEAiWA2Ga2AD7zIP4Kmb9eKnPcLkVOwnGREie7L85CS
MXA4+qKa4saNP3SLNrawqD+gq1T0r7oU4CUjH7mXGc5ajlI76nIZZXS2SXk0oVm3UY9w+nc1u1+K
firWm3WFHZ2KF18p3QdGO8RV90SUzRs5wH6vvTEaV1z1jEVD+AlVzUe+mPhKAIHG2ft6/FGyZGNT
kvxIpxzQIcliBMxaT+koSKdTQObfwknv+qn46blmB7GUWLmoy1ZijJjVHqpLnfjoVv10wgJqWLOD
CEh9onctEqZ9SAjxH8BJ3Cj2UlgyMswG03EQb5Ex5KkvUlWk6ytcuTSy79cl7hrrMOHh7vQGpfLT
QNlzHPlp8M2D26FzvWsiKDc5UdSxYLvlu3rfvtZec7L94KN6rXqskE4PL+K44M+J9gdukZDHP++I
3T0k91yt7+L5b2DpEqrLf/HQ/UBqn8weeSqwXYjIAfF8NkWQWkXL8XM417t8hLYUE6eFYQGIqJIl
iI7vgNPEv37qk3aYfMY55pT+NrRY5VPMXV2DWRvwV01iUi8M86xsBqoeM+9RVFyRWYkQiumrlqlR
PpHkaGi0mqGpdA655KcR0uIC7ugjTovHft/ScSRlwMHM7kL8YfCg53xHVDhNInO5GVtXnKOsfvQm
Kd88i9OtyIlacbdBruGR6g2MVhQB84qvXXe918BXU+nrj23QmD4WN1gLWtX86XaaeeJl5cA5SrDE
Vh6JtdsH8qc+Y4P6SeqgDe0+OR8g/YKoQiOQ3R91SgxMAjicYBb58k/Kd82K5GSn4WNBxpnnTxnA
GMeXoxoae1Oq0ZMc6zqPrVXhk42NYv7A0Mmr1IE/45RL/RvRUk7y6438b+TLoU+HjXHZbksK8JUt
M06TrKYCtmSlXIloUd/SwXG2So++a65/oG5unrtit5R58h4f3V68ZGuR6MOc3LvhbcWuZirAs+Mu
kfNVtkC7VJ+39AGFV+WO025t0Si6Oy7sdZnXi2n7+E/mEkUcC6/QmCJQ/6mmNsp+r9JfZD1+fc11
951Sc0k3ZhZxOHZfMFdx4jJX7ZTma3/TWMuWSHNdbiTDV+qChhj8zzt9CbpFZYb1pa85BiaBlqii
tQEzDZ3jMdWGMzmDxCehL4blBjRw+rKPeF5GlCG9MdmKqRDYk+rRGbwqNacCVbfPuBKnhuJfNk5C
KmP9OFnWYmvene5PKgiC1jxjQ4HOZ5wxO9RrHkGGu+A1JxiKiisahNc9wmn7tw4TR1mcrRE+u9Wb
V3dRMUqxdOWubEnUgYcYZAcAMQOZaqHslCuul4rBAtPG7xmABSf1Q6W+bvc1hIzEDLx3cAJJ2PNX
SzgklNQ8TcS2Hwxo30S/OZw2yGhASBw2JsoeT2k5CKJNWP6CNCodwLcRPe2eHC06HapSetS0fTIT
bRUJgLBkoAYDGX6H2evHIORUrXp3LcLkYdCKkrXQ6T1MkNsAjsjwu1obD2IVd3THgbMTfN38G2jG
dQd2S1qzR64ZXa3Jwg2Yk+odw6TsjQ+fJH6WhnVpfPpfauS1vxgslF4Y6I2XuDkri/45g5KD46/I
I/JDZgx5TSwNlqsxRgSW/7Zfxx7qOAm9cX2mbzVth+xHaj2tVujid4G67Re2bDf4niXNfEXiXLsg
geCTQHcVuWpEqEcQmPivK8agiKNoWabm8ZR58eTcc3aBJ4/KwSWcyFqdYRBmU2ZIqviV4gutUY9u
NIhiLDbvO2fWYpb2BhSyqGNckl/moZJhAfXU9dQR5IyoGRhOLyft36gm526jtAhRP3Pqb6P21GKS
aWlc/eh/MOc8ubrhC5q5HCHzrB3At+dROxsIQLHy6afxdsi4HRidSDywbN1NTC2Dw5UB+9LXJG6i
EnxTAjIsJXEop2clR6/YbFgOrdZcr3UmG8+xvv44GBJINT6LIe+7AJEclnWSbzZuf82TX1GYjvvE
69V8ZFJdtcoQv9eoa10c07ldSiBGZhz5QIF1b2NcORrrGLwUmWQM/afNCSDWayl55KHpdKJ2Cu6F
HhtSTZDMTJ9PHqZ1kQ2VJzCzhoJwh1+SWy5OQdXNKQf3EnFPdiikLoloCXm4K1cGRvUXjcB7jek8
8ag1JjMOdI+a+d+VKY3pInM+gstwd9fx2nnATPHIQJcHtYGrRN5k0mUw5uOkikVcwX6+jqgBE3C9
OIgd8eU//YvfYNESBKM6a1EVv8+aRKLm8zHe7Ph7dAYYn1Tro3hr4xp7z8M4zfOfDrOGcjx3fJLN
FrHILjOFpmWL3yFLsfXK3tKCmMwVDezYmjeHXkff2I33DdNoE4JDOyOnvON1Q3VTcI+FMf3tSiqA
X/paagEmBI9mQoLtWxhFYcRAAO4CmJH0YQ8p7VGkE2A7Z6JZwJjm3BV1M+0V9p6ihPSmkOiYvdy2
9b1NpBSdXse6h80eX3kePholIudrDT7IWrMIie96hcvY9DIZkDgNVTRy6SY0JOgq6SSdHRY0yHOr
St/UOnMfYXPEYVqVLhwRiW48aZO6XdyN5XZm3ldPRPW4RADPcrYomsyfuZkCMCcbccJ74Kurk5fN
O+Y09vmKHkkj55kZhgjrJXXzXFFG4oU1psEfrlHeYuuLQ2FGPevpUm+B5r6B/eF4828g/Pv7zcMV
8fR7AtCYDQQUxBSxTg2bELTWaYg80UYMCMDTF31va69b4x0e8VOQjF8arW+Wn3rsyy5VbMgEyrPb
kag3ItfdVq2CTKIgCB1odQHDMGlzhNdeaazBOYYqFKD8A0Ej4zGCMcWKw8Cs9ULYJ2B+nozNbRe+
aC0WNYKQFAB9RWLSRVyTyqRlve/IKTMtByWeUKevbrBjbQ0qgEv8pFnu0lkPgJXNWaScORAqTb/Z
+hq1P1noDSFaDMQtt2KLKNjtm6/sYc59HYnmPhhtgwi0O4LMU7bwCE9kbWrJN5uNB/SdaM+BlUMw
nvKm/X6Q17Y0vXCco2Ht0FxLwxzgqEibewQYVI4/Hp58g97NvIti6znMUWdDTOi9FZEF+T4NRrwU
r+z9RBrTBKBObuSq+l1rpCM7y/KFuIOl2L3qMKwrh+r8MPcPy2VYzL3q8Q1+mDQ4D9F0Ah6rl0dC
J1aEDzrU/4qMRJd86UduaqPG2i134YuYH2mRMXWFPjZxvmSRn0QvjmgRvNdTwrmMRKtc1G/rFNYY
4n41swhfzYV0wEqZHGCPIrfPzZJI/Wf3C2fZEFZilJ5UzCCs1wuJ2DwcWCpybrfOVgtPvxfXcX5g
sZPULmPOHczeocaxiKJQ87w7+iTWwmohLu1ra1nD3Z71/1Ux3Y5/Z4MGtXHrnVuSnSnrwwHU5Yxy
sbaTSq6v5M3JCOe4OGLEVNCN96Qz2UV8wu0e8/Yz7Nxqb9YPGjo5iQ4tphkPUxdHBQtsufuQHa8i
jDZoq+z14DA9eccOSB2nbQ86koTxVlZYTtv8NYTVY/aI2umCX26uOuJEfFLOA4Dbzlg3IokEU6AU
GNOh9ojDiEPx3xP1rnHlPiC3P+wBryQQAxq3zMfJmh3kJJ+q1lMhvGYmJYPWDnywjgqjyY01XxcX
rdq8kGf5lU1mxTmj+KArpADjq4I7JrTPsgQWZsdpfRQN4Np74UkXCAttNF3eDNMyl/kK08vSWEKN
W2qA2Vf+rOVeHbn9nWMgHxkNeQPPJg3hNfvvkvCYHj2UsJbJ7UhQrKc1kG8mNx/7I0XdxACK2YQ+
1AUviXbpGck8sJ5N873pIJqT2taQU8AMpN/weZPSQR86KI/rKc503G89wRWE6eGSXoln7rCeYNLH
4v1L5KGpvP5UL5mJ/BG5weM8s7QQ0aBk4aiKkK8hUHiBfuyc5gVc2LI2q2R3wTGK/Af9hedVRnXG
pDS0n+V+rrBNrEC/8iRs5863w4FfP6cZxzjWQ+AROep2Rw1yaJjIhJSYMXtZzIMV/aamAdcNdGC+
3W50IoFCUjUj90OblH+vJ1TcGe4hM2dyF23MDhcUrS5cLod4+s+IcLsOgITuzajTgJdth529f5ek
7QSccIPCuBJ5gfB+XtkH2pX/WWj8u/33ePBzpkXfNMfNq+rJWbjzazFMBB66tQxyZsLbNDyKwRix
Wsj5o05PbcUWt5zAG9+NCZFbUpG8MJi7xW7jaADEeveuBJ9+WzOV5h7qh9LBP+xw+LQYQFp6u9PT
n/vmLSbXQW8SyyTWbplWxICkDAHMTc7ctme5FfhozT8JJMT096BCEgLK3eY+AvO4UhF/RXSqX8iS
Xlt6FHTWGR5bCrh73dcpx/DrJtT+SqiIQeKdJgZpQVdiaomt3X9fVvgCQNcAhunz+E/cwwwTLtS9
7/Uu7CYAwGm+fgUv0dR0TVgk9Dt4tXyt3SgkTWhDytWn6mJ1SsuE7lxNW1TDTItXDcHwNA/6ACxP
Y/XqWVvlmIh7ex/yx+tUvQ0FBE5fzV8xlafShwR7tpA3maM2coHcY9j7kfmVH9NcFHNlJfH7OA2k
/C07nTDukpx4UWD2C1kNSivEwar++EApgLzjcnKQady8V4ozrY/J6F0bze+k13en3sT1l6vEUOki
4lcWzW6v9ummD63g+OSpoNbsZ+Us1zNZ3TnZAl4dKMMBsX3UHihHAsxgowD8C8670gIO8YyULpHj
3A2Qa+QQgc9Z22humVgChKe+wOQBBcAxxfwX9ozGQV5297vHKwEW5+4ZxvKA6ntei1DGELDgA+5k
hEu6wvu1Y/lBwT/IjS86jBrK6ytPPc7Ev0B0lhet3vpWFmfdJhheFuF02nRJ5GhIGFAQwTwx96EW
7FhlfysJCHGjKKuE0EdLbD1SpK2CW1r8LyNhHoMTYO5Rz1UN4xh4Gbc7OSFC3RzEHTwZiAcUNh53
3OYrSBU+7X3eK3QSudYNmDR82HfDlCN6EJ1VyRn0+C5LWyUV/5A8SE9FmIjr28gZHDwTCKzcgvzb
bAYRx714pZ4W6aacNs8DtOV0r/o8PIAbEtJn6h7CWwHTAG49Bn1Il1Wd9K8np+SujnAg2du31pkU
iAIeFcSGVJGvy7lXV20x+D/2hU9QM/R3y/1NXpYyRkTUr2mBsx0OkXJjfapb/365dsYtyFhS7kxQ
KMKWWRukI7QOZ9O59ofFZvDasqiHwpiyWb1gLZVDoVTsAUpOMosLSjF/hDzrubRDc2tySnKVse6a
IW1u1iKR9/YXH0xUfJn07COWfacA0ZREaNKJ+y7tfopGsGLZzaoI89X/vpoq6hyk4RfCcKydctu1
gL0maAqkvhs8ZBFGgK3PMeNrfZYKb2APtFAqAbgdVyu6bruTo1k42Q6gehjXQUKaGFjwNaUKc40G
4MAXUFeOScw1movTiMBP4xFspnnV2mH/MBuwmlJdR7vRqSG9ci1A0InflL9DNC9Otk5X+ys2nved
jnOfD91QGwcG2tT2UTL3Y1r9LXSpr+ttjp2zsrV3NhlqtRbcChsqZKQoehXJ6dbgtc7mHHLCBd9j
0WAN+H6GCDqs6Zk/nQBFtwVuAm2n6mFESgSeK7bRakcjdcuV4u+SKA1lf9cdWGU2ttdK7uGGutBI
NeCJ0szeGh9prLc6qBRafDcgId1JalNTkolkHtXl0FC1k3F7qNCTummQLMslQOlQhbWz2bVjqu5j
24i+4jqnvnj2SeCFgGM9W9CaNOLKqqQ36MjWORfRtrtL7oi7i1dlLaDDpj1ow5AE6x4no2+yJufv
K376PwVd3eq1bW5yqSODE1ds+G+NHc7M4qkA1eqTiZNa+SEICx9fryjpZUnwXNFXy3nGdtSlyJKS
SfyT+SQB0fWcDjCvyrNzk48XlZuYl9mnFFmkRSGutH8bXp3+tpxMbju+QElJ4UnJDZxwlksFjBwK
eGQvbGdvLueWPSM27BI0yMAd7OULO+h6+M4djUbTY9iHbr9qGQrnTa+WrMs/knQdBOn1cnCgZNWw
bKIVqDZMxU8iCm6saysjc+vfwGOk9MDrYhNn4iu4WoHqAIH6mHGRSI2WBaa+DCJMP1xm+H8J6LuV
Z1pWWHIuCy/uSbWdmP1Z5EG6zKSII9vgEbC24c3Mu8PGL5YM5gNYHrv867dpsXjYLYrTQfeZEd8w
pnHmB5il+AJK/ThE3Cs7eRe5ykf7wf56sewJcFbM/opob43H8ZHuai/k0WJ7TM7IG0QtFizhThvH
4OJ/N2qfG/PPlkcsa0hwBHDbR68mLvuwAZKwUU55qfV04dUOLKDUSPYUeJKISs4wMbz1dqLaW1Qc
YIyacF7vYUeDN+M89XLo0QpfVYtkXRt6uJYLTQ6uCyQ1NLhXN4jO+ng/JNJV/V3YD0+H+E8sLlgr
gMz5TjSXS+sD6xBHDPf60eExL7prrVS5jnV+bVG3ClXYjA0idlWW/OgNIjuS+VIeSTq6ekIWsa9l
ajHONpJQpeBg61aVCr3+NLgUSkU3ihTpMRsh5Vs4VFyzJ4iCJtGmPt5HUB3Bug1j40zWUKTvPlmH
crvqEws5TRftE9YaICnaZliINc4+UCPevlP7kXXPy8Uezw262dWv7SjB1rovjpjSr/v+Nka/LwVN
MtB4ceW1+xumGcEuKt13rdQv4KygM4cY7RwmWZepG0UfPq9SvQTjz/EEQBhDM2mWpZ2h1dULeSIR
nhuu5UlUak1IdZMrxLO2tVzP/9V9rXOzyB3IOvpu0up0rVYg+9tddXhItOigJIwv51oTU73TyOG5
nXxgiNLnETsDSXUYXAMx0WYBFbOorru29QtuuTqEoTaOQNWRfm69fcS0UrnQMLOypEHz/1+bYpMC
bOd9ezGheHCVgkjVIfOEZLpNyl1v0AR5XSzC3X9Tsk1NR+iHXF5fjPegp0f2WHZaJW15Hrhlsr+t
R9ie5t4lfdiXoGCMm31lYPjxfR9J9vtONyU4yDnwERjy0fooCTxEyneMRWqReXBIk/GtyAYLAt8b
InTTMaiMC36Ly3RYUIfz9omHTR1Lug5EIoSSvERLHKkh5yfwtknkeEKh8k+xi7Mgge0ILJPomewk
rJLaj3URt5xVor26URVtCaeCU2RxBTJp8gqLF/PNTxuJSuLpslab7+YeGGkNtszFlRpYecgWmXNo
bvXQgDgkFV8VmVlJgE0w5AiBauevq775Sl7lW2C3yIfi5CsW1qomFyhVJ9CRjB64hSNHaXdZNkEy
VAQ8qmmUDCzMIHdsylmDozqirQ3/WJXoYZeulVaGO10iwjmApX/XVREAhjtS9lLAj8ZBo6/2CSH4
ir8xV1f49f59F9bNWdlnjWvgAjFvnhO9QiNx9CUMXOUxWwe3vnBfRzkmm9X+AYawbuC8SOzZZE2v
5P3tujyByAhyDPnBdK/qeXNuOk5lx7Zage86jh113ffFq8Wa9e/FKNQjVgv2I6Iel4rXuwoEKrDh
3scL/FvqEtY1e/EDYWlvyXTf0dlgvicmRZrS3foJOMqx7f8P1lnLk6L40GAkUQwyDzUd9RC7yiwD
N0TzcRveY1w5YgdFgy5HsrGztXi4zLE+gsUVrnguH78CtUaOxRNs60QSzgK369cT2S1HhmQeiQgy
lmTiFYIXfRgtTxcmpcjv+eKXs7C2qaaWHyHc3JtgdTWk1aPborRcpn1w0vyM/vK1PQOw6gnkvFwC
O8HxaKjlZ4/Zc0Zrwh6mmeHnfafsXoOzyDAGKlnBiVMx16KOBoy5g45Uj1awBP6/cboiFjxisaqQ
frZIyIlAnO473WUJynaP+WgVWjcYx1xLUKHIvSws6MrpBqLoMpXWjcigZMaZzLBuJlJty5bk3LMf
5b6gxtKOcBOHIDiSlmThSad5tsiSI098py/9FeW9IDQamcnU/sYiSPo2rzbMefx6RcToMinBZZqe
229uL0ARYwEKKcO5/JBWjMr52afObpc8/HKVkDZ/1KzcAjMoCNTDlQQKNpHFrU3+3wrCUJlK1Syg
nnyep2Rzm5Jd8h8vlWQWrnRsZ1ZjY9tD10paaTWmjy88euOMFsSYm6LKQbfK5zdE42QSxPTg63Hk
0Lje5+VjLy+HcQPUXAldu/PAodgZ5Vhpory0mhNVUMBs3mENCz6aCtPUlgzVItW9ELjRGn9RrbDu
mV1GXaeiWEEM5+n4jEmit4SpsHK7nR0Rq5DSfgctkk0GXEAtZw4JwqY/loUIounTYMjH05i4dS9U
rW/R1NizMtDs6Ep3wu54Rl6qGXupjwrlCOgnquSEp08MVIo1cO18TaZxZ8+CdL4JPtggWaejBMfQ
esWML7srHEsnJb1H5qVWeib37LraF7Z/RHY9tw7/7NdPjRpw0rO9E4Y18lOOCZO8dH5kp8+KV8hY
fNC1Tq4neKVqI5n4s/VU+UEjevCYSGnobFr/o9BoAdgsUyYTjbvHTairSpnnRWyd48urdq6brXzj
oK9DG6qECSssFYagqvfzA1gdJX6L08bSyqMgM+MMN5r7OOurLbGC/0emhjjNP/cmfcQws7iclfld
bVjkcCXE9sahleq+VXpEdCEM83JKP5c/UC++fhS8LTpNc+DXVb/lwY/pGjxxiyeOxNb0q89lp7tD
PtXZpZ7hBQRYa+WBL6FpAPkp+NUavHmNjRNgw1z9JGPiy41KZON8ptuYX2Xgf05rUxOLTQQdUAPU
/p1ELKlLx3AppMWsfdM6P5iPhZVXeJ6TQdeuowQlNObkJ2s5sxn7axjIPrNonm1O2j0lMUWAaCRK
ikannakpKJK5RYOnpDDV5BRfm5YChX5DJyRCpbZ8FrkFBqICY1qPlI/Uhnx7srl/N/seAXyNQwht
Ttum+rYbGAitckxtd+EicmFtR+wNR1oxc7cFrBESy8duCMIsDpV++in4GJc2HGaC2UJMKYBNO0ZB
vi9TXUDVaBhNB9JLq8fyw5fet0sGLTVv101vdtkFU5BIx+CYxXu9i/WZkxBoOt0dOUFqOfLVubzm
LuYR+YI4xom2HCCC0HTNppS+M2vswZ4Loq2/c2gVx9GCOb5xEHMAz2rMrkuOxwcTkUGucxhaxm6q
KjAa9XeyJ2byxRPPgsShJdYw5c1TJPOivCBYQJsgT560cyia7jGlNIoPyJA7DP4qWqu2cVA4Oar2
9seE/PE37pbjcHwT8hQDkXJvh+GJr4PcdhbW44QOJGOD6HrobqHKWvzfTg6ccuNqZpoMxvuL4SYU
sFIZwbxmitc0Up13jK9w4xpMeD5OAZJ5HO2PlTtflDOrHu6/zyIIo4vzWYq1Dvrp+0W5VIeG5WPf
p0Y2i3zFwocwrcItd0svUdGzolou9JLECYo3lKsg799JcDJNXWC+hhsdjwUDfojbTpsVwrdZM57V
C7ss5GEy7x/BHRX6bmGTzPXxpjJKsPzC8qacrRRmidOdabIsQ8bn2DExPxkEzAiOTnKGgCPm0llx
V+qRCEX2Gsd7eWbpVDcvV+Wao0WkOF09X4OIkWO0ey3yVtVvKlp0RqbtLEq0rfQ2+WO5n3b9c3R2
UfEp7T6hgF/Njssk/QA+6gL+5ICWm5fwNAo/e+uhqo5QFRDscB/NNHTZ7yOnpJDq6eYklXo3DxOt
uSypU8S34VrYDnWGthXm0Cr6CjhS8h5TVWEBcj3nDysatJMrvV7MbjjrDoZOvmqyOyQHSvNRZEl+
NPaP/Tz9vOScM6TFb/TeHv/FGSHdUABEiIMUyCcwqPe9qt8RvLvV9qMB74Za3mSSMxpRV4euVjJl
JriE2llIzfErmbBUQnGPh5w6fLurMYU7i5Gw6G7ph9jlnpE6kDk75YzEYTkiKY3cShr1qtrfHjDa
yfdfoRRymRVQWPGxcjpjOe8N3YWJ3uNQuArdF7eBP/pGYKo1sdw6INnu+Xb24V1z9eDbRdeXFNdf
KBK+qLqXXwAkCyRDUNauu1SyyVCkMo0auYTVfG7LeTL4d2TXale8wXjOhsGLT3K6H/YMx+ey/XiL
lz/2pFaNR3nAed3HV3z1hsSdGxFfFAp2YVt8khAOgV0EtAnvhC4aVYYtrqY4gK/Uxhq31UNchXgR
PpLBy1lhMIlSoIQGgauqgOazYdFQ4CgvNcwyQ2xEO8hHi8LUnqWBkglFmR7fWmQKlvEl7o9ZHf1Z
7Z2qyI0ORfbY+iuPMf0aQKfZpXroQC2cIEiApjPc5rhgELREeLyOEFFxzh+zzslFvKstaUcbSLY4
NeFQhEvGtQpWv0nQEzx6NRMAlUXcIxZNlLM71dObO2UdI6Ro8l4MTgGjNMSgotL8czGGkCNe2VJq
wIipzBpV42koQUHzvKdmQnzKcsFUoVDBWZW5L/ikLrv9Rtspf8NQqmQ52s8Cdb3GzmZnmANFupB1
iWcUAMESCMiXqRbxo2MX01u4m5ROBf6lHdB4lF5mVC9WdMr8vswyjNHPBJX4ONDiP9qOr/AXbki4
XfoEDf9GRXAt0n+fhkQ+TcMItCF/44eIJxVcxjp8xhEV3Lw6EIY5Tg1dt4G7ESRy3ZXlaR9xr9KV
1Fa51lxsNva9+utijnulEq5kAtGjf6aSua8NL3m3GNf87XKLSxy6VOjPP2JcAy3FlnW5wMWgCY0O
iEAMZz1MaL5mG2jLj6r0uJXLFjHK8ly7WimqBsWDSdmHt40G0uGDbSHLqdmG0I4fY2rTwdxcRhmX
4GYdbpplv2KZrJQjU+4FOwcf+w6Zlb60RNwFYIn96NBisG/q71Jy9Svzfhege6JMUkczA/SvZ2Yb
6Ynuzy2v58hAUqK1FR1V3fspN8xYGBnrUbPUUajz3qoGFiTQ9gaqAqxcJgQqiXC8hwb+/Nfa/mox
BpLDi8sJqciN/nJi4QP3K2SqTe5WM9U9QIyQ3U93SISl3CdJgpc7l7Bwch4tIN34XcFN8XNC+HTr
eCU36hIt6bz5qkN6+b/gGM59+3C4Re4065u5zogpXmMryEB+20tGDyjrM6bFiqbn4KENQedREXSo
MsVNPT8LKWof9lajNz+wq7uhuZ1QtI5otLlpkw322CwP74PN/mdP3pAAeiqgI+BudUUAogSLG2O5
Dt75IZoBD/QzPASGfAuGX3nkSRi58ZsF5yKABZUG/M4zs55qiiGZKciWePhZIGUghyX3nkQn0JY3
slD2dAuDUJgkiVBGv1Gm67LjqXCcSnpVcDv3xfl8DloCrwxxIGyGljdnaD9gQk4QDIboskgMnjNv
XJ+SdKV4pEdhROTkpUOP45JtulFXhRRjFp0TAlrHknpIBe3fBNQhiMM+xr9prjuH2ZY3rxjbUsct
9rE2N674OzkA5ZSKsbCLYmyWPhi8Ebg/YxsN60BxL3roCieOKjmHqD+NkAHIOWUHq7aGQ82V/qTt
D6clDoWarH0ACLSDn90AN9BHlRs4E/rwwa3Qxm/jzKEwoTv50+cp7sAEroLFq6hIdzFBnjG6+mBJ
NJ/Zr/T4ORYFkAnBE23GvJ/qeywP8GCHdhx+PXoTOPIaz0RoqFiuygqIIrO9gA/XtKlxWT7JK1XX
PijSemO7joIHZlTIu70SYML/u+OP6Dm1oVwosIbv+Nc5UYaTXGfqxOT8Co89p2K0u0bZS6wxwPGv
vqPGNL4V4qRThAvWWAUnoEJZELrxtRqtPcox4Ihaxca9q5GWZSDjaOsdjzCVLfyKImNbznUzCAcH
8MIpEX4sCaSZ807w+tapBKnRh2v9wSI5Uqzbij/VmhWs39c42EiFGNS40YeZBstRplRPizRAaSpD
Tc0s5UK99PGZ29TBgOcs+cpxcaE/Oo8tK5fiHI3SO7ul2taI/oG/2VIEBmR3KOsPiNhyqRnMKxM7
uJeMTxBiwk5Z2dWKhhSVB2Aufiv/4Pest+xexYBxLa67aK9lVMfBjmHCapdFPyhUs0PWfkzE9JA2
m+uGlDqdOwwseO/7fWDQi9hl4l2yD58Vq1idarMzrJ991uDWg5VlKFaZGNGbLEkKg6SV19XsVx5J
g9oI/HqtbjqKbG6ggSchWmaDEmlqFhXFFXcZmOmscc99dX6DFutrOYnw+23oHauxEE8UUppErhjB
ZbXqzPQJez5afemMQKn0Wk36bBpejlsGuWPw5THStOI1+9YXYsnIPOp5xFspDpw50W69TQcpGqiF
XOHS7CY2lJq4EQbQinj7rE3MjAhrzVWd9A/njNqrIsXVrmQDpLKOpk+fR/6da2U7k7E7pNQdMef8
I5ikOLhODHFt4uZneb/FnsJTQywzRoJPpkKE8lvcwSTimunzbFn149vJx6VoRAl+NoTcpu78DN+L
Sb2XUWpQJoqlzohbG8KrgfDR8FfcGUQiyS0jJF0ocm6faq9DNVy7xkG6+eg3wma7DICdgN/qaRqE
EIDN0O0MqAk738xhuHOWo2opIOlt6+dFijFE9mEwU10f4XGVBvs6+47q54kKjqGtx85NTNyAumZi
4WHUoErY+A+X7V5NJxpaigrecl4iB1jRHUHfQSIJe0gdqYFt/9rrv2XqgiQ0tgBLTS0PJ92GApnR
xFuvGnpLC0qUYHPbvsEz2cYAMiz6cHfovGisW+a09Dt11tG7jBRrBEO72GI2EBQ8a68q1VPjtm5s
v286PSFv9j2Y60vGNkgrEQXC7Y+G0iKZx+wiSd2+bulow41uwDnuAzN3k9Zp0ZuG4B0zgg+8S+i2
HyTMRp+5RFcHpQsFl0RihVYMb3IZILTh84dQUTrmFSjQIRhBl+swEKM8dWXWzWRfMV8P5TZi3ywy
CsD14PFnGNru7kc3C+x02/YYexwxVxSe9ioIQ1Y3SKOv/sYGeOFoNqYjaOsNhr+eipEYsDqqqveA
/IaccqAbkVzXvCc33oZCxOTz+E0sj+ytOMA8HzUORp+TwmpuXX7s9ypGD6vtunbyB7nrUFfSCETp
R86svNDAqzuaSgqAQp5CULKh4Si7bMK0/sX4mdG2sAYVnbxPfpNaILv8mFtMBCPfyNea8yTxAO1D
OuMPUFQrMrfSQukff91uz7fLFcga7VqJ15xiX1JaFICu5UMIdgvACciINB/mpUsMKiqcntBZ9qOq
v+ovXm6e8OKIPBlLDScL3gDlMDXSrWBbZF4Lcls2QERzi6ovdCQm58YY5MNSGde9b7gx3kVTSWzf
TlZK+hzC43iEC2wtvdj8c46+CmV7D4bYewejVdT92ejMTaE+xnj3oMrI0a1Srp6uxouai4qyUE6m
ucDJjsRQGjR+Rwiil3kh7iZFXuJs1R0/gTU/j4jdiHoV2jPaZ2qevzGBioY4MF6TPqlgtq9PNYhA
sAiOAKsm90DyBJaiOUHsR2QFuS3TVgLWr9LXgxy/5py+FvqJJbJC2inJpmRFBzvseNNrlkkV0iLg
EOy/D/VggolyH4vmQYttVJ4HC0Q+1dRONS9Rex1xuSzdxMYFD1BXqfAUkyDHPNxHxiVVOx+xh0Eh
IILOlT+pHGv8ikEH87m0EIV8BtJmxirRHFRCXX2coqZDU7MQGkz7L1RrFxCzsTkT97On2a6iNxYu
A0qVTb9mcL87D9KaxXsVDXVo0/rdWiBmq+hxsqIHteIiD+QGsBujPbXjHfGh3SJNp2rlFq10/c8q
yZwyqDR5tC2jdzc4F3+kPE+LYgvK7tEiFy2Uylels5GIU2holBXuHi+do58DFSjDYA/OkIzIhjG3
8NEPLacnisz58FYaxr4rCk+d2vITNrep95HfVmb9rDtWuM30wAZqIllZgE3S5njbol98oUQ6ZYKG
M/Up0yiwNCzKawa7BPvZoOujf7lroSpAO1H23m/A88wOdXByKB9Cnj4z6vNt5dyukDvG6NVl8Uqv
/LKuJzc1jjRz3c+VAKxNZsGoLwizf8sxbskzHio061YwtMfqx+jDtlK6nw+cMcEfnrE/m+xEumU9
nz8nA7xPXvZ8wkMnI12Pd8vpSx4RFNjjBOxBLbCQZKJCjCq0a37A69suEy7ZsxjYi8ZX4ES4b6jL
NjlsIGGeCT+dAHWn6yJuJbohyjom2u2jobWcakcibcrjMzc0EDYscSsoo/4HJrWuip7PzukWjWva
UCmR72cHcjTJJxmyHHtE/CJZxwimDuWHztap58vHAgA58QMW/jPtXMwYpqrJZWAL+yxlI/vuYbDv
kMH7uzx5inIFAFbV9eDSDxIMNzp3mNuVwO1Iyr+RXbIaHBlWbFCMcl/9AcfF1Cy031gaqM3oHiBx
cTa9IyNg+S1jtmeAc74GJAq6H0CpxwZ8CBQAGe52KKe0aOcTwMoaCwPjNdDYNv+DRoHDrsWCXiqR
mUsqsp2lm9FqxTYGYtQ2nTiWW8QSkpy8Rmmqbes3EnMAQEAhO7lZ2KpELdaeFv2AQQBVaLTPttFO
WMVbwrASbvDQkCFXAKmDwXtrwcxrjInR0XQAjbkaawnieraRzRQbjd/akqQ6zYwDwFi994PkQLaI
7+DLWKbxqBPZw53zyRIRIkSFDZnT0+9DqM0HC4ITcnYq0XsDpc+rMKxOn48Qe+Kpx8R2OpU9EepJ
1fO1Q+4V6/fmCxVKXnZU/SuVybz82TV+NReR6HS7yDLYJD7fq5GOQfNg8hbubQua9+N93CESIDo4
1MForNmWQP53ltgHcOZp4dOlHyMsJM+NBR4nhnU6BEa9RCV93th8nPzuN1VDK5L8X1bOVkVkmoHS
FRRarvFX7IUbwQEqz2lCcO01JAdV45pr4YYy6WV7o+DjcjTki3hcZWadd1+L7k2xizy34bCvy2t9
mabg+vr7ldN8iUnVMIuEApnKBO5biA/ty4O3X/+nSgtvxxWF1hwj9oEkqVXzf523in6vGEMp7I9a
5Kq3IZUmVQ7aivhA1MYLofvrlH6F2pYCXhrFhwEtR00u7M3nIPugoX2SSIXJ8UJzcGsfWi2em4YO
INpP0MLimC2sAtYSSJ+aoSiKv6Hk3QWL27k+vZfRqR09sje0/PwO2OMc6E7KrtzVBgYugWfO/dJH
SlSan7IgdPCrLObAFltIvQCNPEs8aR5v66+yj6Tp/g6KDrVkTLuNiVtkkhtadv+U2/Tom+849AJ+
G7O5Qvc221o8F5dDYHsTiFtM4ParU5r/zKgceOCPzHzt91K6JqVlnCBLx/OzNRIUB78GFs2H7vFf
Slfx08YfX3cYGrj2O0KricPtmCesOTHvuRPRgGAOhDF0nJkliujSsZ+8MW/P5tSZnnq1Gm7btSl8
BHB+IQ0kbKZjzasxlBCByyZSREld/he6G6kqXyVgYtUKjeKQZhVedyrkcZjuIEXfEDtw1gFEQiwQ
hh94njd5aGwQEU228DxqPrV7n3+ZZtKso1puHEqVDlQRG2+alfNRjxeDmtF2FrfIKrP3tKBm0BQS
2A4xoq7lq5IBUYoeVRn5WWXd5JWjigYmCv3I4yraHBUPcUV7a6lYkC4odWbAmGeUSSFWqXmGhX8t
UshqmHKwGzg32oE48uiMagkN6z1SFX2j+oa12tAsLiwIiKAO7kThbxwOnANJ/aoYiahtvx9LD8mW
dFsjji9tFuc9BUBpImg79g3WvcUTPNZIostBvx1YYdWduAN7+Q7rf3TbdIieL2HPYFBJRyYoXaX8
9nYWum3cN949jPj+bdE5K2NvozQoeed5IicxW2iaKBmKtH4oe8V14KOsyLZMxjlLWhBZcS0D1mUm
dr91X5iTy4mkFw0sXmvj9URU5gRizrAuK2Xqv9qZEgjJDjqWKZ1bZFD9b0W7ytFDWRQTx+kzwB8E
ELxaZriie/JfJ+fEq3+pIpNVK4jemG6SSaD5R+g6ST16KIK6+OEli6DB/M040aMCN/z30Dmd2HLV
r4LLtvYyYRYVw0dfh/xo8qJX4KVO+nHuJ8K6iUrl6OQ7cOPMb+a855r6xy4GSAty/rYnTPV7h4RN
dGjRO0ekyL9tAOeTbx/ETjyApIOOSrK6eVIMOxh2Xx8b+WxvK3Tu3YdE0jTQtq8oXX1/Q6OueTlL
axIQgncPgAQTECgm/ppfcIdpHxRN8BMjgF8VutDFwRqUFPzgXDwAuIH8akL7p5obAawEbaFc3lCo
K1zLXe7n50OLwN82i0jqjSe8q15JB/jixQwVI3fqWG2RKKw1tKbMZJp+mhjFWtq4jr/STOVEd4SN
JsX9whE+H6CRqe7ceItV/Yte3CgAqQgg+0cpIR6WABP2OFN7BW13QDOREGXa3fIH3GFDR7VQ2a4M
ZxBRpBC5qJ36DCN7PcJWQArb+CzW1T2FtKIDCw+uuFLiYwmjqFCty8exfX1q+k+L/5UfWgbS4QrD
ZxpwfEJzhoF+P0Hum8f47idvkWUUAaluwb2jGHjIXlIbK/3zN6eYF0e7OA4LCKgKVMIcEZYlytI8
3dS387B/t1syrVY34NySnkZxDnVR4P5smkjWFTKnTuD3hfND5Yl/hXoixnPS1gmS93662rWt6G9J
TRBMMJf00K69hehBfrhL8ErLvjNUGd1k5NIHB/vzEzigvk4oF0qRVMPpMW2w2DAxkJTIdLYiTyHk
h5nnO+SZcAekUt9NDIDtJ/o7oAS/kKVMFQXXUagGkTIV1RcsBxRFkQOvvVXh2mZN+hv7J84LQpmi
NdPN2wkWJG+EARDjZXOI0ReQnlB575hGhChSgKQg1nZ1NY3WMsEAhOWrxZqRXDCG3SnORmgvgOtG
EAmyr/1sR4TpNJMojHvFVUFrUS/gIAElnReUm4xxpj5kWA2EsQRe08KTuzQrGekWxrFRcFU2ltGQ
TJej8VJhc8mYjgUbJhzZBhddsARssb2zvukLijICM21hAb6Kasw0S95jN7ilqoS4fM3kx/RZvLWx
ZZiVdObd3rk7NEx7ISs0iOylhfItMb1EF+35Pvyq/Zjru5GQ+5aKyWE7IuJUNO+WVAGKWsgdXpZP
MldT3FBv/mFCK2Pv3J9gMUJyuXgjxhg35kY3e3B3iZ9Hbj5rjcEf4p7ATdTW3UUlyprqlrAaybXS
kkcABI6wr411ap6grrY7Jy+xfgVsnqP2u0xQk6jqFfk98a0BY1z3mQSfIcFM3TfQrhm2XQx2nPWH
ZYj4q7A8C/AsoNUtQa/S6OIiTdOpCNnqZxgtXDbBQ9eTF/vg+OJAwskDZ9XvxKUCvU7zKXXZ1YDI
0dU1X1iVW6rec+BQAxm9fCZVL1uDEkpU2voc/wlMaDb+29OEnZ7iiyFm+GjDzcsapYk+op7OxhAU
lriQMqi3g6t3FmGHcFX9+pjxQNDP8Kh60trMhe4AhtBVNku0mD2IrcKlq9mTCOgEg0ysEWesiZiX
+iCYVD254uZOPVcZ7PKpfx5kvXgMOlZ7gIuC11cAeuSNl1SibnB+X71gxe0tXVd5ldeRB8vgC7yb
KdNO3RzjiRc2vkPrpTYxBHf6D/rUzxI54bjIAuHixr7rLdWOxYuUQTbrFeLw46SExY4TpWL8pb0q
YKc20Cf42i+UAHY5ou8889SlkCcCCS9BIOPjERCVEUEU7MNTykfVoriSokKk6oAb/C77Xm11rCvs
JlKjFCaVSVe52smfrdpkhhh1L+dcoSWjD+2Jtuv2Cafcg/Cj1xwgKstW8nvRrXorZXDENlObfV4s
1GTr5YdRLbnHfhced2Kj+D4r3JHi90hXktPlez9ITxK9IIjJ25EgqpnVv6UWcLdAriDcheJ5E/eJ
4gE1q+ebx0nKgP91Vgvipz4G9adSw7n1XutZzRhf45ZKbWvUSqtDA7oBlQrqklvLelAKajkGu6nV
NEntiAMd37djqLVuwIVA64oFOzHhU9eifvQGXg4NbvwPMPJ/Tc0eh0gWnPhXR/AmpHft55ra3/OZ
SEkFTlYHzGasBnCCd0CRDYsbxmb5mIRHF/w5P2tSzUfzTVKXrLmpJTpSWbq1TL8X3iMLGv62j19A
/W2+x0Ol8RUMbU7JmxMQYOdVmfA034f8C+x0X97GG17hNf3s3Fj2yeGOZRSeT6D/v8MZ+MfCM6Qy
K+QcPrt3ieEvkNo/a/uqzSqzPhDLqD5A8IohbdEehMJ97KQFNdPH0TOVWtcSkjWnn4e/lKZylBJ/
1BwbQ6Mb/LW1Y1ZLLJoDqb85WnoEK9PK2J8K50AQGkiJUZjRJzroEMu8dFtW1OUqG6ksk7yFR2v+
GvjMuBWrWrwQYoH/EeWmFrksZ07Jo1hBozMLhkjbyEKOKEif722sypsMCmBO77GbLgkYEqUSdadU
bxRER3QONSgCRwpZK5XU4xuq23Ps1NKxA0JmXO75fvjMCTqhuuBsVpwGjA1vc+WDGcUV5Jwx9YqG
DyicOkmRHubduBDRhnIxDTx6oINX2Vyxhks0SVfMvUsLgjyxeq+zQyPaJR4gD2AmzQeZVZrCAFnx
n6BSHLeBex6k0U/0+Q6Nmcnud2k4rucy2PdHkDmMXZzeTT/0wO2H9SpA6mYvb+ApsPyn3ccsyALO
Karty/U+eJ0BgzYGIsE1DqWFeuV4oBAsxl11zuXwPbMiB4T6fW0oLJA9u2yQl59fxzsW/BCGZYxe
A7fZ87ZKwYKWQwLccIo+yJvuTKuxBc20gG6iiZNmNRjuYoNW/YiSF0f3mPki2AvyK/guCEefUNKF
90urCaxms8cXpXyerYtRlduaZx72KiOL04LVjB12+GRRaOQ+Puu6/1gJ+iZKyyzEeY507nH+fmxe
hY/AvTPAwWH7xdxyCuppyqTi+noBTYWtDKGcst4pZxiIiW4RLeN7qPTND83mi8n3ktrkiRO2pTwX
0EDOHqaaH3xXlkP0F1ee08Ag9pjR09mR5imNeCLhxOhyjxNyfSPC37ivSX4kRPBRRga8eJ+gePGC
JR9/+xvXkLeSAGcMQqPRqAxkBiICrM4sSNvkMePu/iDgR4p1alkYUZ6ZxvGu/Lg4/A6m+pDBxhZF
HuYaPAqdwynJTTboS8X4wAsRB1dze9P6LzomZ3ewuPH18rJ/NJsXKnBsktY/zDfczWlMCYxuMdF3
6PlUkf2gujIolC10NeNmTvksguYzVOkBllQ7MAOv5L7EusGiFGoWBGMd2tc1VMn0Lf5RKeNh20jv
be6bT4Xp6CrvisGZ/Imy2TpfqP9AZl8Fi4SEizSgooroLTnKUXzOJfkNXGe6FWsfi6k+yUpLEIbX
9Gz7wB8x47CQnh2nIcRqGJkYTwJDl2RVJ55dbJemBTgm3mTtH79nHG94A7gXn+Dl6eh9RRONmTju
QxA68d5Lj6sZiHce+g3Hrnbnf0qFO1jc6C3zuV1IZqXJE5oM61+7C7yPNsNuxIBTip3GFsjFo9S2
S+WJTghsrfeTvKbvtzHwB15eClmerQof9wRCX3YpasF+qrNVi5lFKFOr7HCsC5V8+cecfGJq/5Jw
TIWwd0ePto67T025MwaOtN7VOSwzJBIZ2/jeHNfZathMEPbvKDJJReQ2OwDafxtPh975riQ5Z+of
hJv452UpvQT0jDhgiMfTHw2Hsf3JnED8pI/ipyfqcIaV9ixL3jS4MUWcTCIABFpi/TZyQ5gZ8yHm
m8BtWds7JfrpklC5nGAz2RYPWKkZjXkKWUV2O3OLk2BEa5nYJZBCkNY9/st/guoC+5be5R0tVl38
HhFWcQrCRVcIfv031dGB/wHA0vanouhi80N6bwUXCugNf8GvYhA795vkNQgYIvY10mntyXDAUrkn
KdvSQAPJDQ+wUaUKNtwSOnlOgZioufzDTgFXereuh3lpCwvVpflt/l5tXH89UOv+oGxzvfiBHYdg
Az//2RZmDQpn5w4BYDMAHyugFg3/qhBonDvAgyRXeklzRPCGvXJRraO4Ym59OLqntilWn/Np/CgO
VUMwjxcwdr6JGf163fZm5l4VmGQ7p/asHq/7pKp8uxHopbqSmPVhSSP5wPBaxE8nbl6PUA7alaLU
ea4MT6+iiaeHXf9GihvuQAv6CXgVRcCvtiAdjIjAev1ndgYDswMPh7UwXGzXC5w9kggcRGI/8ptC
jMFdJSDcmH2oWBfOR7z/EV4/7xmML7sghlAuqyabKzRz9e9lJW9UOfHNjNeqxqv2i1RReFmO/p2l
NDOPYHM9ffQ+YBPPS7v80dhWAtMQLRasSix9A5Qpzusu1VWbUtfQbcPEiZ0J+S23DSOVnXkWdsGt
EthUS6U5encwZEGmar3cmZ+zc7vN/tz550KLmogtuj1qkFASLjf2LhuBTyoauZKL6dZbGEak6QgT
4hC+5+9J4mgmEtHnU42WDiW961Qau5CJjzEbPnb0XY61cgVcopBP4xi5jkhrUfy10OVXQUN1ChBc
nelkhUMfizZB6Suom0wYA7wyA7jbbgbEB9mZZJo/xMLdzsp38eN7IU6Y8cYNa956m82HvhBFRpbt
dUew2ZPg6Qag/WO1svw4q2lmykKDjcgbVAYcbDb/qjw1qhFJ/NjmNHarANobKxViMe2D19bYKGvo
nHibS2Eit1tGdOF0/CWIX1a8qvxpFF3vEfuy7BkWurqqhiMpw1fqceJbCgfRk0YGuXtoKKpx8299
B0JsHqXjhF9CeveCV91QyQ4D5kZ2OQXIB2pSgH66K2S3pANV/sSQ2ucChP8C7RpytjfmabuCT2es
8RrD48VGNnm8oSSLlMwpbaLsUUeJ5A4uVMOjO2F96Y5H/WJfR1G+ExB3XYGJryz4sfWFnsv4gFuI
f6bcuAyc/R6XRx+6hTlUPKjMj9C8wnTzytEd6LRmjBNXYsnXv1Z1uJh1tZLkQeQdjWH7B/Ie2hv/
wFWcaV4j8kjRI/DEdVURnvx1ixNGyRJPLzt53SO9hMdtgdNNe1amZwo42bllB3mglFd9u3Aw8BNa
IwKqm+XW/lhS8G9WxJGLY/GgzCCwl1wKOl8o8GsrrkPCWjOLxGpS2mC3rTL6AAJvbU0DwYvEljy9
DtlwArM7mGwZa2ucpRA6HBvhhKlwI50pVgpEGSN0yLOJL7BWoo6EI4PnZRCUbSxPR+1FjVZv8APs
5Evy23IsWnNjPwe8yWoaa/uLPzXBotZUuqiftbfH1UbSQ7G6493/PFt0gsYlu0CCbYSNARSFuXa7
+TJXR5MmgfW3aEiPS127J5kyOIa7enCK2aIml6E4ZhvKtwMmR0a367iEB/AA47KOZ9d2LXtfD8Wj
COYDgoe2NijCTSq9xuSk6Tf+ao2RgwvdyZ+SVxrWk710SnzEYOci6lEeZBro7MMSaLJpjVj3cQ+s
ZAO0CX3pDLg6X+hrCwNzAB4jgmwM0vT1z+lOu1o1FSGSNkCVzReIpqfHEnqu8cSm8E10otLTGKcy
OCmE8iYQiAKljVN0m+yJDF/PlcFXro83E2ho3OVrkzdZuH5M6uk9fR8CREaGMfUPEVOmxBm9N077
rjQO/oVRXR6JuKG+2mbgRwxjN6iuhwJhZd1jdeePBnz7g30pqs+IxBtZHbyQPCYvnD8XjRnJwtGG
XGWKNb9NNYrQzF2sbhOPhg58VOD/6cUF3kh46qmk75qs5zDzvhbAlSTMkBXcykHhUKFnMQ2Dnt3e
tJlmFX1RyM8ivhY8dwmVFMtlzsj9de0l8afjMY0dfIdfIiS8nEWcQesK09fsU/DL3+cBkDqYA+ds
BxiMYCgVSuPO8QXDoyFKi/7JGWdi9kc7oVZYGJyP1GCGJLoNjYbX1YxZEAdqigtmPR8fV4MCMhGg
KECAYmVf0H8goeH/sAWxr/ZqwBNw9bA7HSfaCHfq01tgKGW28ndCh68UiKdb/ZjbZlf6m20HquU5
2mUU6UEAbKfU+amaZ3v9t8g91J4f0zDjJx/X3LHc/1SSqm8RCCx4BKD5IzVgBUoerZr6i64dI4W6
TEmrRjs1/JfDjmdkw9kGjoJDMavZN+pHqoqZ76Z1uAgeTQlKAZAdTGk9HDsD/VAeCY4P71aI6adN
BIts+E5Go5tKNlaLhCrl3XxOcK6CIrdU2xu4FZfPYV/agcrniNLNXLm1T4fsZYMh4XJ5J+vzcUFA
D8NVES9ETKYM4LIxjua97dQXALqnBPkBdNGMA4fVDvqREzFRQdnsDVH9JSupK5QUARmLXp6RMeNu
DfsM+g5qXsKztp/uOFvuNhlrCCd1z5tdZfw3ga9UtJ+wKZJPFrB2q0m1ZvqEYF5vBGw+8IomWN41
io4QuPPYGz6L7uYe3O1P4CA+3rX1oFDHS36SLlI3jSPo4EuJEt2jdiRCsruwclbIotkhzjisu+pL
DXkaiR8Bw+8Z7Tbt6921mN0Fa7u2cdow1YrQJwBQjLmI9sw3eBCVMoALsC5zDooa3JRqJxKFdnua
7DU/OadM8NHV8+KfmxIxp96XCFv0uzRf5l/DXP+RyDn6QgLAzpc5SA/4lYU1dlvdZkQ7oAy4ZSnQ
WZvLhsNfht0h5R/MHUKk9lD8FPUJhSoVmJuGxUnBW1Nkji3VnFsfBVT2lT8LH2GDZPD/BPiFsjHt
/ok/YTyLL/wtKKDF5raySXEj4xMNyehnbBQb//RyMGTIdY6vPnN/feJ9Y4i3a8dFPkBXJdeGof2/
dtnd+Vhsjhm0WJViUBaXAztMwzeOpTfBqDin79COi0338wavkV+inaA+vr0wMVx8aFXpUIBh2M6D
yhtvNjAtZ5UcSzkonC3Olx4QjiF6IKZ322dSkzLi7LYovmYYt6ms48U8/tEXJQ0NxNxNzQu01/dh
nlJZzxJkcnsFIczL9eHzGhqpx2rva8NzLg2z1ZtdoPx1WNMzTTZSJsaCy7grTqr85F1knvxZj9Jh
PTu9gPcVDtSCo7MG6Zhj1WlQKhkaj83MksKBcJE+lMXsryf93ri+3bBf8tw65LhSGvzpqVhGPHeg
8GxpdLwI1PHU6QcCUDKC+TfSh/6NUb//6a17fU55tL3ZFExguUcm9taeeicjV+SwbCvC/weAY5+m
ghUyFuqNU9ptwO3MM09Eh+38VlOxiKf+CDDFZ6dezM76HC2YYhrnDqjmQs6LAGddGig/06rAd/A7
3s2O+rLswoEyIK5jSUorjIVk/N0FPxvgWxxHf7UTc/QX5RjAhtdcXo2Rm3wkx+2pOaeCDSyqPt+7
LDit8/IRSVYgCFpmgnE2vACeD9MbktQjF+XfTDDRooGd0a/KG693ElJZkWwW1hVDYjX/M4bsZhU6
0zXi/Z3sQte1XyZhsT/LkX9itbHEmu3EnMVU1rsEQ++vDU710oS04xqrboFBA96KkgLtBC2H7pqD
fBwC6R7nli3uAAlocs7/DSTV92dB5rueocj/ursp5KjYzA10T/xa017TUVey5TvrR65FfbwEemlq
HFgGBQxtvSg8va/Cofu6tmSOmKHbM9RtDfSKwtPtb2poQHGTkUGmEgNkSjXObtE52CkGFL5S3zEn
Q7slWSzNt6zewVy2q4vwtRGenugRcfmElTsJIlmfFUN/JPojrnXMlScVWSQAPAVZT6q/1w0WbBKm
qdBBsOZ7/3xKMPvquLCroORfI5BeEmcTXDvrF88PYEK2vroZcPLL85TnQyP+o5OoxQ2omTSiQyAu
CA2kiq9EJ2R1//0kvryJr9KPBUIOzkrwsGOgjc8TrTe1SuI18mRZmi3PwIwmB33U0Q0LQx7IOgHA
EmK+Rpo4zmEy867teoki+BBL8tg9YBlsNd+hJAmXSULhQamO4k4h9WivDs8HEcS1Vk8L5pGI8Meu
zizE7ZxkO6liOcRgwxWXypmOiccsi27wnZScIIVclKtjOdIw/e0l9yjdeTAag4CJ1ljsa0NVGkSP
6iRSTz0t27brzZ/OcDfm33T31cq4s2qX1lKudEdmItul0RFckKD7jfj9crIuZInHd4yZXssFe3Cm
Cz6fZ//nGqkdBazIgxJadqUe2F/hWRREm9m1T/Tjl9AMYXu2hqv7b7pJod3EsVKjtt1V5DM9Qj/u
rb0PJ1qpJUBRwNXjY4hdo39UXO5jJwRJnNKPtWVSm6y9oVvjSdXvnjzL2K/M1Pr6MkD/wpOyXPY3
xU7drspDVR8sqAvhH0fu/grJ6zDfV5UX/L5STfWAtjeVQb2HLmS3f/6zu1luTtPZigSjXFaTRzP/
BrKNMPndjuKulMc9qhcDhVtMrNPxOGsqqQ2Sfvq+JWWaYVbLPGxvD8tav501ZI+2DohgTnzoyigH
vwqZceJA0s9XL2t1Vr37BRVgRgAglah+zJVWjUQOJkuJ5+nwPzCOsf8aL7ZNHOnGsloDCuLF0xPM
ZpMBPDc5ByZBIszasTkN+Xwzqp/CYoWfrAUUWEZDu463WDZBT+u/vozLsyfJkJJISWT4T1gi3ur1
Tzg9LRBX1bUWjYiEPpUwO8mC9eocCO68mLNrRB7anbngDuM6WZ4dgWbX2H1DeWLeZLyDeIrlax1G
LudKRNsz4MuP/aPGgUeJgqNXvgBXD4flD6JuzaHTmPPmUBbITxwaOSEutCcF1XMSs8p+NQKUFvHH
pF2VYTI1icv6drfKYdvUUT2qdkWowUoSRAnrX2Vc+8uGxKhBtnRKQm4RQpwIiD+afEjzUl42RLyj
7S0LpkqBZdeVE6XIeDtef4IwLDVmZY64n+R5HAYOr2RXiPjxnBlvGX1Hhe5FOiwLPVv5Li6ZsZJz
rg3dzb7yz/SGu4eNsB1jhsZAHCq03hjymQIQBqybuwl10lHHArqABSQyIVexX5LPGRAggDZQlrtQ
ZQUYqnW7+5rwVv+iBSw++2PQKnuOwofVUS3jwGwOuDZ38VWfkgGTnoVq9Fz2W9JynpvcSZS9ZTHN
rkO+nRSRWQn9tf+pnp00Ed2ziRIDJUqzBpDvweKwkIMGm378EtOadSwk36QkPiBdSjdIxOuFrcH6
Buyo/OaD5uPsXQuxtA6YEuwycdLfrdHMFUk90bgOMcCLy9lZEchn6MrSnAeTUuyBz8dKXYTXqkHc
omf3I9KghpbRVSGWH+FmguyzB9govqxx34S+b7r2zj9/Xd4z542WLwNm+StrWD6P1OLf8CCidlm6
uQE0n+nOsX7mU8+N+pvgwWNFXnu59Yjn9J6pV1XNMJH+ZyGTYedz8v+Bw0OqDl16SDlNDY2ozY6v
Qe35qdGhkHtFpNRmKvtbFrFJdD71XNeoWjGlYXmSAJ8KtOsP6IXT/cUKLxpqs8dYn6rnsPZtTtIR
5/YE5O5ewcmxn+omPxC4hnT2DoGAWnMMdl6VHQNyc5I95Vxgr942f1rU1fP6u25XqsoWubh9/9F1
TkjfN4/amItvXAlC0nRT3j0OZKUsLYOQlgpEXnG1aHXgfie4G3i5IPCm7UkhHbiB/eFWd+4qKqdL
1X1XzniUMAGxb/ZAFn7Oh8BKFKkNH759zCX1KtW368TH1I/oCDqOvo4AS339Pm8PaC9QuIxW9wjI
9/6mGHj1ny6SXSh9Nj7BkXrnKWoCQtLj6L9fYK0sGRs0HkU1ZCqq7XoOUEUjDPPmT+TiR7kI+RR2
eJQbD6uxkTOM9FUkkOBLa+02gO1mvg6gkiG16xnjQsqQiv1G1EiCabdAdTdQIq4UtYc8/K0FDodw
6uTPaFYKRw3MfjKmrTuClPwKDcxhZH6l92Vcc5gPftfVYTasTi1fm4kkF6g8fZ3RoE6BjNW6ftlu
t6kEqlP95Atg6TAe/6sEiXASS3ZJPtsPAm3mRuNy+FItrXYsf1I9PQ+WSn5j+LbndOiEe9xBJdF2
jp4W6fbtj0hi4EOE/EOblRJCEnSL67JSkTlEjk4uqc8N2C70R4ejk0K1CnKhSBQn+v6pEifRJtOE
HI4lN8ucr5w27ta2XBuPsMDB3TTKw5HrYdwXf4YDYUw4aaiOXw7WELT59/whNB1GmwAxSXl1S6Hc
akOnv8zFsbQJsigyHDaGVApi8hhgVzpms+4+MxHKEHuHSX6iDb8izEw/wrrZF8y3eej3UtKylS0z
fia12WpEY898njgqq9IaIziRKuZ0qDvb0cXclB9edKhXZzaWU7OMEEs4oCXvIahObZ0alSTymiaT
rNm+4qzOLXUU8U29lqRv5E33YdTIDaS0kj5m/8kKtk5TIGTvHmpEV8ee5OQiUiB8t5VGpKN1R79b
DfjDSZNQHWkQT1f9ZiTPK8FO+2idsylmvZjIM12S1/rXawTrOnrcXOl/+UVFkQ3Ru5T9f8uvImr7
5tgB5KiczCBLnSVDBRYbRA8wyJ0OwFjGH5Ymhs4LjrAcdQW8ncZHffu0p0Upnp7V9vsXKoe84OuG
L86ViO8/mj5J/l6M0BwS4FbycUrG4G54REDVFctRQ7ZW+AhtEvDD6hWpKCRa2Igc9t5Zw/nXKexb
K4S12J2FLMIGVoebYmNZvmgooIEzGJ8QbGYRYZ8vI6XCylqGFxyhb9JBhSDIB8osWGzR5kLBP14i
JCXKSUhqIWkmPYyBL2krVNf5kEj0ghH6YOdYyGVO98994CY8+lCw9mDzUhzdEl+FWpAKVtZ/o4g2
Oz0AbLTzBAJPa9/fLmIBDlJRgvJPhAp5hCt+6vThqHH6JsHPp+I/3fh85pLGyYS3Ud9OwWWZ0qFD
jzFI6k6ehdOpusJCbWus735zuKE5CjCiN6ZdMyQy2A0OALQ6KMMjNyY1ziS+0M39TKYgXyRGO5e1
c03AHuSO312PI+G0RiDxtVJjcaUFsDmToC+oTh37hNx+OUFRFoBpEnCs6ZkpZoIpC+OHBLQr+HqW
yl+FQbdAxpxF0UYAXEEb22iouxEUz42kR9qYy36ua9m/rjlF5MUHvZulbYQCTAHMk7sIzFcvQ1+M
272KNqGxLYARL6xkR2BhKerXcoaWLBfbvSn78HUwJjm7j5F65JPlw+ovQVVXR5lp5dMNV+FKDf/l
+LbJEsKiGx083xzf9S5YOVRdgdNcqRjagaJ8V6PxbW2mQ7GwvrC7X7gT7PthTIK4NvH3eeMwYa98
8T9tKD2mA/DUePobdUw/hMXtPynub8mwX0pag3ntxg866qqnpGSgYCz/h6ug2Jo3ME9RHKpm7sDb
H7W1FKwPoGHjXmYouJvk2IyDhntmK+Wu7RxpZdIenlD8xHfvwF7WiHve62IXgGMx58YhPVESYHTf
hB5vCiYcm/J9KcHoqyfo2LojinfU4H5fIvNbnelwQpsnmObX3OLRoLogVFQf7BIKYrVK4/lNRoRw
I1FeNipsV/tVs5X1oZSHudYgSbNP0YPKata0YCx1gjX6vZjv6X6oqzYt3cSy2koQoZsm8XGRxcgB
bNGr4AQd9AiWeHnm3eoZDtyvK+8koElfQpcUT5jXcqXMRNK3LVziyG2AspYx3lYSLb88MmW/Vf59
QargToIkqnJqQNpbviTmM+l7UF2nhep8CZYPiKqZ1k+cfupWJC2MbKN2gCv9vptyhtyr1PTErlQZ
nvrcqOgtt5nyXvBRLeNP8Ql4OLS22dGMqUHMO+RGn/Zd7PqHRm9/32aMJVT4SbGzzs3DaKUVBZo8
O8z5pq4itRmE0VjLRDJHddCFgVoZv1LWjMCeLZYnLH+xJXwhUZ6pdXYenF+2/aeVboMe0sEPVQ//
VXaQSOcdCCz0Sc0u/ZMEJ1GbaR+ED75rCRnPDYauimf0apnG1jbsXeFPV5KLK9Gb1ncjBuoe4AFf
XcYLITCBFDGzvzP+NBkAci45zCvgngTTEJKzFgpwLKUuVJYHdOGORiY3zDFOZp9dFTT/qBFhW9qH
Eti2l1Dl0YK6AhFCl15GXRG0o0JDrCNCvgJ3+3P9xvekgMGWGccOyePN45njAK5iN9IcAvRErgz6
pLoWrP+kmetYqi2Zu0Juv7/IDQ4IhXZ6AJ8dFzoD92vC5m2PHE4iWuFBEhMK1K0s/1TdXU0itkY3
n1QzDLV4qwzdw+yutGepJ8wZONXKli95vKrrQCe5Jqss1Ko2upfVAZUHrmAAEET/REjkWhG8xgRc
F/iqxRbuktgKFx+P/dk4Wkg5wT0yy6BPlMXSGTwlU7zbIwV8MJdvXuoywEuvY0/hR9dUsYhLwDZO
tK8CP1pmwWXMN1x1JR4clsVZ8cyDh9F3db2Xiq0RvugsEcYIQ79rEl41HHEgAfWSdmklzj/dzNt9
HttPs4q4/r0ng98NpCUwI2s5ClgeJn16yHhfOro1dtUIvtJgq15x0YLuQDbm3S/JEdsuc4n6WnOq
wNSDte3UBjLfNRWDA69hO0b1L1fZ7yZbp2rkOw6rHD6OP4A6De8PKdVe08L1FHJzyIP1AXVaoh1r
tIUPYbVip1petxOHUSj0ggq+Gk5K0SZeYdDqSj2Bu+U1nfNuyaftTkNnKh5dBYtwIYh3xZiHeWEu
WkdC63CktKf1TJv3AOdSuZlye8knlL27lgDzKzKjmmRFaRtzgFvorjVKwpvH+yFBTdjLGfwd5fvv
MaLJjnA7o1LlpCGjdPUW0IrhPo8teYcuGEzo3dey3Kc5//MZKf4+p7KwNdTvoJ9+D28zxLz2fft6
BLcedVJB0c1uajKlAPBecIupRv7uBOrhq6NQEfGQYH+cs89ooVruqVlg/KOvFnS8EgKkxwm/QSJr
EXc5NX5eMHGHW+IDYp5qdWManQ7BbZj8XTOLcAK4jjHUXzOJur8omJfB/gCYktiE7R/rS1UQlPeY
63OoWxfmbbmkqWHb00uCclH11e0yiTMmbGlfJvQ0s9FIwJgZXwVfhqT4D/yPl0bAXeKDsA0bOl6I
HeqIv9RuCqWsLfg/I28mOpCVviGOcVyr2zZ+nRlMst+5zLA99lk61GoARlsImltmJGHIvqFi17AH
mOj74sMA8QEPo+5Ru39dR7Y6xfsQKx7ZIFTS5jDKzpl3CoPmBtKynyMPnOLwdj9BdQAAYnB1S/PT
p/GAzpJHoGkYzHAj7r8bmbk4eKPpy79QH6pzow9KuyQg2R4es/RdOi6vv6TO31GXr9JhJs8MMjli
Y6/dHXhuXPuEpMiQZUlMzfMmXhjQCmws6lZojKUygbW6OkVkiFS+rJM6+0VPT/YAxhdZ4ovUd3OJ
dNIvPVgfplLbIllBsAioOpigNk5xDJVyVwHZWU6+3Y4Baian37Y5IeGDO8WbzSVUhpDl0eTA68yQ
lAmuKfYFqAlblR2w6xXDvd2VLhg1WceKvvHGmRycDyr0w7LRtN4sWYmSqYUuzQHz67rMO7Q/E2rc
YgdDVrB3Rq1BTPPjmTe+tXbeFvHMD9EkkBGUlE51BdfN1lv7CNKdJ2fzJAqoeTMctp7digkxclaS
fKd4nWS8yYdjnNPco660kIIrJcMwpDrhZjKIk4QQlSs1nH5ZitCcjTymWa7V494jgTJnL2CyzI8c
5CjkShUEkNdhyTt19Qr0oPK1MDeGEIdX9+06Nw0vUCSAH1MUW3wso9TS9XohT8hmTQrubQzNpuJc
wskjEFPR/UrqG7+cWEeIouqm414+q9eMxbdMQC7kDyoKDMdjdpHhF/BNXlFIs2bfs4DK4j+R83QO
ty4s+IWkJ+WqHZX+KbYrFheJgQ2uz6PAfkiWWjxGNoKVHUjkDIMXH6y8izcrHivQVNmo+zdHreQW
etb3lNcFYjqWxZ7gHcF1oLKlt3vXjwbjyOMvMuE9jhRpAPCvbeXYy9A7gVQt/iAxBWz5hOs0ZGMS
aOpRXPbJ179NaxCH0c0BpHJAwEDJdsoy/ccp2zENLaEDv2oEuONDDz+B1HxNUeM/hLMG0j4Js5wu
vAzMx8uQAzqU6pfOAJDF/DzU+lgF1YUy27nIYlMbVpowEKkqkAiz11hVGLovlk9r5UaOe3NQDsp8
re+HcpdYoWTPv8OJDupoPVguudT3JoDfR1jdMv/Oh2I3RmnHc4zjw4fVGsS9bCY5YX9OyPRYEzZ4
q8jAjtgt74AD/2y0OWrVLLlTOZylss8OyOKxy4tGDS8AGYxwTpYPkxznIEZBEHuIOWnNRGkc84K8
QmexBKr2O09ESpf1Rrz9JIlWOV6pW6liTYfopY18WooA7YWnHxvAZWg6h59QieFgPaikdQJx/biU
3L2GYZplV9eUstXwvCexHZJT5QrvaUdrqHoWLqthVAsG+wwiviBHsc0ZUFs0MOZgQHzR9/yBcRLi
EnbxYnJ23mF3QHStLO21X9s46CGbYamrWUdvipqx1J/TRbb4vpr97tJYsUKZmFqtjHX/E5dhI5Jc
bjODMQobpt7zMv/IUDK5DsC0cs6GC/5gSqE/QfLpg5X3GfPJVBjcZrJ9ImKDKd6NJbydfjtulMp9
x/wfYXfo7lRY4qZidSkxrjVKTqfe/R4rp1+JTr3VdlKdBROfQ0Xu7p1+jDp0b1e2cf+Ra4VbZeyy
YWRNr3xc6qLXX73PJsPR19mnOoJ3pW62aaMQfKhKk3bAb+oxK22zroL96YBNH93EPQwMMqW1NTIG
KJnx4w4zk14CPn3hmxJYrEXqD7IlB7elnUXAckXCVMmqaBhIrIOqsXLpat/OrE1pFwsxQwjr4d1E
zk5alZn2csTrXeKk6oKiwHfe90hpIjYYs/aZw/TNtCRnPABWIPAGBbI5F6dEcZPTXAGUrsH+T9m2
tfdwhP2A2Co8INGjIuFY5ApJBJHhMgGuDI/3oKSWEFSN99qmarpySfrH9lOaWxO6thBEitO1FrTc
r5EePy1Q5fc+y9sFtCj0pnDcmVCEhxm5ljPtJdoBEPMdlxr6jS3skkfr1HbWI6h6dujX6QGp57gC
yZCJgVUeo3qCFiS1puVAopE0TpLaUtSLL2XpsPCv2QXVWrtem6sJLEheB7TrQ5yN897SCeuFWMDw
p3ZPBImYaa0hEM8pWI4L3xUryd/PCxQJ6R5VyMZ+tvndxyY7nihhOVJN4x3eLSUk8ncgN497rp2a
1IvW4P4RNazZMtNrmSQV8A0OHU7UxCiR7NNV7s+COdUqOgbE/gfVO7lwWE1/LYUyFZeuDr6CoL3J
0uRH142Op/nhVKIGpKml0wtLwJ4yaUayWN/7OwFJ9dEY+0q/rar+zJzmWgRgfEoWUCsND6ccFX44
U55aO5aEDteBKGwfIYcb4/wwvg5N0vDh9wA8LRO4mBHOsRGpUNEcsrV/SXmBkiD99Im8V3laj0n1
ZDWTh5/9tvST+azcVrMZ3QhkX+TXh0XolNrCKe3eOFBj1dsJXbHVMqHJv+I1hzAHv2vuGnz1fwcl
kpyVCn7AKQZVJlTWs/ziWJJGPGS2qOQPkPjeprXWXS0Axg/GHABbWwn6EloUDpG7wCBXdnOHuCKm
QdZgY9/Kobelzb1yMNb81Pihb4kNwPFi4k7uccg8agfQX+cXMh32pi6lQTG5fckPUGPA/TGbtZ2b
KNGGGlBmCH+qX70jc7CtVLora58IBUkEZDTxCs/N2WT1iWbcAaIhMmHzJ4Hm7VMm9H7RYdAaR8jy
MJn/E2eNl5sPscYqB7tzqmMmUZ3zz1J1KdXochU7MM88bCp03Ch8xQV9DihwU2WgWW8InI/hpL/n
C0AqYKXKqPtDL7QdzxSwj5SO9bzvubVzABNROVGrKCtXdngh8lk53mt+J/3Sq9wKSO1fno5f/XyK
f+Z68kCggQVGAEnObk9EmPjQhdqwzgiZGvJuHEDeXGPMrofYgwo3cuDVXWw12hOnR4JuUr5sOOYS
bliOT2oEw5C+vKBYQIkxzyzM/hnipc3Tbwz+OJ7KDtJXFHatVlz+IChXndul6+UmD7sPzt+Z+0r+
YBM6f3W/bAz7dJHZe2amrK11/WSTXq4bQnX1XPnZgTUERdMYr+JW5zf+uTLw0wdfRYikW58rL8tz
+o1aSAHN48JCHOC8lRcula+eEJfrKso9CRjVGX7m8wj8QAonldcqRHLKjUcuBjhpE1DBkVW6cjAh
H3uTkGaNbcWThP12LRINoM3wphJRUBeYpnbbhJLW5Xh+F+9aZTWYZTp6f//Dsj44vPt5XRYX2zEn
xKgO5CjdlbylrtA2Za4pSWafsr64gLHihVL5k4dPyFGxFfKkHmsTWXULPO/SHJlhPmxXebGaS7ua
iMaR7GuklPCW9szeEOzjGL5KzphhhtIc+hK6kX6rEV00EGRWQrT77qHjBlSQIRXgAJSuzfbpLeS9
Y6bcP2k3o7EME+a8JwQyU8najpaOcOCKC6LldVwo/MOJYSQUqJDDRUoFZub77YxvhRmrSy9aOFVC
BGWYkOB1me1yv9KmmYimRNSCb4NANuy6KWDdvQFddAHk0ObDY28cyBFeYWrylC1T69KSM7lxa7h2
g3o8BSm95R0rJreTN3GEVnBmeg1If4J4l/oB/bsoU1Fn6RrPrxr3rJ3MPUJmkfkJEDRIYFEhOrqU
Ox6YArIfLS3HGlLd9GqfICyA8oTmN0tQWVULqi8FRjKTx8RH++BgCtnV8exxXKvBXmjTBcMwotGS
vJ5rv/IOJV6hhNR1rC4D9CQF0idnd47ircf20XE5B2E+yvy58cT/8ky4RZDEu4M1mq3JgxHzqJw/
vdnGugvhKvLe7zFFePN8uCKX5jRelo3SwEnCX9gYXCY9D1314nQE2/k+ecjOa4+rfaaatSfKFuZC
HY2C8jFH+WTf2rkspmZiLN7xmrnJD9V2NedJv6JfdxnHaVdlyvuiuE7TOhU/BX7uQ2kJ2v1AMNbt
0HiIgRmsbxSwWYbZt+o5NgUu5Ob5VLkCwbb+xtI/OzYZzozY+ADtcPdUYdWtNlNjhScE5JTCrDeh
o341r8CvAWsHePg/5KbmTEnPS0/pqFuSObPbD6+Qy6axYe6ejo462DAiOaYf0b7l32mOOBmdeqGl
rT43WsFWRWpOCruzLhg5bx+ivFl3Ox80yED7XrTchSvVQANwGXd5PV8l2oGTBaZ7jSpL60wPSrYa
g56NN+HB6NhQT5p/OBCT+ACt9zYNZmq2JZnabX7JnHsIFlv49SLXzNwh3vPfmiq+u0tz8qULVmlq
rsaLocsTz8BDsgoue46VAY7GbKMf33W04s2qbTIrx38I6ovPOT/lpp9mnS9pJu8eR/JoIJDxQW/D
ilKlbigDnvHQ4W+mb0OUElOi2WU0R+Tv3zZi6jWkL/Q/9K6FnlfCpYNDgv4pYAbhWvpaDIhIw1I2
UxjIvDwrbCRrwTsLY+QXZNZ3SpYvRKivpCOVf6r4ly3oJ4xya7xWXFEt6QNgImLbwiYPz5vDg+Ma
aqb11iARokrqHkADDrlHRD02keBBC9u+iLGjid4jYbrBLsa9/GM6Iupir5WkQSfdxZ7EmOc20dqx
+vzJEpQ+BzNXknmG9N/UkF1Y7o3BFFcL/GEcp07S6kh4zWgqqGvDtAJTl2Wc7SCOemPf1gJia/XG
rbc+uLUh09B7r6RVZvck5yO81E044WtOWS99iGxBs0Tb6pN+1FSiVgS0t1g+oNvJSBlcUT0cL7nj
jEK/FxAljnMhrZWbbAZgwd4Yc7v098ITuaK6v4lF+Opnkp2kco3+VEoCcMLfadAe8Bv5dy35Pn6A
EBILL3974fYYQDg6+vEdbufX+nX8vdeSPIpns+rZ6QPyQMHmwgSYD4jEd12PjaUNnOKUUyAmWsD1
X3NHTzl4kHhfvrn/DBTL5m2XuwLjwx/pzW9H4pqg0Gn0L1MnhJVm7WQKPDM1s2L0+jmIsNZIjXup
mc+oN2KUb8NCa3u2eDy8KugL9hBPEzUwkCZfJQL0w7jF6AtgX93+lzVuGUasl3UUpSAIB2X23IH9
dDJOtWQaQKs80/n8Iw+o/7FU+A3RSwg1590sKMs2pl+QVbFZVv6FLs6kAbCbZxzYUYJNaMWDHNmR
DT1L8Stl2rXqFEVGIjOxncmzn/K3Tw8AvqXPxjLacg4LK6nmPbHdu1vxJ24mncGqUYI5XQ+XQYE5
u6DABSu1nHw0J7l4ToqqoY8jAniZyyLlRoyFZBu+Qqz8U1pEsf1mLF8TWZ1+nSVn4pa0cChjaNkO
x9IUCAZ+FcGeQOrakQIG/0kOZF0VqyuUHhmI8QseTvS51VP9USDn2FavKBYBqaRMG9r/CbdpeJOC
+xP2I4JnppB0Fg7OHjsLKtH33uBf/97YAozPI1wA36D3bTSMy06ywHUHVN1amD3IZAkk2xP4ZnqZ
0bIgW/rkB8yyX2osfhVNHrVKXv/YQGOezRfof7Ojkl7MuYIUviLS2ZTrNWR9PKl5r/rHbCMUSLxj
l3fQPqEiZZMbTnzMtB+cdWkrZBapp2N8dLFi0WIAvRtutw2vOc6+WogwBN5onAHqOtYzxGqHBdxn
LSW2vnHI6PA55bujJJl1zVJuhOLXdIGhx5MSK+m9HV485suiTQmYCZTbqO9H6xKHXr+GFQrkdhyz
8YQcVdzx5ftqAqP9cGdFxMe6a/ybHm1k1Pq5XI/FvwAF46iNM23Mv7Wjq6Pu8EIwAROQNOv+49Kv
xpdR4e7gS1zouA9XguY5E/Ks881nJsZNuIlO5rriaUYmsW9z6LbpaEDhKSfINWAVV8SJ1cLts3Zw
X81qmUQUqT9E9JBurCS90AhFJ0+crPqqhaAlRD6eYs2ToL4Vl3/Nc7BhIU8d+/ujbJ7DR1oEWZKI
mGTBfiuemIchy0wsVZ6AL9stD/sIQNEbPq1FKstKs+p98G0WqrToQIJ+dh9giBR5noppSsuM/Va9
5gOfrrqr9oyNtB0u5QrkcKAD54JxjB1De/7Ynd3MHK3A0RH9zCLFhRRUPZuENUaIUeWddZ5NB8Zn
Yq8FxmIEOaNxE5pgm/WuJ2twt8ODIiZDHifed9MnCJx1TDKM/OfOsFRWfiMXOWegMKHPvFMvpck+
arYDL4dIJdCWBj0TwCllheWNAIyo9zbuTFuor9ySeYPH+c9NsYo56/eNGYUfNqzdoIYujmubRqsM
nlHiRTRDWijK+GypyVUw1P8i9gW8/cLh+d+4S0gPzQFJmPaog3QPvXs52+D0Wvs3oCtRvJmyGtrT
3Sfq7YiGIar3xZzOLjeG1tJu1a+0XySYUeDUjhuWCzSYYNzTpFaD/mpvTOZnAaib/c3JDBNTkRuA
/ltX6A7NOmLfynYj6K5J+/3eoPj/414Sq8EqHmW1gaMF3ozrMl9YfXvlWRBVpOv4HyXNix1VuQMH
x6h9ihFgAcFn2oeFZqEJp2gZ0AD2BdcfIthtFo8GqgIU3Nt/13PrFag8Yj8IkHpFTWeC5dfESwDh
F2iimlvPIKUyIvdv++92uOSXCiaiEGz8R+Dh7WNyYpttAg31A/5CHnWFZnIktJpxyW+wUoCkweh3
7lo0cOtss682DRdq5vytJuU/JO441H0Zy9hLYhKSYHfN4zSH4PdOpKuEl+jPK8dmVY7xBzz0l7gn
qKba+EpcWfNstN0O5cbH+wTVadjnN78eOrNj77HqE/kdX6L63LB3MQpiEeVcf5mgi4YqGDk/wsYp
IZ0d3ki84rlMixs4LuTy2CsVpl0zt0TF+3nGWCgq69X+Gkzxd8431DFw7Ofj+X8mUWn8RWpC/C7B
DI7U/ACXeB1AUBC7yBt6n+APkvmt/UkVdilwmCEdA3mv2Fwjujb0X/T5ooNctD7OBt+Aw7R0Bd9y
lBauBcMhV1m0wDsyCqUr/iEunBTvfG6f/od8GgFWtN5l6VroXOFEYThpRKg1Qq5mQKGRgaOW/JDF
HT473i8ev/woNq5dCnpx/SDYQGUXEqHhS+2Po53rBixZg8N4oU0K+tPvvM3AIKMDVRbLMA7m0Qmz
YaaiggRi07xOBkUq+vrDNeDd9w2FnGx7hoCTCLMjFJKm00D+LBuVRwOieBZhg4/oPQko6SK3OHxI
uFluU3R5/fzijzdxFn41eCF3HZBt2AVy+1WCcoYmwBgh1vJWLPWoIP8ty21JeZ6fge6vkW5NZEd8
SnqqJ5tyP2quW1Mm7vrR5tKXXpUn8GXD9DK3lt4K//dS+stiJsW5v84d84gV7k1LwURILmuHsOim
o8vywAUjT2xKzeKitOfrcgcZsneKCzGKNx3ADGR1EEMivnROCbQz77Ja5KKzCENtQbjLkatjOyQ5
d2qBHzntv6E6UZNg2fxXC1b/+WIySbAMVTgcfymcLE7XP1C03xqichjastTI9AmQ1mno4nxvP44h
OPDKuHf4yiS0xxcn+CB6X6XIryELEQjc/8+iXTy7bTfxaAO4SMuTf1lFDSLHTVAO+Vm7Oy8d6+6b
SYjJwePJr/lS7f1F3gqFTY7jr1sxUdkbPe5nkwZSEYTQomNJ2Hdhouk9W8T+aGiF5qm8B4Cc/xm7
CG9ild8dYzQGY6+wryN02YDbhhoz9vEJg0SiJCn5Heg8FuuCJcxzgqBwsylkTchmK2+bzBM/iVAR
6vI8zh+DeZ8SgaXTYDf1vGQ6xvU6EqdLpe3u40DhQx6H8LNess2vzEyDWQEdnazC9Ic08v33293S
uPIq1/Pcg+kQas75mSH5+sElTb/i7z7EFvwQw11nq+7clZvRFNVcnuVclsWtdHrDHLXQhiVsvEMd
+daoAmIzH5xs6hKJiZlHV0ZIRvPEtGWFilthCx0Mk5ny1+YdQd+xkT0KQl/QLaUwsUGnqq+MnCmV
orlxgtaSkRKndHjAmVrfYinRCJiEfptctn5e/Zc4C9jI7k+xN30jIOOjMRbdzAjirflrQcDbcaQ1
0ofSfa0AMUy/K2BeveHAJvaw1PoDJaKVu/QjTsRxTCFfj1eXR7iAMXWf7cSOCYWsLeZ8/BO9bRsq
Nz9Fm6TLxw1nwu+VODc2WBehD1JG5NP+EFyozOvnyFJSXw7acnwI6j6OGIpFWLp44OkexTT0MKwF
a+hVoUNWe8XqdpFbtWD5FMp4PUbfX5yvB5A691I8jV3LvGDF3t9Rydwmlo2aOp7f/izdhe8vF8Nc
UY6gA7JcW+re3o35lrlblI2Jvhedrmnc2b+C3Q31YASHpCUYVf26RQBI+6f1eXG3gQT1ojWqnhiA
rLECrFdOuwjuDK0iPl7yDUygOzxPX7BrXfiDZ/fjppHPWyfvSafjEMAaslfGR+FzzAXcZ3lAYm6z
QirrhO6bg7tn47lnon6winYl1SY3Zl8LdwNowXJzNOQQ+BkOBkrO2XSW8UJUpaj1NoSBa1uzVFoI
LmpBoj4g1PDA0tDhnkCwDBpq2Xn/VRNEL7pLSD+N3dbx8uEul72QEo6LmMUYjaDp5LDhfwYkaBKw
bgn4/0TeMpO8QCYQRSIIKqEGK0KthYkTCLCROeCO/sWbkX8JaS+/3Puy6oq4sasiktcfvSsw18nO
cTtpujZ9vRJAQzRWvQck4R0BO2s3zugwxS38R2rb8QZhuYLqGvs8ibYe6qnkEVWhHIw4CxTPCT7Q
DD9ataG4HL8Uo1P1A/yolLWQJk5RefUTg+8QRjC2QfmPN0TYa4S7v3CKIorvE1lHqezD/hX1ZVQX
0yelCZK7Qzc7NsKnXPq4kDHe6nmQgBocoCrgPB0EcSXK/eBgBzZO/+IPtOF64UkUao6KKVt0eaQB
m4hrzB/1arSxo4yt840q07WNO/Vf5hZBtKVzv0x5jihdgMuQRL8tzD4zLaMzKcZbJB/CVQU09tqP
WBQXfFetpKbW86GdS2skUO0T3uqZGdudzVHCdQhcTpJYPvscnIsqyv/Q2AuDC+VWDn5h5tonrzA+
cgFQ6ZNyb8r8UpmNKBFU7NUC4I3CdA70GLkiHy2t74rK0BD5kcXglKp2u2Q3erHIvz8hhaFaNsNN
IpWaEbC+rQYwrG2xNVBzyDXu357MypDhDkxMn1budX647WutGLT6wTdX7I58lttG2wgPfYv7hO4J
TDaWuAZ85Q8UwZnkkXSwIsrKZyWOdHCHF7+OThWvf+bBViUnfyo2JOtEVALicpbtT9KlF6OzwUi8
8XO6oh0tCq+G+mR6dUWJxK7/AnIxKlJYxlG4kmduTVgDlaAP+L+90Ky2+1rl3MrRUtUhlFuVX8FR
qf0YY4Zb3SQJWkyov/TnvoDhrEbmXahWdpc7x9GVy2fZiUYnZjAAQQczssrMX7N0n7Q2ay3UMa1/
oCMu/I46hxUJm/PVC0ACHuwMRXnIm/XKwcq8tN5ZFD0OGHjAZzgyX/ILVUwu4awxNImTZc5e8mYy
2wRMM+QLoBtK3LwVE2vWm+8l2bT4E4w63p32vrbMMNdrycwe9O+DcSRD04mexIPYRH+4bdMyts5T
rfkRBWV+1xnIimo6mhIjxJxfs/Gh4RmY3S3JNhXXqvx0hnDCqAZEToMvrk5m/5owcI1g75xTYLCH
naYWACcJvP2hJiaLAKOAOg9SxACt39ASeGM5+VXLZuGUDE1pHmkDujNShObwGsZnavq6XFnCE9ZQ
i2SVWLVwZXP99tXBgd28SrDU2mCIrCKGMcXx9wKOGvUi8M9aCpO98mByJxWHjzsfWHm3Re3w6z34
x1ktn7jEeY6qHdgqQsW+xWAsJNbP1bF4WW8zbOIuDrr7XQYKdQwwTxJOkWgEKeqPaMDmC6DYdAHG
mxPTYyLuO0J9UWOTbjOiZSXvee4OdUXO5xz75ISBKaikL9mZBKWn9iMcPStiLuleIHgqSq6qSCik
tcSfku8C2aksGQcg48HMmaGKDsx+zzzNrwYcZBJfrIIDsG5u8to0YsK0aiQKknvxvXseq9/BXHX4
/9EntVUiePlW+OKaWf+Ns3S8FzWv3HIPtwAETsdyB1BmgieqfQ81wCbsp1V79YmPLkF4zOkCPgql
j1XbmIVDW9JRJGuAqZ5f8jnSYwn96auPb0B73cvlnJEJud1U4Z0VpjLwRfW7MYyJ1O8b+rHKqDz+
NmZLfEN+2jbzCcMHiWex4izapYb5ZM2k+PclJF92jnx3II6bsibbQwcQ8IuO8mWjeDCXzbLX96DG
6jNTAp843qIrXrmo5P63Uwr6cRsz/W+VUnT99H7dr/zuR+23f7PU1Che2kECvy2nXkFz0pXvIFDh
i33GeQ2xVeC22LJTGapiKJorPQETfsfyUioWBDW2HX11ngQXrOhwHdr90OYl3SPbKzmPsIuQnvDK
4WmHaqxjL12n7bcZH2Wsng+W2tGkheG+gj+fRbeL+Qke+n56Zvylwu4xiz8DHz5QuXDdw1/lC/y8
cfdpNmk5LAF1Eve4IIhfVulMN3gIwzYzhohsWk4aTnqb2niUwGV89hgeKBB64pUSQrY6NLqIeN6N
hPm41KTnNRC7BG/jSxz/5XiZ1IM4TIPsWxxIBdtZYUktiCEcBh+7qvwHTWi+BjEtI22oMLFt4Xci
X+pvGr5MNeuXbkcA7KgZ86r9R1X6+TFOl9IoLJaHDv0Lk26fNP1gvPMb95mmCLffpft+w2/cY1tx
PhgDUTXtimf6xDTHwQfXhNE14jNv+7mRyV4ERh6UJFuRzAmyYuazG3y2zOQCNJNeoZQ6njEybX+S
CHWCeptiqmwMQxYbwMRDfp5/B2VihrkD7Pwy8mv1H+Kx1teZYSY4R4wE26tIft+bHXVgu/lspjNG
ZF+yKuOW0fBVphy36B8mc0GNiwLhejawd7VuQN4rNc0wL7ZC28IM+NMlhNfrl1fOuoUIHQJag/YF
GTbYn7e3qfvkyPDP3LEyeIHX5PZVOZ1P5fZUyPuYqm6VcETmOKemHqdSksm8SrX9LBKX2Hd7Mdpr
WgO0ZmE5qRd7mG8T6FAas8GbCnERAs9sd5siZuIJ2AxpjGpnLdA4cRu2IPME9qkXxwh1XusFS0VY
YfHyPBCW01ZZFl5a1r8+I2UQuOKGEy41hasU6qYJo+dgOe12hNGE0E/TZHhqavh03KvGFk3unv4d
AP/gxv5faAqLNjasjSd0X68XRmjxmZUs6FACgBN6nOLWxmHPdK7fS/H8beTmHMckQ9cGwV2LHAi+
/d//s4X0mxvNYYSq4ygNfGIA1vH1qvR1eBoeG1UOGi3l0wBh8HnjLYQHrlYyD3kGxDY3xtH/X9Vw
3Z8JZsQdH3YamLhiIOWrboGoWe6le5R0GK8gfhk5ym9WqRyryZGvdETwZY+WYIiGMtTLu0sVWyzd
WYahVWWOFrvCD4KpIYhisEu3jmztCIa742GDKdlifGHMYjqxctuCkgt46qFtNbmqSYDYbsKXyXV/
45r3xAPy2gVhYIv4/VePp4oUWZUM5x9mRUHD5t84rOQVp+PjpvNOivp4Ff/wSP+2hhC664whlVkP
xyfKYDU4+Vw7G0E1BgjO4bIfZKw3fYoQTDaqODVnB6VxDe+F5SZOf/ZLmlOLuEScpaofmE7mPVqk
Vkh52dGIn68hrAi97sE5IAI9Cwu0kHOeWpOCZzEXm/fRn8UoJa/orL0VoKkCwhwpCPc9YNNXBDZ7
H+ch6X6oqQgghbwONBt+JbTM3ic9vfTvCYoZgVyeb3pmc6m5NvyiWhOhy3ulza+PDMmDx5nTWR9y
CWM8cCQZ7e80IQ5gELTuToNkph9/OFCoKpzylUjYGIvyh6CFyvuIbhitlqSgul3Az4V2CIRijkv3
Xf+hsFcAeoI8wSsRSVhY27Gq3nJ34gF4M9ZNVAfBIXdRoRsabY19U0ijoo/zLkyOIq7J6YtLjkMS
N6nliYFWL9LCkPggGx/zt1iE2Tul1zWLDfvvNo9vj/7cNJ4IAY7QbvLFUP0+h6sd/68scf2H3z0m
uJwCLz777tBId+Ay6BJ9MvsBHfKYO4UF9Qs+A59tXBySl2ewG8swGaka56T7bhXAsO7Pq5euLo76
uHvfYIHQc5/2OWmcohLOeY8UrbySaO9ZvDMAPvjhEhc3+FM54RVySdGeOlEa1O0e19JHnbXpMA84
citbRKVomB0VscRJI+yvibQI6Oqw76zL7Wi+eIdCcfq/ljOgaR0LO8CA51pp25z02GVxw7wKJqE/
9Uiy+N61/FeJfA/F5Bqlo9prbf1pOA56Iunf3l+7lL5gnilON1XyIxXEimzlDXwKCrJTWezWyzVz
wnisds6mvyDJhx964l2GIgstgmxv9Ka0hOKn+chvV6MU8F31rIs22Ay3nzqeCjssFYO0mjB7yLda
5aRLq64HeMITFtgUjDGj+ztSlRogm4Z1I5ZW6B061/89ZoH1s/M/6B3HcRI6IH/8tb1x8/QhVJzY
4qSBQigFUGaGGbNWscADPWFXRrSzF6DG5STgp6fBzGySjecgnY95LWYjRKRtO7eTN8XtFBsyu4l6
VZKU0/JHxGEltwrRY2Q6bIpEbzGa3vc60Vlmx/cLxDDJngNgKhN/p2054dmYMPqnB+hrqOaepreG
KJ8weDwKarabasUoNuXJMtQEH5iWLwB2KYy5inXK13USWgtiWV7JVmLvUom3XvQla8z9icxuaX0H
Xxxp+SCJCIlu1TVJHz3kAvCGUpUYXPLudmGzReoxPudnsH68E8s+YMReBZHWy39IpPISKCLDp9UP
hJrxTKT9/+z8uTsaaBVr0+b1hcvPnIskIe5nR+t8yJQjfdEVgzDzTdy0X7ECQkbKsvR07qtVDqpl
26oFCSwFWGZTdxXNsPW/J1vVKjVcIqRn0TO5p1OsMlVYG6U/OmXzsdyZQm32jXzlWPt1VBK4X7jI
QupieNzra9Z1OIXQr7XGPc+/Cv9hRJPTPN9HuukY5/BJOBmBXFgeAEpLhRgu995lXcb17BICzhUt
7icX5dMJybaCaxM+ZKTCPh0BLbY6zfWZR8vVFLbiODVeJXi/Bmh2AGEUJjbRZ81ZMBJ0gqcnG7ru
civNCJdTdkXC4/z75ZgPneU06zZdBrbte5riNZ/sVRoqEgd8rGnczgPmsc0Qm7iVeTVKc4LReejs
1VS18OzwC+7YXbKCs0EOQOqkPdMyVZBMWkIBy9ynbolblNiIBES3JbcgM1KiXaA7slUPcY7wxjB9
SHK6nZfdSn+wibz7O3VKoyRD0FwPum1SGMejxKbT4Jhi/DBQHNHJX0wOooXYHAdZJuYZekKSvoCI
THGTn20V/n0eo/VigNM5OAQ/AymyBk3NYA3FvvgyGURb3Y/yWB5IFeigGzoCCbydS40JYSLR8W+V
JR76aCOMjtSaLOphMPdOUGxJhrW9ijxFSpmWMN8iyecxVMV4YfQ+JoOvriDNhOhyRxdfG8DuncMf
Gc1Qayr8Fpdus4prFLzzoLPkEKrP4kK/AgI+SG1cMMa59whma52Su/3RKuq+CFXR9yjcwW1Qax7K
8kgfCRgDqdZs1Su5g2uBYDRTw2EDb4BBuY/ZiP5UF4nvYb0xJ3iBE+hNEU0goLrFzodbwNNFq7B/
Wu9+rblhOyiJL+G8UpX45R98y9mmyN1D2Q6mUHycHSAR0BcabpPi6iCka+2XEf18Pqa4+lf6d22K
Xau/M9JAFplHWh4ezjAibA2PeB/6F7QmTQVwvXL87N5EJnNB4cy0JqukvPEN2DKDVeqWNzbki7no
qWgRFfu2Cs73PRLBsAZnQ25RZICQ/P5Xp6ufosoMkFX8PUp+8BLOuaXKE7rN9HzMLpRBCHU0d/pE
ExuBXrGIDkTpMlILrndaZwYdWsBiD0ct22r/0U5dU2ZELNlZ7hAskcLkfrGueLCqZxNQ1HNbrgK3
7OIrlxE8wmyNzr/9qHVEUw3A1Xr1VVekR4x1iNrS68ELIiTsBcvYa5qSdi7xeSa9KHNACUXvL+CQ
UevghWpeKvNrFYRGGm0+GMz7K0voSr9GLqmikvHRYRiws52eBBrO/aU8zJtuHGnKwUjy2SuLi7hF
2n++KOvMIhEHD3f0TiKUl22yfZBj80P/QkzA1e8KbZnwPi58d/Htf9cr7NwRVNGamSV1qUTrSxTZ
0gtE4hLSEN5/n5IhbulXZq7Tp+gO30P/9Iy64WifI3C2o+MUtHcvKnrhk0mLDO/lwlsD6eACOgWZ
ae508rtn/wLFVUkPJvzTeW7EccbD9lZrilabItuhf5depGD2Z2WbvbgCxPITdgcJHvrlJFTzttv0
G3Ue8J8rvCIeLIjW1IXpqHpKEyCDNss4u5d8eyQndoPB0E7rmCPz7dO7GM2j/OqGMSTQkOh0q4IS
0CgqYxCuzymzzQr+RlasCmgbGmM4GPO/PEq3gZ2RDG8giuP0AyK8b1P/O4sNbX8OjUXccvrzkw0Q
ZPAR1RACaeGvvazy6hn232tQ2VWToQqWxQsGRS81EnLGS2H2Dh7kRRjDYMdyKG0eXo3Js0Z7lV+E
WCCSEJKSZkgUBmpjUsxmYaYTZSSIik8hshBUQf9/JKxj7GHpz5p2FeVR56P+5/1IpX1m8dbgB1Sk
xrc/KzV1bp2jlqaWNMA2XO26VXR8qM9sejH7FCbwXP8e/46a6GnRDn6nzv5XVwjjbfj25YE1OLno
XWPxCck6eJw2nE4X9OhZqNVgICkS43EuJ0m3JtAdTBsdn19qJRKZgOOIV5fIvDfo4TtkmpBohS85
THoeIJWPG6dCwZZrcPgd2Vfc2n/LqyB3wjTRb/u8IdmheQ+vrKG1xpva/Po0AqK/vWNNvHzTWYuM
645jWXeXlgvoNX/noDbIq2OhHoQCSwReTJiZ4LNN6SYgADNnWtWOfZUURSWMAZpyBowG38ELFAZB
DxJLK7fKtrWaRhF/67jkfp7TWG9mHX33921rMh1iWFeiib3Fr6gr3/BrCNPO4ekxZG6pi7kTmgBi
OY8s7oiwQXnLZFWlcFHYA9lSW+2gSd1NdY/Gy2R4fgZrNhz25kxzF8K9Qf9vCU+11UoTmNfscRG/
bOd2MiBmW9MP4+XZxfhD0PS1f9WUBX4irsuP14tWlBs67LagvbxolLnfTBnRutD9GDuftBpy7zDy
2gvGXHIJpDcJ+HhRFh7azacyGdtKwwiqV1FRbKonTAMxuP4d3aqm6jm7evoLdpPWgM0xEjWHevGC
LaGYf17NH4Wm0sIjZpQA1kuYX6fQC069t/WFbTyCCVO5pVhjNxof0zknHDgu1vBk9yRaYsVljUrU
2vDHLMXa4znAa7bN8UxcpB5gOT2MGGR2iRtd8J0ZAdX1P63ADGe0QpzT9QgswwLrLj9BJl6Wy/DM
bgPnMBpWR39oe4G5n+vJODHejM3XsHGi47U27FnMv4JYfvgp9PKIb70DgZ8LeJCl9l7DvzOQ/xYc
5W7FDt6qMv3m30QlTsJclcrBYi7gDQTA84mFkCWiloP6pYjO/0CWKtyqqMDTVciEely4uqsvAlue
f7IkGUO9XKq2twpr9QeMwFJN/xCoJ8gPTZ0gphkdL6ScQIIofOa6Lx42/yerXBi1QlKXvBREAXxA
cSCnqtVaa6pHbpK28EWrRm+y+viyisHZtXwrSR3/UXYZwZ2xWtE0dZHTqlL5mrl3XO4BQpA70oMk
Jyh0Zkbhpx/Csu4HgwT2IZ3Eo5nw9bPABbYBe/2vJMqDIYGBjijJrATPHWma8DM7drIuz8koONJH
x8rjT7OdldU7oVGNOx8GQhvwbTyEcecfe2BwcjZN7VloONI1KOAD/Kg8hcw5c8sXfil40pEzD+mD
iha1ObcyGVFtEgYSRpWPULwRLVXQW1AiMjDheLk1IOs5CnaIbz2f/3ZYEQPh/27rnfbDoFrd9dKo
joRjA1MxwD39tcqqdqEzOqWshQbTDY/7Xj7h0hi63ZWnaSXPakklfEY9nXfs9gZFQqY3QVvVrhSb
UlrkjHJpKZsSWZo99VtHtvTX7MaRS4RnMAjMnIlDs+9wabThTKhRjd8NpxfN4VsPNdNQ8YpO9jCk
NU3Fk8HCmJsi/PnKYH7X0mAVLUKKZg30ZDLXcfNhghbG0QZ6mc5SKK3kdI+Mf+YRjjQQ1YXAMZoX
3ytAZIXli9R4wDykoYcIn4x8OBpL0d0yZOMp0LXECmAmMFLlzcd3O4DIYseGs0AKturSxlsEVSMV
UPUlKaMBvSpYya3I7X9KfYDK7Nkg2f+Za1MLJyo3RT53Rv2PrbiGIB3r9BEIGctIhGX6f63MWbum
hwEwxa/7zkdbjZLMdefe10WKkQu13k1Ya1rKbu3vp1sTS6UMeqrLyZFv8h32FQuPHzoLxFSIm2Tw
Fx2pykV2+MVFMWG9nhsT5wWKfIJVzLb8l5noFAWl3RnbIxNLRUgfm+xhxqcHd6VBSveyZApSKOyp
uNlVfIvkmvcl9KMU2hBxDuLU21byCcFs9aoCiMsCpAu5l7pLqHUBFz3omiq+FQEBa5zcr66Ok7ZK
W9mdnRrlA7lZxvjOsoUsKpYtA03wI4u+6si1QXF762S0eH/eTpEB1AAF9XcZ5b1HJL4QmT6MDXa1
A/blaVGYzzk64fAeou1qyDtPuP46ubaekwh/xP7gm/YBcM5rE4I2Y3eZntBLlHNiInFacaU4THt7
8o4ezs2nhUfMsR5Y4ReaIUqbB+4G1DEYD5hE0mpNOyiu0nzL0c5FBR+qfHvFtYZzsxmTjguJsaj9
J7Saq2TOun2WGGKGuvdaLKAHB6FiP/Q2n2CLaHH3mHXQ/jCqktnpNejrXX9uUYeZTlUb57Y/S6Rb
Zhw8NpSoFnUrLHY12p8Ek68LHMdZpeM9mPsporg1FsrSVY6zJouoUtheMp3gBXofkOSV3bcO8urR
RfyBLivVGVGuTJhISO7QNsjQeJ2Ju4g0JaswgXWJsmdxwG0QyqsdiaPKXtTQX0CS2VTh7Vl7nEnh
9r0uD8sFr2sCN3WUPx0KF6cSTvm/uHFGDmvyzgTOeIYoeZ+rMi7hYdqTRHhlkDQWj6FPWOdnt71o
M+K2aygeQMT3KSzQcCW35IpS86Q8a1gpKkuGALdmhVks+rqcUQKtasmoXLgmymse88vc6a8u+oeN
IFwoXwsQg4hnmApR+rVlAaS+NY+RrktQ5LdHFJIqMvAUrg0jUeDMPW18dxQxokrFgRmVUJQTKyYn
JXz0F6a0s6V+VFnIhqGRSxRXMOXCvMDOJ2wYopNHqT3llpfLFC2DqZgoMdQRaCjnkc6tNBZKNV8Y
WQ7oRSzkCWP8LwRxjY10PeXp052XfvRCmQtthSkbY1r4WyxyQlL7slJ3QkEY0TM3W2Bo3+nc9Ht7
9MizGSa7xc+OzTF7kFmLmcLAa2eprbr2aOoZCwR6zya33CFEA8TAVvdpaBPZsJGM+f/YsCIhNOfk
PtsiMMaR29i8Ycb9VBitvmoAcW6g+mZETvHCJQTA4TO1igNwZHubZbQ2Bfz6p/hKtTFNQSw/aEuq
3fibhFuNxWY8Kowb/ns8kaaYOITfFOS2OYzvS71dLlC6SOeALELf0LBT3yt2gwOwUMzkw7hq9MRh
jSb4d1eYNvtJZXcFwkCJc0RBgBnFWaoP9Yi9PHhC5gzHTdrPdM+2EotRUgg/I/n0EFqhGpZCtMWQ
fyvzPrr+/wuxPEuFRg91qKdJ+f82vtQtsewMj8jcWcB1HcTA+caRLYqHtHA3tk76r2NJY+FfhsFA
QVKouom+e4lysRYCs0nafSBecTKFMcqiOXTt4Kz6YO/Pzi2Qmdp4TFDae+XJPPtpjE+khx2OhFuG
r9VgTrSf6w3S5z+HXfa9gollqnNB9y4NzlGql4+ZLjdQqFOjMgcWPWTuy4sI+QqP9IksosDYZ2AC
BMp1w0+pI4m1btRYFJuN7NIJROlekO4MqeClkvVU0ls9eOENm4Ze0dsRk4/xUw0GilXnBUT03UnE
LCQrHye/2KN8XPYWZRhZqhEtFcyi1DXME91uYVG990eqQrzM0GUxh3IExWlvudt+daRoGgiljS4K
YdcN4nbiGUhiozgaioJhxbTH570OmHjEiLWZGkQaqFDHUwcJryz0sXHd7j3BSyki6M1nFg5b9BBt
vWbsWgZY2HlHk+5wi6XHweE2Vki0BicHRgdGUEdcpcksYtYcmVYjPSbiJB75pwJdbxCW6rzBUBNn
q47GdlEuXgmKRINhZ6T3WP0exSAT5xx3G8Z19HxQt4+As4NOx698rBsBFt0T8YvWa/j8QNWf4eJk
UNKUXtuJS14Qt0UXbz91rcmJKY2R40uavq+7iV/h/VD5oA82gWQx9injP8YCfWE09FqpKQ5z1pLY
xzY6HPET0xyBLDXxzAijls1rN9yMeZyRzfnPk8Rv+1nYte6m2dxBwbS5KdIaeylK4hw1ouALeOD5
6yw7h/TibAJ4O3eEW6iwNRssm/SgvozeIMaaoMt6kFmhbF23LXF2T6t42dRHSeji+jJkZ8K+KATp
FFF+fILusmrhU/JCTb39AmUJw5iVgHpmQRfOCCSJYRvaHAtzCBlD/qSAryZvZ9fR1J3wtoHc/rzs
VqxJKpw53dyqB7HcJI84u9GbNoaS9AFYJ4uwFgA5yaYVF8Znug/MIZrWh6NaKsbBpEkb15Zhr4ui
+aHIly+OXuujzSWPeLsi8x/OdeS9EM8/AFT5vyMxzK4bsfoblAbrX6OJjYKQ0bxSa8fSaDw5YvrY
Ae9tNVxUI1ane92tFzKpju9j9EWx13Aw5NLravdTYR53B9oiXnttsLzCczSfGHDhcI6I1d1eEaJ2
W9lneCRRZQi871D+B9WfTpxRF3vp8dhUNB5qeUTArGeTZA82roYh5PSIipPeeY0rfMu8tYljqDwy
32iiFicC9xNxhu9kGbn+L6omvRwFT/taRi6nzUTKbAcPGIEP8LQsdwZuNyp0LznQNJmaRSTAkuTy
/DZh/uuu+8RTod96Lw4mOOtK4nYoqd9kFOSKTj3f4WdYcGFsszxAq6tAU1w2tM768hjLzlvOcnlz
p3s9HPlu/YwzH/fp37m6hVnz0q6xYXusUinEhvPvs1EOpqjfKN4z02JyMObNm1BMgDsq/K/b0MTe
Xg0deveD53iQPoYJW8h3qyMkFPiYmb6nSNrHIKjfLIvxRReK6RTVIbKrjSjVgd2/9F7kUedpLS27
xVgaHoPWpUo19HLja1EHj8WVsNnk9/K9b8N6LBzsjxvKbN7OdhpMKobuCBXTojOZ+Z70suXcudhQ
gcJndSY/1fGwnqBKuaGkTnfDh3obklyv9oHQFKmNNQCV556sXokqWT+jizPkr+oqJESGecmZixpW
xNesbyy949pZ0pPfHczaA6gNibVK1DIN5WFLomA4ZhLSsH/MX+GeT1N1gq4CLrRXAmyvIBZPQyFY
YG+dchMv/xd8AB3ILOP+XqAnDHy6mA0OMcBhCjvhqnHYyuGVX2Z5x5EjGfFi5m76EFLX7inVPFPm
Czica5SiCbh5VgmC3zU4XW4tAIVbmRrLWt4JF5B3L+EPJxkZqEAWa9CpqJRQ+eSljN79E7tB7OoM
4ntHPM7zqTrGP1MaJZqohVojEaX0q8YMhRjuFkqkdtBC8yhpXSdWOGLS5CAtyJxdbyMXpxbKIfNF
3SptRJTlrWFVVt7OwKwcpEKUq25TunCuYdoqCSG/Tal4TWzz/MKLsR3nhXvubXOJSgDkF9dWX79Y
UjuCOMQGW73p/ILt6es+5awvMyRC1Tkzb3xiyf5QaQbnUDzuH9veaikQ2n7maYPidJsSe/0nN2YQ
Pbkzlugdh0bPgtly8vDHK1WtmS8AVro7n1UIygC67Hv25mYjJEYYAF9ppwLscsyViYPoBvCFTDJx
sUVzqtOpPhQ07ixXWPHjQpLIGnfVu/SbM9VGBY+OfWfuA8HKaoEA56ZYfQ7DcI6CHMp5VGKopVeP
i53aaMBHbWb4D26QKCbQnkAMjXyt9ubbrAUP5p8fww1JQZjqguAKKZ5ic+aU3BK6IQKChKLQQsvk
LOIEx+FH17284SYM0oXE9NVi8n8bS62VDILHMtTwWEmSoMxzvCsI7FCZXhlJrP5dPINhGyra6s9K
sYWzg6TA2zAne3GPQZiV3ysCimdIa35LwkXWKII00yt9Flad9glsEy9xIUAdmHJDCHOXwmKBzAyt
cvFzy54G+llek5LnnANG0tZtIX5jInkc8D8EZpZy5SeOcfjsp2mFOfQ95iHIW253qwRvFwLuI15h
tROyT1EW6j9IZNVhAjcsoAha3+acqoSiTPC0QWTuKcrwg1xQEVaHIFYdyeg4moU/i7ZgF5n84JwQ
Sa37n4m7whD02zLsbxwGN4iRcmHHo7Gjrl/AKXFpHfFUeALaoggg32Ysq8HT+e+Y+ln1ZG2EAGJb
YCoJzSRreWhqBidZXfZClJgX8r/dLXvEICymTXI6HlomFiq6KxNNW2MXxjuYItEh/8HPG458EoFm
NdsjmAKjxKvqwRQY0wNOxKMF7gZidBDu90MGCsfh8rrszq9NV/xe5cp11aSur4DAZ+hRd8s0Fr+Z
4gzRV8haHQxvtn5W/nmXVtj/dgo/UtlLiDshnHJmuogBhmBR70IkPMZ0/bJdIsNd4mxwgrXpMgj2
urziV+NawlH+8+cMDZnRjuqoelbXDPgbeN9sVCVKcbgq6ueqpGnD8odkRNM2+kpzWRM6CgP4BPGb
8OjeSD9Hc0jxGv11c/yzTQOaDFerTBl7m/6qqRpH9TU0lc+xKhMr3+Dv8Ez6LAOfxDus/2oibiy6
NgultJKKOe26iV9uoHOhMT9HlEIJGRYdZbAIymMQTBnQ0WJga7F3Iw3UZMH+GtbMcNVwNoZ692fu
XjwwkDUqF3SYJvuTfMvxxxemwWiFvDXE5FfSwHI0/sKhNkyMHEPpZtLFhaq17tWqnIAvKRvMTG7A
+l3WY0W80k5i1kTeYfv2f7TiiqgDNrYMs9jlGZSRszN06oSowmmJtUK2wEiqckajyRqLduGQz5iU
wQ/nj2T78LDXEddoEYfrAdRqbGMIUsPKAoK+3xQHimN/wWv/gVZntW2cD2/5khST0W3pbkN4AFB7
uivfD5HcotNJQje4iXQCAKPSZyrFaxJ6HoSs4XrlK+GvGGRJ6sYbrfa3stN1P9n1Ih7QgRu/4jGj
VMZkwcy/O3fZoQ16omu1/31z7mK6oP12zUT9EK7fnA30Rhm58npBj9Q6Rdl61JKg5nZFxdGBdBtM
gYH4nlkWK0b30B+KiJBIYkTk6CRsdDYVMN8ImZ9Kf3pHdqgYzlqbwm912M2AbWlPsgFYnNOMPOws
ywO87iiADXfk40LHR+Hr62eAmR4I766UOTfbSeYp9LGv0tF7SBzU//B7ayHl/akIMqSD0/ivgP8y
Ez9KrgIra/wohozqOJqsEuUSa4J0oW901cny/JaMOUmyp/PlUrkimqXg7SEEvT3CQklY83OB2OMI
H2NYkgryuR68WoK81verSGyQr93CLjAe7U8tFOFHN7lA7LZlMKbi5YskqX7n/L2rRAIVxVJk6Cja
/Hm60u51Jhafe9SbO6VWnYX1YzidIKRwXk5v9n5Lq9BAPopL9okqxbeLB9g5Bn4aAGfSog7S7rJ6
ACjYByXW7pin/nragwStC2T2uEizEjBvSQcjEHbEA+Rqme+JxCyb9QwNyt3p+l1m0gRQTw2k9PYm
6wMctEjAIH6HftxdXyOs6JW/gB5pYIselDoqBBlv+HUrXeEUf1uuWc4vErNl1xoroFuON5W5lL0n
BQ4UGw6yL2P+Pjaw2pnbXWgLlrghnNpiN7TuwL3imBBOTgUG9pKC7meM7mvlBK+SYGjArWiqnvRj
eLKQVO5Ro5BDUF4TLNQTfmZZce6jIxhQu/gCsixVLtHUZKQgrYlVvNFs4xTFto+94zltGEOR2Pik
EVGZu3yDkT1lCBKSDO41Gq+ZYBIe71p99nh71Yim3zzGDaWdfOdtZFQdrZhq6xtW2XYD5IpQLNRs
vjprlq7FPWDG5dIJTZWMSVrVUNxmj2lCvyQZdC00rZAkoSb+SGlnPmpVBmnZh5vol1AT4yZTod4W
PYXbzTutKYHzR8qVFo5nUJaWo9ft5BJobU04So97IDxPYtx4beg22EXgu+KtL0QBh3Qn1gwB+8pI
XCWX3LViT10DuUJn2mQgwtANJRuaP+nLMCmjRM+kLU3q5dgguPYm4AhO5smbE/P7zxvxnrBbH74o
fnjKMBPzAFhoSM4nANAwZKeugMsHVbe3ZnsAWUCm26C++aUcJlfB+OT51FRj89Qqrj7eUASKNoNu
K4XR4L8EN8/EwpdMogkCDDzvSnn3OKdhoDCSFy6gUNJkfYs2tTFt0S4ghiVVDbWEgaMMeBG5Ouc9
aTxab8+rdaGQ9lXfuN7+FA9wlLDgtyZ+evdiNcl7fYW10t6lRBtuzck7cvL5lZpJ4RGN/xk2yfgH
h0yu/NU5GvcLN0xzhbc+noY2lRGHZ/4WI73xy6gGFzGvDHfl895Fcu1MULLV4r+R/FUqyrDEMoj/
EoZ/jeKuOkxabeR7iiSpjJkAU8S8kPQEipotua1xDNk7Qoklig6NEd4my21AoFKkPFuASapyMEMA
tFD8smTGyq6pb1pQCAcDexWoem526TA9ynL/mYwaTB8UQYyUn16FqwjulgJaEbvrhTpd+bNG34cP
FcPM8h4ognWD1NENsuwbODPLTewbZHSxk7k5Y6JRJgZEPp0POxzIpjodpDIPJzOAVOuCzF9Jtuha
QyO89wh2aNGjXNMqYfkUskviAIzWXkJaKfqHI7JnkOLNGQg1GOR3wl3f9XhjSn7TPb4Fyu3IahEV
EmwdjywF+fUbXnS3LZjKSPPFOAAjJQrZPSH9dZdgGbkmoYzZA5zANutoFChvo77fPbHcrVdwpbCE
UxtYSNq/ZmheZ25I95kbv7FhOGvCWo1gguKbUpnJhgcS07I8u3Qr91kMd0U8voTvU8YxYQDyyuad
Lpr/gpxM/FG+R3wJXgum6wQMnZYn2ie9tU9hxymxEo8+/+irgnh/xAL2cqYfVlniiW4zTIG03gXR
FeLodLCmWK+c6FhL0w50EaE3ksWKIGGdNV2bmIat/eethctGmpMZs9tPG9z8uy2p58tz8Nmuudrk
YNQBpYu7JhCIuyGNLratdh5wJRF9MaV4edXsMn9Kpd+q/eQ/q1L5dnEmv0QdWlVe6iGaB9l8M/o2
0dC1ivbIVdghV/Fp0BfhQbq//F8/UJxFAxnHaHeEll3crkQQ6zG6+cF/BV6eLFtaJ6TJKDL797WV
ay2yqpGQ0bb7DTp/aWiFeoU5a08rYXicrgRiNvnjhfKzn3phhtYAZJW1alhx1JMmV+OzdX27JCBt
XraqpppiAiQOeuB7dEILSZyI18tr2hc0Y/3HulhR3HG3An4OUjOEfK0R3Nu3RKSuRdHLxvGm0Cdb
36XVAO+1VsRtiG4TJnMjNgdoT3cN+BwJACR3yLHqQYWlKtSoto5bOOgX4isF7Z0AOzjK7AIQcu5+
RSSE5ggVwYuKtlaC2ayQT0dGddjDIGTOIN+y4qqAepuwkcVkgoDdo7xfzhRoGQmSCWeJrGrjrFlI
SJc4XLFFCdZXuL1RqN2uQcD/E2wi/ltaeDnPf4Jg3X9UJcHTG9yycB2xcbTB3aKLvnQ1RrRRGkij
NDDrFdpLYgU2KR+eylgzp6xRsdFhx0iXv3oWfQorahNkPgHnvXPdDEGuaqK4Kwzg2xzQ4TgZ+J+x
n1jsZF8YPhvhhJkfVUI6hS0VWq/8H68R2tEKkoFpfbH0Jj3cTpOhi6pkV/YMEWrNz7iO+pO4BZJN
Shx9qhCOREGiWJbUrbJX+YyOEdxuVpKzw8vZlY/+6ofMlyQe7k2FekOGzQF60anSmm8b2SHHnvl0
Eh7vce13P1RxuLrR9QYWuYD0gfAYBPbdBo+guXKgz8vhokoo+AEslW7sKwUP3XnW9XJzAPa5TzmM
RzPUQRyk7Y22J6atY13wp/KQiSbdBD9zajC6ECYMsj1B3ugQAxXvy2DZ4/kWisPVYfKFZuF6kp4t
Ta9jvbHFECFtODyt/t5mIl3yxVdkB3qGK0Mp6mvJKCfKnDaXhatPVLcwGXC0rmjUeQOM6YHirCiE
MdlydpWlOduL5NJ/t8pyhPNKFu1yniOJJs+9dP5tCkkufz+24R56RwWX5HXlSA5hwpkXjGcEvMoa
JFPVd7c/CMtPGInAMSJvnRdsKe00Fc5K6JWLHJEyMxbnNfrlge1O0+WJF1Y3Tzkt3vf0whbbOFfC
ul5td8qByefmTe94dTtTkt5PEo6GVwM2mma0bSSggwQKiVUrZljcOu02dfGDFEIeM5PMZ4gOpT8E
A4csGyV4rmRXC/HdhCWMiakqSeFktF0S+DQnQERqfwYd5FI7YMeqDNl4CUR8NfTgbljUXk61o5uC
S3ZOwAVn+prCof6TnfZeDV2jVcbkrcmrlIIpc4dfcy4m7x+tLFAktvHsjuogVFszDQCjZLcW+MAi
1qVxnxr3fLy26lJ5u0apIA/7GXIfiyq3mZu7AvqTGjGS2ozphsZFbdoPFyEB5fS2B2Vn5RB6Jkne
+/X8s49qDR9D0YViAt7obGzbmaExpUdpz8izjeSRpJsKyXMzs4uwyX9XGxtAvCwfDhI5d1hcG6LI
OPSywaFNLBgnMzXIVC06kFpOen8MoKuKmqQKjSzjbV6eZwhhQCbIFJu51PA4rEdMrEnqpQzgQUiu
ME4GjWUcpAvrP8q+Btk1IOsqBxSTZ5nz6athpmYnXNENR9faqUapGphka9t8H3WCBVXQKCCl/XVt
BJJryXFJ1+mJaQdUPCtjsd0zOMKsLUgqon70LhNaiCjykNDAa2ALupoVSn7fZsz5weqA5lXA3aIH
6VXAigsyRvjClaWJK3u56et17rJ74LBpDTeL2krxuaKYMQtnqPBRH+LYAyF1swfChv2QnFAoCCJH
d4FDc1eBku681+4HYmI2w+/+om+JmufIHjWC6xAoux8Q+9qkhqn7J+ReTjhocHe+mshGqHnyE97p
pDLIupNv6ml3VqYc6hVu2UY8sBVRRuYNmkJE9EYqjIHGtxhPi2FE9kXLzic+yxll7OU/IZdC6z9G
Z2fgrXugzUlCvPWiOTHiYJkSU82/q5mOjX2yD2ZCNuvhFLv6tRgzW+SjuTD53f54z8WqfefnYp6B
2nvity8dykbEs0Bv2+Nohvkg82EEGVidIPrbDP1Lha6A1xSxbDo5lTVU0hX5DSd04SvHnQbekIlr
CHaXJeytY3/nHrnbZX7boqvF6igCW1stlrI7caIuTWODNocByuQGHQz21CnZdj69RqVq/X+dF15J
RNrC7AiF71FrIqV7eNhzJ1nLmImCP5aH5xhL1pww95vhNhPQwwhtFw0DjotnEOZaasIIHyq6ABwC
dHwr2OO+ddkSDU0fU/IjPH1Q5Ss51O8kXiHBXAvQsMCGemG8Q2hdNx3qD4ooGkeHnDXP9imYV6mF
4S4tVadKWLpn1j+uE2r10YnQesDAWfrD0G8XIG7iJsy8hJY0j1zoJ5zLWzkbWdx+a5Dbts3GdsD8
hNLVKlbDYpVPayvtJ9oaWB1eUGL3m7yFRZoyS7Mnyt6nAdvu4aNhsbWs3B8E2prH8Ur5Ps0fQqd9
Cw5biSGpY37DO8hdB5UMhHR+cSu1xsemgF35o2S7GW3z0zZ3JY3uIi8ZKtgnRx7FZjyakSyLsoUq
YrBTmXOmmeZaNNcdJRqUrIwExOW3wl+QIq6pKtKfg+YNoA/2zCPItD02eDfrLQj8as6B6I79i0hK
9pvG5ffs9kiCR1YvBDhRWVnYCpz/UCFpu9vJky06gN3lTqJ1ntt/NmH77DHofkAIW3KEorzAqy7C
s39Z+cg82FIKANWv/aMI2bfM/ISci9IQXpQdMriGXlrZu9QVsMFs8I/xKk4pDcVG2elxGksH9RBT
gX5PkPTmuTwm24e+3o72ku6W+AIIx+dbtALOFUWltauPcgIsFsrpg3VpLv3PtSUELtApLjQ7cOMo
KpfdRxseIxKc07+lqmU1W1EnEmrXsPCa0aVeXcVYw1pCNAiiWyEEsFXnT0KNu9Z0xX41+bzWi8pY
oYDzSWrOuV2T2mJcTN/qdaj8jUxBO6cSmio4piCpNO58nnYLm/mTLfiEcvSfkfJmTiXcIfUmQBMz
JdouWh88j6a48mueofk0Jxat/QuaUZ9DE2NumSxi5QdxswxCKqL47ZNPGC7Rr73YkPhawddBpQD8
d9G8SLuKJFkRLHIbhrc3gOq5CjKF4tbiCN7Hl7h/ZxB/3XKhyxb6y9f4KBFJDY3TkmjPlSKKfjzO
zJNqoykP9A+jxN9X2qJ2PT3KCQ9/qLaNOHMpq+DkqaqIjA1Bl9c7WjRz4wYtDpOF+vDpVFv4FBkF
/MH15E0rjo8KYspeCXImaB9qF8kE819NJjx+I/MGNdiHX3rtaqn/FS3mpdDJudmlrjcRvl+gbVfY
nfz2Aa3+3SZl0lmfgqKzYo+Au8U8PWxAZMUU9RnI6O1neZ5J1VpJF7pl39npPpA6vr7U+q8rvV8P
5kewbkO99hNxZnameuVt2u6ORcLEQ4ju98Cf+/kYJh5Go7ZUafgOEbhBHXtV6R5Z/9G2ialxD6LN
GB37+hA+VsJVB8gMhMnDJ8ZHnXbpuzh0TM4AbH87SbHJO2P1JbKbrTKz1VdGHj46EMv9jPcf+sBe
O3ra5svBF8BcpHcDPFw9TB/GDV0K8IYbxpFicUa1S2qpV1RdjWY3hUjTH+bWnAzyzpchlOkx0N7/
FiVI74Kg3RtqQlYZchpODat3zlbAkvjXlymyNktXFTqHDHvfmRhBAHXssRQZ1+TYDBrzvDTI1oXd
Sy/gVHLZAva6vid5mP/DNgLVHdHQQsNNL0TAxQkpbdMfYz3Pms/J09HnhC6+A+qXO1f5CNblxSR4
okil7ieeiwyFoRxaubLvNuuTpfO9wLD1+SWFjeW/0ct8io7NpGIyZ4fV8HDZ8jUsYZy+iy+6xRQW
FO00eZr+7dMRHKoTIe9xGdsZliSA8dwY0szqMp1o4jPGTHiYCu0gngHeg0/Z+4cwwdUrNXyTCO4N
79N8hzUkA9mYU7m+RQtl7KMQvaQHy762fqNgdEjvYTi03G/J9prCPQfhSm2gEKxJ5cewfHTPHVGA
t4ZWxJGkHyFcFBwNEdF/42AJp0L78cyNwuzTv4q1MxumoR62kNvCF6CvZJcrLEeJPocLMlMJrnvn
UH8h3ntbCNPrFt+iP3ER9MweqamPtT9Mh4nIw9cxjGElp0s1Bou46p1Skdb60lS3pb7ukvNR6bgn
oWaXQjbUPZDhdzUq1Y7rCTgzDXkbv3pigsl0I9Dw6ArNxnX3T3E1Rrvt7WNVB/RSPPOiUa5Mm1ra
AnlU5kGFAvOYIWJnZk1+x/rQxOUgG14Kbq3XzYtmOP5kVkFrFrekgL9RSYyc5JMsBu1R5Vlusq5i
OwYkfHXmaREfi3YeKVRRcE5Lp/Es4gX69Bi714fE0/x5+H47Bg9LIfUT/eZY5aFMdOdjE5O9TS/S
pc5cmOWI8KSzKtIxxQ5oukhK0Hf1133rqw+iN6fz4+5VaRNVaV1pOmQo9YqbvxsruYYBpwtSDzVa
6cp1Jj++QWQsubFA0nXswC+r3MQR7eJcM2Nx0yppjiBZQgTDRzwRLqDnaZxAqOa7gI5QE90P9uIR
1SAF2GMYW2Dv6VYoiPHTMZlcsCmKWKxruRomlvUhrFuMgh7aJ4SAacsTQ9zjwuFjJi07qbou17IC
g5lNGlJLrnx6aW6g9BUFADF4v3TaHklV586HYvNL1LxVfm1DNmvAoXhFxDZ7TQcbqAJ5zYplsOGG
Hok2Lv7MB2n2ylUvJmme3lgIcDBHUKeazsnbdbFrkvfQQcmJiFTlOAlIV2fBRSWrXkXM+ctP2/Xl
/TerEeT0cnuapu2G9IML20Vr5CAeF7fjkSrqRfq8UzqULdvwxR/WtWUNpBuC7a8QW3Rsw7+apnwa
3eEOWSghLxhRWLbsLLl61ZyqfrCBk71WkSdp5K9inGV/SY8MlzT3jIsgzb4I8fgFjwCJxjF0m5ci
BrKnt+NnVxu7Dq5QV1IBKs44VUeCUDCXeeHkb7bAUnN2IstSqDTEcW1avYHHUcfDS/T2Ihtbpq77
0hqqb9IJylkdfvl4ss0HBwQ15MdQRkPkhcljyJoTyhiZmrrNMFQcrozHTyE9pjI0R0nAt4ErS5y1
SxnHqph7MUi5To44MXXJHhUFLDYIOObeDMlkwQpYQdVy/FauuWPm7A9vsMlGkDP7iZf0f3Fm28N4
c9o6LaKD0Ku2T8fZdKVMV8wP1eTcjCUdNCHBAwnAWLQgwwth7wiv8FJ6Ww/UzidIbEHu3ffyks5j
7LPKfhw9+IHTJd0FyfTGgecvGf7b7okyeGEr4j+CuV9Bqb+O77CuoDJ6ET/+3n+jpsAW4b5qf9ew
tbfkPElGiVbPj1SaRbP6MS1gdDUY9fsQCljeFO1YKSxDSIKl+bVXWhgsC6oDicpwbdAMN6Ycj6tG
FVio5dN9Z4PVSfwwqrWJvLLA1oekw65hzJRFHYFtkz7hjtnQ/jdFRh5i8P9EDqkzceOQ/Fu6yUKt
sg6KudR7nOLFXYl07Zzk9/pzuYOsrPx2jezD+hSnoPtS7Qf+V0kGPLI3XdEZvD3Yeh6h9ZTRjanM
SRjirrnGuz6erz/cIx/tDr7vgjDU9pjlgmK12vzfTzlSP+ZHejNTiF0umeKGWV5Hx5DoLpFE1y/x
Lxy4hosV29WBdywd1BMfmSSo+/Ty+ITG54biU1rSVA8ixTi2BRVnOA1z+Agn3f/tH//J85clldpK
TNX9qpV+y21doYL2KlLSzLej7oNYxoC6mKidBSLsFIxVsxrGKuDMx4Vo90YLmRU8bVVNgzhVOyT+
1BWKHfWY3uPydD8GfI3aLmVp4Wy4bnljAL5Tvxj08pRtbL3oiXVuBBvccUP4Cu9dTb8o5G2QrJgq
twp5iVaer7AVUEZcq7nwXsHYO61J1yj5+eOW0wElev4QVODCzhmozirBm3EhQE3hdyNg2v5a/RmD
8DEmE3WVxbNIDJhThFFBBePF1KX6dYTt514xjsROrjsCDVQMFvIEBEJ96wlKKFQ5jynaKeJs+YcD
J1MMjgHfrHhsncAJlsEOhmOL9K3+ucgp7qXXMldsc+MwyeAn+8uP6VclMLbD7SwFQnYIBtvHtOaN
yaFQmEZcbIN5nsFoxylubkmQ1OMV9UyuegdpuwTHYCeHtYAfcb4fP/0GiL651VWAPwqfQ5UiqX5w
j5FDyHE7w4Ir5T8QwxW5sTz1j6Kx0N4NKHb1zxshlXxOeK/Sa2dR0Jk3i81npZTIF/sPxUf/qKs4
MtD3nvucr3sGtJ+jNJokTOCFR3P8cRpwHDWADFSPbb79lNE6oUqIcLfVgcKJPaqBmyzlJWOlTQih
ab8NbGSkF4ilYgTetKJtCul+a7qoSrewmvkrpEDTN+AMXx3875ZUemYXIhKn9XK9iKV9+XgFya4J
ZT3FD2dQY4g4MMTTETcnqN4YECRMTyMO6S74XxfQ8rDdyI+jERseiycULBvfvCM5f2vMbCGcaJAk
4RaSmgJ5B4gFYmCzZIajM1DYmyfQr3C8KdCX2Nzz6vpRjZBUKqzIZGWQDqwzl5cwEQe+5pVLqIuY
nZbitykzq0L/dCYSSW6a3WaPDc9hLr6KnMve2SmGquy4adpkTCpg3N/qf43PN6BfN6Ms42vOI+pH
Lb/yVZeWxR7gbRhrlDHvkQbqjwC6J3StrrwWogpddMP5KC5a+uumITlVKV+qmuc3NZe3A7fVqx2N
8SpVgDrVq87WU+eYDudgKNXOd114lhonplOqZHDG1KtjNYiebTRtpCTjf1ghKiLKb/h+sl6Pwacu
7aKSHB9klfdtyrz4lejUxiKU7aG4Ne71rjBn92spW3aibXVWPOFPLu2BMdWclDiuE3xtAl6QtIdF
b4myQ6pNVTjgrr7h+isGuKk91TGB2WOo4jBxsncgr/AUB9Jy/KCHJtQqpn8BbWyR2JOK8gYe5j4z
zcdG7FLlxFz5GpBz9fdCyOaiNvygOpZaQCkv6wNCv1ceG3k5ybe1Ur0+IhAEBnJHHYShO+vrQ7O7
C6snXIWFG6JD8jJDChW2jeFKgmuipLGfcH3E3Xyo1+UH2ScGPi5xaDZPicZhXnyOIBtGZzQ+5rfQ
Z4L+CdYjdybgkIj+Y9hJcggBGbrqZz4UXJ1w8Ej9NvBv5Rkz691n2C6Il1b1TGajLmG8TgOVwsin
Lzr94Fhvd07e/XmIinTiDW0U5AQS2mlOnfp/3VMZg+EhQ+/aaRdk7CDfAJFBqBPLHCJjRfGUp5Qc
6kEjNqp0Rwpg/8C38e89o2q3myEF+EYvnWYKU80F5raVT/eZS/gf8O8wzpPjEvwTd2yUeMGUDxOV
yrK3xHFVz8JXjGx2cErwsEs1jtTIwETE3D2HOYS7ErOWFptl+RgB80eI5w99GoQYK2mHp7z/tTI+
qWTmf/biJk5DDWW4MW/qN9pFnrufVMCIkEEENp2Y3iXbW/J3Yht/+fyF58MbgB8hbTG7oRG6pS7J
od844uJ+FzVJujHuh2WI0e1qgZWQMi1fnVQab0atH6BH+STC1jmGredOzWzxmkIGYbDP+hCHYCWZ
0SWQG6J1Kd6u59gyNk01ll/9tLfc8AFMXWS9Ie5+U49lhAyaTAWypZUHqOA8ArBBM6PugRc32koE
l3AClBBwSxdCna0oTj4nTx/M6o+skwymo4BFTOKC7TvXMACNUFE3RVJmI4tl2FmkZxNjQKQpD13x
HG2RYgWcaLvEvDer9MP0i4YgUipm0MslfasxiTM23g0PzYolzcj1mZ6a+NkwpCYjB/MELw9PwvKE
FMouNsrWuYFUUYx18M467EjKEeJ6PtZP/dSY5mSkWYaHuY8y0lmeDIlWSEre2AnjMY/ACPhQLqVl
lNvrC+/n7OKYS2GhS8XyeEhfukBuckiIsbN5H71FyOB5z0GfxoidA2a8XFzfP0Sck2eqG8n0YqYZ
ixGmF9h/zdMU/f0uNT7GEXG/1D6U1574xljPF2FviW2IEevPFCNOiag6WzRZx8KuLqmMRWFYB6eS
06PO8gtPOQeF7Lt8uD8T+r7DRP9fLiGfo2y1dY0NA4v/a0xKTNM06UsVLFwIiD7D2aLLpZtOUZtp
09oTI6Z0gGVVCPX/pnWA0DNKekP/PuEVSRluKWKUCvgT7jGHkYUojmeIaFgM3w4KwjhURLqDxcp5
9s2kOboYIUgWaCKnYKp+M0cVIabXAukhlPUJoy8FdRL4CHcIkMvltRAx8SITP2QvfMZ35Ho2cela
yWgZ+lVJMJBt/T7YM9syddJpfr/jOITkGi6u9tfVak2B5HGUJiHnVewyAmRirlDOzu9pwzEcAXVo
voSa099CVuGMBr8kvmQMTlO7oqeGQb6DrRrE0C/q0F574Kv0EL9qOOLVfcAT+CiXhKpB5J+EhaKS
9dF0luTeyruCmodDecKBUsaNXp2P7W22a51Avjn4Hzvfr2rPaRSmiubxCxwIfBKYi7xZtjpw119i
0dQh9+xUEmWxxyhz43JW5FsZF7ESwtcEG9KYriAQjspLximwfPfPrP9YJsLr1Gzn035+1+ZElwcN
2eTGJCkAdH1r31qjExct4+bfisrOKaahZpmR+VYCSqn5E+aNaFtvi9GCMhctDRyCzBKf1X0fX2aT
HQ0XSCFeCtTv+I+lVFN9v0hDgZa1rl5FR7GnZwiHdlYvc06wCKzumBslJSmM7WbISOPa8QPVlf2Q
nhFw6pwHK4En7VDL69SKVkTUGGC5B1eyCaH5WX7mriOuviPXnrmHrUO59fp97vVXU+59SQnq3czR
jpQoCDLwNAN6McxPGYCXK8ojOM4LKWBvXfBVzx88lcHeFF922n3oLolSIAiyMdwUqUv6uUtv4VbT
8Ss2+6uA7kBxC+XRhJZYbYoOqjYGrueLkSLvAmVxpzUTJvx3RW2X2VNVlHYij1Hm2G09flohvg3+
+6XJnmfqNPuPADoMRkk5VrveAvXmJZvCho1emYKj92kwF9PgyuOSKX4ATe2iYULwQalra93lhTfZ
dc8yp6Wfth1e1pY8aGjmO4scyubE+fOAlmEhmoLrEnKqU6FdOhWFoyH7RoIsWGTaSGcSeGFctp5Q
tiK0XtoHtYffCs2v3xabncuJhyC+88iDAN6K8wLHMxJirXekpjdgtC6zOhCkFhAMfXUnpEFm1rYv
g82ubY4898OKTKEQK0VmyPSA3RzdzEz/ezazjjgZ30pQjTGmstAf47v+V4NAFePJSQRi3BIXn7pP
bUxngoy4gFn1Ei2zoPrQjyINQCYvKyrUBYh0nltwqvxxg+h3OBuhouRcxz9BeEW3s9d7rO6fMKBu
fpQyigDErnP0w7+K6quNR17ID104W5JZgtwDUnGgEvfO2DM1F7nGNiBr7OVrtvaK8k0U9uJaN1aN
oxX3gOPun8u8rkkn3MtoU+FCmM/agcXElUIm6HqcMH/hDja0BgahHY+L50KeE03o7VSToM0yjJOd
eaKPan374m7ud+46VuW0+feib39odarGuSSrHa5DUFFr7w4/P+RR6W38scHWTwNDv7YgWhnKYGTO
UYlm57sX54lz2aFgDP6jghuDAlk+zR9a3rC9qCbtMxLiNHBkaXX18FAS/4EGLCAACCqS4L1cF8Or
xdpl5wwHCV1+8CbrFfIOVQXQZyrgF+/2cKmIhZTbRIbehVul5BQkj0fPR8TAvuQGzWBW+a+dJ675
04d2XzorRG0AQpgF9AFWDIukYhoOQBgUw9VFr6B1J1S1tjhkIvijDlJ3uhkeo3bIsVutOlD/86hH
GWCPBL2eWJuHsdW9mvLfdLXKmNWMS4l1Y3b908pw0j9f+LcZ9kSnvEWjPB1duHaYnZPJVBayKfIP
7TvgKLndk3N6hIxjiqtJFzcuytjcW5kWmeXJ+x9S/89vLH0mFMbdvnIvPpoNy5/YkuvB15726eB8
//QSYgESfA4NZps5DkFnsC5VqHGbVqycaZCjAolMgugWvuVc0z1s/szrdVkd8spLTUqiEyydZhNa
SWYFyz771qvgCKqUGBxhHc52/chNkGWhA9P493dpuWWv7TrPYwR8eRYxfYo3JOxb/7gVZptrV8wc
bI+9FPwHDDki4sP//IGmGCFNsTYc7z+sFcHKkEln1CD2bU7mrLsYPuYBLg5osJxYM9F7Ix4t6ISa
UXGr3MD4r+x7PnFPUe4p+IWpdd5KAXrgau51nSv5wrvIVKSJ5e4p/9386JWvCs6fT3L6vox7Z0Wg
LSXjV+m8puWWBd7LBx3yoraW6xosyOk76/oyASB0n2vv1sG41g0KMhAz2xxCHft7BuabTUWWypBd
w0Fcfnat2Mfs3axWErv+/aDD1sbnaQH4DarZLBDPmVJqJ7x++5Y4ICHmi47LVLJTyQDAwY+NqI9t
JdokKwnRtCnIanLi+3rfJMiKug5UaNN5COtXHI6rn7ckuM/STee19lGxOnosTAoIHiblnaFHEZhs
huuWoIPnagNSHktTrfbC8vDEvbe/SrxMKdrL3b5MHgsWkGz9wnx1KSFb8X1ZssJfx8FocqdCOI6t
HwgL0ooxwZOXHFhxEDZvzd5WHRSbj3Bs3pa82VawgyCTSNRlct4Hfy41rF8qSyXo0PxmexS8AhaM
lVcGstT0+QfQvz7GCi0KmgdPnBICKBzKoqeGtKL9toXu8SbifLiHqNkJs9H9x30SD7FEvZgS58+q
f4o4rxRmvPXfvSYxPatbrYLDLrFTmNMcsG6vDbXDcjIc8mlQTF9pZLkMRPEP2YWuJDZTbitmR/We
BP3GUHefZiuu+wSejSyIirmyOQi2oNF8dBe/BSKM485D2z126/TYbRk3c/RbjJaUJagKC260yOEw
bN1/v+TrM0jBQajQBmrFlqssZ7c3iB7cEq55h94Yrm0Wu7TNZUzk6IVTCrfapIJoLVxxUVvpBOVs
s7toM0dDE5P3qJIQrFRlbYFol/uxoKHJrBNBHmhUtqdNQCLHAF4JH1KYPX5ng/2IBfsYUnIVmwLV
PNS7gNc5d7rxq4hzsLtGB7PKqbnCAgF3S927svPxOGOInmJ9CAP9o4U/KgtNgJhXAkUElnmrzM8Q
2T1CWys7RN2R8Cj4v4FNz29iFcamx4HxNrp7nBwSoHR8YM747tMtbsDRoRPOxVlq2BjGzgrhR0zx
wg1zniaS759Xu5PzUX1WukWQgG+WKyA3TDTIMX6d0FyXqwFfGukfoX6cJFIPRx3MiZgVoc1H4U/2
srPHXBtRh+y6gBgdjW6qlJpoGdFDMmoaZPqyK1qHx/GeotOlNuhJXgTTp+U1cl3szDp+vnSxo4O7
tpDtACV7peK2ooEAkgRxyrDjIqWCteZdfa77r1FmC/ko2NqarPn67YJ8i6ZJ1kWUHb8v/0nPCDod
vNKjs1sckoHeNQE5nnX4RXI8Ro9ggwKtRHlzbwGogxc8cB2YMN419BS7f5NNNCXfVn5HpeTn1Rza
W4MU1I6ac++RCX2g+yGEs3IbMSZuSKLPz9anMOdi3mgWAi5NvWoG+GjFEcLpbtFJYE3U+H9WebaV
bp1d0Fb5hatUbbnOQpwYF6hKCsIZ7e8/+Rl/Uh//C0jpRjDhF3rQeF1Wr+g83KVn3qNN2o59ziKp
MAC6kD/PNVXTzdzSBQfxADOP3rAkPrIQG+XpWr7T4zfHkWOAUuDKVVeIU2PGg5TYy2AHg/HPk9jr
hIMrOcC/OpHXiXLggH8q8TuI32SjWtYaU5sTQfQMfVj3gI/7otIRjNOl92w/gjLDEcAYcJKJdUrW
mNXD5lUXyyo38YqYAmgp/N4vBcLu7AA7QxskyKzKJMZEs/l04h2Qlnil68ews+/kfxS92NGL/XLJ
k8y8qmf3NwQUvJs0HZWodH9HJy+I+2MCnprrn5YY7UbNvuMcsf5kocNpJqK/jMFmFtAyAREsH29P
ywccKAzxOeNIuYdLBuwWaTYlAwWr1YtIlq762YCBjVY0Bsz5myNB4zZODBqhxaAgLubtFpNAF3mj
Xq4FEs0rSg1g1Rr40KFpRClYrToWFcLonZqXTpQhaVePz0A4eXUfZxeJytawqA7nIlFNK27TV/7Y
sxCc2iu8wvRX4b5g7g1V2Zt/ewippu45BQiQ7nuFRJU17wAwYjqkS+UiYx6X2Z4Z8PekSZbkY5n9
HEc5LDaCLFEpH+7Fyo8cxayORM3oWBl+4OWCeQVhC2eYKd9jBvZj9FJKJxuOA4usL2CRoq+DjB4L
QsfFeI95WhXz4GIHb/J/JTIQLfN8k8oLpOMGkrGQfySXfkchTfbNxJUhIM5eSPUdpH2+GP9rQIGP
3kyTNS0w3Zxymzuyprdw8/wIiwmarokCkHweQrhZnz4kgRKgoixlxdbSkFV9JnZVUs7MtKmbYI0o
FZl0GeVwS7oM8KUXOigDGAbQG/JIKKtBLQuLNdjO4ymtlU52/ky8CFo4YOxIl0KfggjHBlltQFA5
wSAqPcJFtnPpBwTNs0dkzU+MI1zQQokm3F/d2puGdC3altVt0EpsfJSsBX/djfXEjz+ynusLluSC
OO7lK05RNzQyKxwU4UuV1uplR78oGos7FUSD1OgP0GOV/+KuHJhRAg3mJHjiuql4Jl3Tj4HO6Zqq
AXvRRTcqvpY81XrtEJHwL+Fv5jgOh3LQjQCRwKDTDuEjbU92ummT4/ACPcTQGYAsNpGB2HnED8Qy
3Ey7f2KrM6A7ZKnoWp2AxbE85sbGpjRLqOaa0GfqMS3kakA8ame48w8lVTWvbFtGEoWjzNwPsZvD
zzV48wabzplqK6Jvkjw2IASzixlt4IL2cF3j30uP+fU31hzDR/MBNoYC7MacVN9NX6ltAopytLLK
NXKoNWiV8h5CTKVZAMBIFErsLfHVBue70ZKB2Ucv+ubgv816l6oOa/udc3Rvoik8qqvqk9QXtM4e
50iAvFyfp6qifPWWxvkNRoL3oxCZIT3bHyQoywatFnqIIZMryykFVsbz+PgSCckmv2VDS2gcSbjj
yyNbZDgBagxmK1hv1GbuVFiuqJziWyXkbwdIinqrL1INjfWz2be82XnoViBkDSnlul+OHJTgfsYl
RgfLyUbxldXrVGLXgpjUjRZmndtqKAWyBFbAK2aj8wn4Oe0EbNRk3/Q4S5TshEq4dltrsQJoBGFi
URH/MLHhcRu7zJJP89t4YiC9ZafnDII7uZ3F7Wt6oFlHtoa9KmxaPLwr7bZ5m44md4f9HtlAPSxk
WfM4qCbEsG6bCjxyhLjNc8Mf76vLVvKZy19zwZbRw3RCj6VPf6T1+yBWhWnBK4lm3Xgj/ijAo56P
QLIu4JzycUkUI4w6GQb1oA02oMMyFNFDT7RFtWwkB/f9s7zSBdEG7+TpW/OUxWpXfPN+9D+sg7Xd
EH3vH+QMRBhyKao5CaZkfgf3c39v9aDKI2zy7ZgOUuTMMgh5QuFmDUXOzm/XmuCAzPCJKCJhwyqq
kghwP2DWUTqu/+gErR6KcpfpGJbYjc1h0rozswiTE2/EHoObhuOqzKWpLRsInX19vyZP/iDxMOOm
2i7Ho2tAXkwYiTRnJCoNO9mgZ0qzS6g/HDDiqjStSYzkytCMMhHsHz/vGE8AARuSZbPvDoidq5XB
01O1F8izVbu7zs5Mpc9dSMl0tdPhW+kw7CG61wvB3BEZl6GEgDgikAe9kjz7uPeV7bOvvRmTv3Ak
P2NJaEKVsYFZUl0vTMI3dR33WftZek44ww5LEW+jqTOUnvy+Y5188XU9Mk1nJd1EdSeFvBV3skFo
1H4+bcZdGnB93VxnD8d9l3sK9l2+yMBGcJNrOzN9l8i+NENYx7ld+a30449qlQNFAXJsWxEDqqKo
MKfc5/gD0/xprAcGLnKWsfZAlSo2DCv/4qgXLXzyRIxTby6Or5g1HRrt+UqrmuPC+a43p8A6qVTB
b3iVA6vm88mlG4TaV1q4VlZgXcpXZmdPgyenSSTCUSxboBIS1TFP98SxjMosStcC2rHVwcn8TH4A
UxncbxipXoK6ajCeOFORWs5yRHI3sOc3Si9EEIioStWj2CyZVZyEgWOJ0mckW0j6/2fQT1un0uWA
TmKnbF2o2wqOB7q4W2N0y2KImBL1w/kIWzwGp1+24hbgwTppowGGi9MNuWbCDPB70xrd1fLLVnGW
lBn7HEi9HybDVaP/U2ANDsQINHodbT5pOXg/eVNWCKeyMUWdxc4/DMkisqavLfEDyykPrQKnnUl3
nbyp9u/266kBj11IizWOrHJ9f+C7pCFrZO1I0eJOikHlWaPu/VzjMQ01AxvGWr5CkK1zKJ8fjDgq
BFw1Uk8Fz/zbu66sEJmjIY3koWZDX0skqdtFQAzdSc3AxerBEV7LFWrdwVcy3tj3turq/N5E6LEx
LyEA/rIr7oQbOBekqZME6IZi4qgl9El3HFvNyWIQrdYkqRT4ez+jg1QUYtAiknfDw9L1DIxgGMSO
I7je0N3YXy2B6ttZxiuoU8WgrnLj2NxF/jqLVUrLNld5poPVQ7f59xikgwi7lOuYtjnldng7DnFL
Y19qbppTQcwoWC4Vr8SIUCTfprVNmfc/k+oO0qkvN5gKQ6xhQUb+i3aIohPyzQfV//aiJRMp3lpR
o3G1LPEX63kriXvxPgz6icRhdh832MAF6DKRJL17KH1mcW8WNug7kd7h6xbzPWVcATMyxF+1QqLm
sKzTxufFHOFHj8StheB7KDkj4XilweApLmHgzghg0UrvDf7TJg6MXdZco0rPEfYt/ya+Uwcp9KPn
gS1jtBYSLoscUp/QE0PeaTGeNkvqEV6dlu9yxsE8m5BjZRuWwGMvR9Gk8jzquCeOL31lkkoIQzf5
ohXURk5V2Ug5uy6HZWODE0P67p1zRntUn+sy1Me2FhCT56/ZDQJMBT7HELvdKluko4OJDaMgbLrg
HLFXpTkK+WVQWHIU932OaaM+l6RnHECxpOsdAvwytp4p2IDiuIT8W9jTV3OYcwOpTs1kS1pvsl8i
w6opyx533CYmeFVKzw5pH/Dg3sjAzPJHPrZ8QaZD9z3oo4NZ9x4+1HFYM5IWMDNjZ99JKFQIomRI
SLmTo3g5jQwKwgxqUg34oPb50mqVAHwHP59vqAPjEs7ri0waSBxYXXZmu7TqVfVzxA==
`pragma protect end_protected
