`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FhZzrgSh8OPLnztyUZFhrhJo3xch/bTsmJfqAzmX065l6CdVuFpVgrKGULMQEJ1ys7XqxFY7emfB
WIXjPRMd6Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gFX5jfk/AtzbIDwK41g5tNqVz/VZklNdIMtZqCRTBlNmbvXCwfDAed188EPD5XEbLJ0qsVg7x45G
NoGrcPkUugPXEc7gcDLBRTJIy6jDrN390uyG2A3n/rFVveh6leWOTpXF6BuB+ahUx+DzrqjVRlJ+
ELrbTl5yr4YH4dGZw0Q=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
H3OqSET2gCchlD37lXc1bMABSFAJz5x07fu1LMiEU28xF+/hqHMhYhbDbyxGRNc3b+c3LG4JkrfI
2S25b4vX7tIs0W+nRSiXE7GDOlH2AH/FvSkr4rJDHatzxXHkwjMFNsWh11KDGWJCdBWoiL2IQA43
C/ws0W4W+aHXN8p6DR+tk5hU6S63m/71gP3a0v3iRzxsJdUAs1aqPKEdNPa3CYOi5SkB0pB3Lm3g
deYJqGW6Y39u6YPox1OKkjaVQ7tQW6AOmVDgZCayw9bV3Glc6pT6WS1OH5IsuvDwnSnwtFO8lAPg
oo0d8vnywZ1NGufF8dwGYx11dMfG7m04z5U75A==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Yiplpz0y5VoKgRNw/JFl1cz8trozfHRAcuplGlkytSGxFZJq4OQbLGvsfV9dGiNmOjEdHccgvcDL
MDFwUnbx4E7uGet54Q/JiLDNIMlEePU3cpJtqEPatvKWj5jDP5ymLN+slEFKbo3i9RSiVVuhmFxB
u6pb4BT7+Mor94A2ml1nIKO8hK1IHX4T9xsedR15G+cjlZWXfIlMciZLiYIeDcCaeiVRTTre/Q3o
L2MACWvH1JXQCIN/tRe7va9F6PJr1x4z/H1T/PsJ62UgP3Zl9DJVuiZMo7/8pr6jiWhIuNRZe1/H
KgvBLrIqnE9mCOZpi1C9+FbKEPGzkaQJmIr3aw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYrRrgTX9TeoOzXxehPIFgBOr8WABrM0PlMgLC2xgLBhiVADpzC9JCNgwdH41b7NgvVEeFA8jTGh
y2MQhjHUaR+1raRx/gHHVFVAo0NZXl9CqcnYbv/meU0zkJRES9gSghWCAMSCVU5fNlDS6MxUxtRD
cagVQq2b3RpYOQLHvz4+nC8sUNjkw1vSCM03vd9ZdU/rjTyGN7F/LcXayvpX5K+7jncQGlTXlbrX
wqKuksHdtdSf/99Odo6ERN8mhN8cpow8uVtcf/PQKdcX1eXLCogOygJ/SjMhLNltxqTh5wbwFPzv
cUW8B0vg7xQRcgxck4AJtXuC+OYviaC1NECmMA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nOUGCmVwWwwTcRnoxTFYwWaBWIxepQyRY25WDrt/txHgY8x8FfAGSfw9jcwCVOdXr1QGhXxKJgwc
DF0kgDHz+pyv4liA4NroqbkJrZKGk3t8OE0WgB/qMov0acdtx1CJhhwtt2pZEGZB0s24NhZolXIA
87c26v3XFh2f7wY2XzM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gJC43rWQOdIrsnf0yF3xT2Inssolfj/Y1c2kb7j6XuC1DYjicNBp5fNt5GE3qy+dl6PRq+u0wyGR
J1CJFI6ZXXE3RRw3Jvs4Lv92BL6A1/+7lauMpeoBpCUwkuDBa6fumcydNTQav44SGmVUqQo+hkdW
57/3TVppH2VjkPcqLf+ftwCgc20g9FeNCbSj9i5o7HfNpETn4+lV1KC3VzqCiEhfBPGUBxFEWHk3
bNZHLOsBsRf5aXqKNItCuqGoR+rl2x1fTza3d1y5f0JmIZLlND2F6NkDAsobyMyxF3pm5VdoO/jE
c5vVIaPD/H5Pa2lXqKha7K6xWIKRilD2i9945A==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
HGjAmlPUKcMH7gI/f2nhktRPAgsh0yTOp/Br3k3fEMreBMGSMgfIMSX/J1KqekIhKui+utI3Y0Am
P+dOdDmTxE0qr1Ucsrw8/U41qjWiPywP/J1P1nx4r191H/DjppSB/jbNyH613Jx1BjOdshucTSFT
ytDF4lVE3No3ZUD2ik0dS4mxCTsBziN3YsmbTBdv3PX3gdRFf0JC4UT0OOylCpyvYUdOtYDbeh+o
TjSnjiI+xhJYTTiMFRcmAcW78uqojCWgp76vheFvUTqiSAF9L7GvtkldXGLVcUq/46kTLz5dJMUO
3Nsa5fltFURbpd2+PlAlxyQEYR0qDsXHD6a8ww==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 7440)
`pragma protect data_block
mMlusbO7+khIDW9cgdhi5LuOnFHLlJ85XWXf8pZhmI5TB4zy88EjY0Qf61TR9Mp4mLv967cFAJYI
WmFUi4u68hWrMSyV64hH1pcoxfW7j62s3YQYoTDWF/aa4D+OOU/3fCcHfbmOmJvVL0TI/kQL7yhB
a+trVbBBlPP1ZIOZXF2j4pXML6Umq/An7NKmQavy1NCBaehFja2Ht3cM+LeMwoblk+5KJ4fjYhA7
Cu7WCRO+QXxzbF+aAnPD4LOzrxVXef4Jg0lxNFWxsFbN72l6mlijdrWXazmDeFCVmB3UIflRk4K7
ZymkO+F8kM0kq/gJ1zrUkex+Q6x8jyMpIQ89csyEpEbkfIIh2ye7nQvJ7oeo8lg8UXpFWgN5w2qq
/LzjDKMZLiiwBL/G1s0v74ua6kCAYzQGGNHdMGAKtXCw8an4EzODVfrRKoNTv8mXCVTUX28/w1+E
F/iVlcYNTqioANB0g5SuP/sezK3i4pjgML8ADMzJjeOq/wifeg46S8UMIQ9NdyQINvJKtXnhrz2A
TqIay3pfRm4E0Gpn3lvqkQGq4TCQ8Md61RxRMuK57CuIywRimHsokHhOr+688i7nAKyEqsj5JzVm
c2VePy78ZGOfSnoua9ZwW+uFKirQY1S6q1MLQoMZrzj/j+97CqCENkOkTfwGv1FKReuFLWwytAfa
+ek7UnqEcCXnk2tC0N8o135EkwwS9Be7gFm0AN2GHtOXhx6TqN5CIAzACsqmHuT7bdx5B7KRbY2W
mOepN9UaQLMmBrwIz1PXLEX79oMLgibH8Ncust9jPG/CeQ59BNVylfu7MvKV4XLDMOUGg4OrMKdj
OX7MP5FqzV9EQ7nq4v+8LKh4iL3ge0ZvKpnWVzDESpJQCM5x+7eS7rgVsFGM+mtFRyFs84kJxXp1
pa022oJtTtjxwjARk1LMYzIkC6SyWutAlsAM6Z4DuftzOGrwx7xidk9ZTk1touOkrU+n7J0o5P/o
MDnIzoDbzIY4Us34giqpuB/5LR6j2iMyN6QZv9HAJfm4sEvgcdS2Waxb2tPyWrDgubfNaerUROg8
+tt+ZesATPuzq0ZVvXJpkzv8wqJmcHEbKAMLcOYFUwxFGcOFlFDS0adU2YYtrYyRebLZqiorZKCF
1h/D/2+N4VWCzybx06QcY1gdS8ZV3MtSwWaCVn/2gt4Ddef0Z7t78eOGXxuwTrVDolMQKkrub+Aa
ktx/J4iX7S1vFrnTTD8QF1OCT5yzq+yyuMeCHPdK0TsY8MBDHUAo0oF5V9yMOPu4HkVb4iXVe7RY
vUQIL9pS17AGC9UHQvbYYb+3IMf1l/jK8wRqEJfPCnG2/k315c3QI4K9X1k6mpZZE87DdTxAAmEL
5ORHqrRnGNQ+KAF8vK4x+tq/YULVsP45aOd0X0yZ7DkM91fRv25bYp1v7+rBtcP4WmcI4l5OBd+E
OscX3Jo/0Nvjx4wVxugP8R5ZmIUWxHyS2tmCcG5IURwdCArx1aKk6rTCvIQqjMkw0s/PMm1dFIEZ
E0V67a8+VFPGqIEzlxMRzYgsMRYJan+ob64SCbcOXhOaHhu2jBai6+xMe5URMrufpNUebMSWAEwK
7xohl4fT1rSZlW+9pgeTcWOiLkxTVPWW55blMuZg0bj5P21Lx3H2xun1CiXrDiSyTR/ei7+SwOvs
9b+lPj8cq+vSqyMvfsPaPiWEk26L+d3fK2PyFNA3qRvNkL6/+9d9bo+IaQyRUxVpp7yUJV3ASMU4
hCxTN/1hOHm2k0BWoM2L2p0AiIuISpGH/m71W8byLKsZs6JNmlaFCuKOV5Bg1PgtpGNX/OjHiWAX
mgm8x0seT8/f5hYv8Sk5glsFRUhYZg23mrHRffZGhzteZuYOtgdkcJn5uhkzNNBj0zpvp8q3L+H9
PA4c+WTDX4x+nXcjJ6d9ZHhVcEet5NhtW2D58M1VNf2mvKs63iPVlOLxgygt3kw1TqhsoD3UPiFU
W8HLlgv8LMyOXgToCQ4jofadrValTCBrwF5J2HnSN/hIvdiVbAnOlY2ERMYCnM9qMw8+/iXuL7i5
3fD076FFy5H4RiTPm6QWxeFC8XztUcqmK2YmrUWQB6AjScCCzKpkbbJ0qE9tRZHixNR/cI/5phGX
HS1v8sEJojaZIWfNtNRDSlDtBsjWtD7h8UwtMnKVqt3K3KSuckn/C7H3OGu3S0CiseVIK73tQiAl
QB9jj9IsJdYyt38kbtPFiOXHBbllVWHfbCCs9v083zZ4IyKckpOIXv0bxQvGhFciEyvC3wL26ktM
oBtVSlFq8KDtxxy0m1SqbTaN4jzEMoaHdi+M5RfOfT8TwF9Urfsovq/mvvqW+UcXHjA2Qxqoen3x
wM3L4JfYH8UIntjJn/7XwABctWk0T9Z5rAcBMs5AvTdk5AJa01Bpd7+vR2dPY3U+zmZLl4Mkvc9C
ITAZxik/ManLscyUKE8kkJVWToXnBSAakfdCZEhyuc7kmnS78pt5rutLNJTaAu/vF6kkwBB7KcrE
JhvSbmV0vNaGdmMZAZ1BPW+AbX+HMOBjoR39a7KNsI/u+eIz4qCyAYhLZn9YDNqOr2BBP9OZQQPu
REw70FfpKc8lnCyv6cQEGp9qChejbc/9WlmcEVqI3BvSHJikt8iI0B/lUc407aKICx2UGqwyviZo
WngI/4iK8aPsDW5o/zOZDMH06l0f8HzjLihqUIjwsIrxmtNWfeUpXC+BnztfobibF5fYKO9gn0y0
VtXm7wwOy95tALFGPc9AeL2pYnpUoxuI0Vt6APKQHGfXkQpFeP6CdDvmYG95fHkHF+clEVAdmQKp
Ly2NHmvGvtJthG5i4Jqt67esrKVcvVXOFSJAhagXVwheKqsFCSXzz6eDNovLzmHFj+EGsMpNvWfs
gE0MrkP9X0U247CwajyEj33NqJkaMjTU/GYoMGsTAvcjb/eHZ6wzBqeBcGpFeon94yeO6Savl5HW
MpP7v7TS8qdoLFaJPuFEPgYCwp5HyCfiIXdY+E4DJ7Rt/Sx5MIYtM4A5260jSyUY7zMOqe5vJS66
1BEG6K07Uzwy8UCLYRPGuX1z0FAWEUzLuxyx2qJfxS7QsPPXH29MRAoLeK2wY5zQ38wH8tCDLi6Q
DP0WdSoNOrKtid8NEgW+RpWo3VhTsbIFlpPJUoiP50ynBiL1ZHNi3GFPcaFSBmciB6zXvEzi59dN
1f02mJQRsxKXOQqmQoIJna4XNZqcvaMEkeamAhR+dxI95cp38UR0iFgAZXCkyaulWGuEb8XJRYrw
Xuq2KroxNxBqmFu60M6AeYZUH77Wg/8jFwbXK3hhTTGKOmJp73a14aLUDfVNFewrx+SQomAyZ9U+
dBuQG/OXsWfkpjeBoFIlB5WgJsB66lo1ouC8AJqy/WLSvfGqxLWXWmcLx7Nw9RcojjZzKosQFaf5
IlPwB1msZKNIhGdhiX2eY6hqqZ3B8dgkjlhM/JLKKsmOsf/ho0EuAdnTTTgKXs3Hczb8QXu3vU5o
ZrJ7RhWd9LvrJg0VR95d89ZVfPjfkL2oKNH/AHqHydxfjEJG5U9thevkVmUJJ3apD7XrGU8DyVBN
YgFDRPtk2hndhCglNABNFFxp2UlA0ot8Vo7a8AIqbFTRBiXFcF3bRqMLtac10nfHCASGaxklaZBH
sCusEnFo6qmSeTAoOmlOtUPj0g4Eu6k69h4sK4E7baCoZ4tFJ7lpYgTanV1bYLwZ+nkdQEmMaetx
43AdBpEgw9hOwnrz60K+OvNo2/qtPG2wj2wHz9pYOBu0scRNbxVDH5u1W3E6+hqLShgLPuiZP+PL
oUNlx3JoCHjzhja7nqlSwEfn1wfT3jXXs2SD8RfeIgvXkxOeGrqfmvF5/FIXNLjndUpheUXk3Zgb
tdslo43t/3pJqs1qYwtoTWeJy0ckqJSR23LB4W5B2RqGzGtbTKY20EgUzkzhyL6ypH0DXrsdEJ82
M05I6XAPXWXSIHNznjSR4SnQ0oLhjLhsGOFRMR9SDGh0vcxFct0jYMSvqKHIdXHySj34DTDvbTeU
zO+gSlFiWpcjIG2Gu5BSUPkGOIeZNO89TZmzLWVpSs5AILw98QdG+2UPGuK6u1zm9xu3dMFjdYMa
Xx/229taeChDQIQIXtUHMyFoUEM9WUYlvB0765AGRWql5gbjSpqO6uiLsi51dgyrJr03O/kjSn1B
qy0ijNicWgjjRQRK03AI6Ow2P6oRvmZB2HL/1zL3TZXMQhGlnUoqhx2/JiebM5bZKEZg1ofep5dr
DsUya3ZrXFBhvXvgMDiBseC7gmg6iNu50w/Ndh36cypMUHkBOpPrPXtNT5HntSi8VbSBiqEh2FuE
IXl8xti/Qr/JRJ4xpc6QCS8AKUYoKifQo2RNvHAfSRXpGmj5ZCq8KlRQkLfL6RQZKYSvcuvGLkmz
3Nb2xVOASVOofoQw7R5Of3EwkxOsTWoTKVCJx8fa6EzXdjT3KebsFDQYW0ky/E3ArtG2iRoAcxQ+
vDzmEzs+Rq6Ac2w9mYg5yRSjRAkGW05x+hyHsA4dQF5aJ9Rcrd6MBOdcwWVdeWO5UZkingr+UEpi
ItFps3akmdHX8aYyvqxYFNTa7zhdelEGB8QZRSG8U51lpTy2sf1zaoqOY2V0j6RLle2mN3Nxya9k
IS/m9OF5RFE4fUWPReLWmd811gMRmA2vwO2rlPexDD/IivKc9pybmCamuaTWWN1jqWYq17E+IjH7
5kr3alZAJCtDOuQ36BGzAIRw15aZp4N6HANIBRiY0QL3jfCSetiI/cCW1hdWR1wCuwAQW4dTBtVP
SioKnDov4mpxGYlujnXAL3BznZ1etdz+FjCeyDhGyfelgLTZHdQE5XtqXYzIJ9yR27pf7dUzS5Mk
oqJh4gBAXE96ByhqB4zi7RxsIwzqkVcfyrkCrjmBm+909vvfyfpVOTmn4rHoiOlRF7ytctUdSg2L
chGN/xuuJs2OfphO7n3LqKQ/xOYgBMTNi6nE6JpChBSzO2eGgtxbAHx8/CYnVOb9miT0/7/1azs2
iDGf2CevaIYhqKkJ7arKnkVVxGqYQyvBqVHWmqh5dNmyHUxAa18P9g9NmPlb351GAQF5YeKYzhj+
dCyjrCSbrmTVcF82BDpXgT2zBfUjShQU7bZb3GbafERlElD7rSZsdQ9Vcf+7Few5EnXF/CA1zKBN
4JqaI9R0F9A9cl2LcAfhAdutm02pug+YNeo1+IlY2Z77+E3WsV1aAnGtn7NYRzy11E7OtPh5ncJ6
JKadALugyiAiM+Qu4FbcnNWxA6PMX9wZrR/AbIgNvPNBIxEMl8jRk57naAIhF3CnyfQw2KBlluFa
a0aZHSI2Pt4RSrUH8iF4K8dr/X4gqlI6KiOueEaJRqdh6v/CgPhhSUmr0FJQwWWMIC9xw74RfHNg
B0xJ2e+WY7BXSb4MxdE9NIGEe1p7Xvcsgt7FGX1QoQJIVvWbtNJue84voMqrxR+oTTJqA/Ar8mgq
aZ2dX1GY4pK7TgDUowOpfJ+1u+OS/YIBj0mhUVLL3OTgB4xx5X+NZQuDxrGJEL6KbCZvsTbDDyy6
a5rDL5mRxMAVTFRdaMQd8MZBr1LCxffqNisI4buI6JbpZfCuMzV4P8ZdhuNaoH8cxh2T6w1PBYVZ
4+i3wKjbe8UsTKLK+QEZ3fJYLob5Bs5JvhCVfQlAfOSp1XUBUu+3VAVWbN2kNzerBGQcDOXT7aiX
kZXc9xxn+R9Gg089vlw8XUqsIBZkjU/zlVvdYZzurJc47tB6LpjTX31WfQkeN2EN8n2Lsu+c8Ufm
5g3GOtqeYT+TX1HbpVAOnZOl3menER1+a6/WMBRyURwVzluEHRpMLoY8un9uXhUhRma2G3WuhdZw
m9Kpi0oKY704TVxBfyLU5PLDxOJJF63T1Nqq6bNBs9FTsp4C2QZ+M4BO9Ainmcsuq4Mr6UPcrU6u
eRZBsZcnfh4UYuqPw18p4VXOnh4Z6tBNEAOD17OQ8CoBJ/kK3aONdy2QLPHjxzIo7MFIgAiFctPV
y8hvNBy3EM8pFQrY/CCSGpWO0fdO+qH490Dx7jUsF8zpvI2k1eUO3rSmZcvvLJLRQak+cbmTgX0+
x+Cbc4VOr9032aOoYwLpocRXPTLN+Z3L/47giptAUdbBqc0GgBa6L5xMkcjiw0ybJrWbOwtuV74K
HATXXmbjvRpFSly9XBtK9LmdqrknMxs8SOEj0y4lxUWYZu1dcgkbUxEFtjWu+lRthBTCA90EXms/
3gf5fB5ePPAg7ZPuHUq3HnE/DqUVXe1bRwtfVgaJ0QeCNmlqyez6RiK5ncH3lAk73UQJIzBQTPo/
1Q8dgUUspasQSInoteYN/7SkdOXL4TKm9VuEuWr6Z+ElICIPvifGPRN9rzqGbEY85mkQRu1O/tMs
E6EkTpWReObfa0X829Y7r8KljwvSnJ9KDRCiwututnhLHc5Tbu9g44UsltbYjqIbwHDBWKuGPxAX
CdGWOT70oziXeX8BsWqt+Buafby56opTHbtjQZc/x5y0DeKnUlDhwKbCLHspzxPtuK4jzi3yxkMa
ahtd9VLwKG/C3S1Gf5G2GQYQxkOwTftbP4EeIBTonzSGWqvCfwziueBzAatRWs4qD8t/YbkUW0qo
Sp0pAkS4fqBhyzAJfLvYqVFoNyVThKilC/dhcEYnvVQr3fGhTd/y3Sj1cZ6w1yVnKNeViurfSMik
mJSZwcsBAPueR31vbwIrXch5TxFnuujixubYx5pfQte70AfaZjxq+8BK7MK6Hro8p/XuI9kJ3tpA
RgbGw+DcWI1r6eWfkTidOS74cVcQN7O1Qaj3vggHY1vxHTU8+ujHfSMJkIE20JIh1qfln2siviox
w8EZgwJ9+rJNgU004SqrixGGMR8k+cJ4ygZ7S5AzpMlpzpgzTmVOmgng+SzKJRloCmh6jnA15+f+
VkL/o62CYl2CmrUZVT3QMk1DAI4r9hlF3KfoYFh43Qo9sRYvq3m5RVV3lDU542Czww8aYuAdlEDx
wZzm759U9wSWQW0DU30Z5Q0qet0V8wJAREDK9nkz0wMgYD2z9HwF2erGnXf4u5M+u9NU0UBruZTx
EOcNCFLSUicIXy372csq55+ReWtYS991NBFfL+dy5YZX0YZiMiXv+VPTrpTTAbq7TBLSQ5ggLTsu
DU6+RKIp05wqMXgMHN2FmJFrDPjPie34x/1OqaG5QYiJoPKZaYILRPNAdrV4uzcx/U+fptCYG9wl
JJrAJJbuIQ08GYfX+u1vy6UUOaSMoN6k3ViPlxAtUsOJket71srFDHt1LrooomLzI6eNqykUr6Wz
kbaY+C3uEitmiG57ItEP+NQo8KU90cqtY8GPb9SNgnzr20HzYJmZJtbZaSZjdHtJTPU9GBBLBa+u
2+mIp9NR11/Np6eVDHTroeiKKqkejmwn64uysnM0wTYMymeGOUcQcxFZppzQJg8QemIOCe0olwqD
gL5t4ux2mDFjBfAJF0plBcnBUo1yB9yAaRDGDBA20HdZwSwKeE3IHqYRQXxJE1UgcS4lQG8O8iVS
ywsbAvyzlyRRK08FIbrMmXGLG+LZklDYZDUCVC8ZaKOoZvPSnxgT9kj56EpEv92YQ3wgmhkvXKkU
tGNB/NcIQKlWp9DZmx58KUeujmYdmlAyjFd4DyQW/1Nyn+HhGPa8c8asK+1J+/2wP1z7cM7zMNET
rJsru6oDVtunumLp/iVhUitFDR0hVfsU24ZVt5HjPQTP0C83Ks0rpl9A7lUT0w4HI7muWR4yVszM
NivDZLnckcJPoXiE+KFdkC1zHkCr/zf8dkva2hem296NwifqLZBNmA1I2pE3UDYgJw33NIQ7leBy
uNV0tz0osC/JZBwUBPgr1B/IXU3KOV2oW33dQ+/IEFfr0G1KEWy2hTejmqBVB3LKclXkD4pdFwVV
y75R5gSuqD19KwsqAGWogvKcErCC7GbTLVEmao2/wYVV5tY4xffnzASzPSx9V6YFtLxmJotZ2JQT
v9TmpjldpcJX6vaLjQ0cKu3yNJ21TTe1fl2QXdNRkDnX8wHqpdXc3XHVh9SWLY67N4MtkVErVTP2
fYmoPh2Qv3XKt7iVt3F0mCNqR6FYAO1N1igNdTTEZy6rNxfGiFVAh4fne2N7R0L2C9ykJPtRPQ+W
L9CSLZdlEgn/om4inCF6+PPfiIJIQQx4g0+/BtF4d2kCd5wJscAWWbi5mWCnVwFMC3EfJ5EnKEtx
VjmD1OX8byt6i9dFEtmS45qe1h79qKx1aEnzJsA4mculngnkGiZJgApVbx0N6W/tuFv1fx1q3JDx
9ORja+frRF2UJRLl8e6uisY65+dbXpmWDn8dNE8J/mkJkuSQRbEcaA2V0k/Tfr/P6rTyvo2udfb2
8Lc1tikeBegy9OSaCPn/FFJoCoW7SORmWZ4Rs4IyqFkYD7JL4xPTk9XDURcoAo0yq0P3+NKFePjo
8MUXhGE8hXOnYIE1uJ+w1PZF5okN5ylSUQEAuou/IlojYqJiNHQFuuvSqvqq04eMzuwUansWPv0T
ejZw3gNPKgY8cfG8BjM/r2GbgJuFBM31zhjuzJmqG1iO57k7XfBWHURJ7zQ3p+b8kMHlyok8PrxW
IvtTXfiPLiGJ+4eBdEUFFQqSd2YDEWdN3M8KdL0FYP8uqTeqbK8LfSxdZE2ak9upyooipi5cP+O6
db7R2KCTAmWIDcAus3sFuZ2PZKnlpI0kCXXzVDauSCTdTL9Nm7D2VjXxYLE30XOXvxBqQ1rWKRXG
OohdpyR8AizKkrV9WsKMCxYxlJ+BYzYWBkmJUbPPL3sD2On4TFjJkd9tIdIS3xQBrjx0yshxPm2d
xpxgtinJi5bvJZUNeRhW5V7+dsCVedbJcZNr8RHw66lsEYYHoCJthH2yOcWLMixYFAzKRaIOXDYh
mKMXfgWw89Nixjb8DpYdYpz2fKRbIp4P+Omp/w+Z3YfEuown9NwMzZjW9fq0qhx9bQLDI87h1tOi
Ej8IGEkz42auwXbIGOh92XmV2e25IpKvuHMVGScDbBg37JhiuVo9htkhVGQClx8e+p5CPJ6E3dt5
Bw9XmG3fnoNCE3VldOCpmmk6rsJZ6jZV8S+Sqsm994glp0z4r61hQmx2Ank5xS5aVR8CxbT1JU+k
GKjZEOIW0QW48DjoFgONzWXdzk/xr+2Cy27sbXONp5jpwLMloW/FFchoEFo5kAcp07XDQfB+PkJr
YyXT+zNQ5u0fbq0cbm1YkjTzlKRnww6Y9Ik3Alzw/+yMG6R7jyxVdShIUDkmk3fy6nc/o3E5pPrF
2aDm5TIaobSYliOJkMMNz6IaLgngvH3S9s8Cx09bKpg9Xqlq4mEUO8/E9rL8f92j4IgGYbwPxOhQ
cI1Kh1dj5pFK0DAT7rniK4BUOOndKXiKR2Y0zpfUp0v1PNWkLOg6Q78VOCwVFQE3ri34BRrfOE2p
I9NCwgjbYa4SYXPhExySHRZeh5eKqMsYF0Dq3LEnsoawPgYMbJ7S1U1uSIm88Uhpiyn88hGhclnL
g8bcbDxncGfaB56QSQuTiOMWCWfpTXpM4Ti4ySnjP582rMQt4Lhm0Y70svvdb+J9p0/qUNPo+GQT
DpVtKv8wO9IZpBKnYt58XTufdww7pkLFHdzA9gyrH6/XNZlGppQ7bBQjYXlrp7AioiRKBtd5F/Gm
BZZ38ZNoa8BuKmpFIhkHGREFHD9Cw7PKDJXHARJsr9qUN5godqDjQJyx1NncVQYStdmuqJkG8GH6
f6bnKgAqqCfGYr2mAIWyy4lno/PIu7+a5CPxjZ1Uqiaa/urABHD0NUe+dGCxdnMVEskk+Xf8By2d
W18f5VLfYY0N/bPlv3/hI8MdCnhsgF0OJyudkdwLf975jLHSjXuheSPCcGLp2s7rvOmmTUKQDDqv
kP95TlsJbCCtDH9BnQdrjUB+Tn2D2emewgHDkulk
`pragma protect end_protected
