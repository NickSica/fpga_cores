//wire gt_refclk0;
wire  q1_altclk_m;
wire [31:0] q1_apb3prdata_m;
wire  q1_apb3pready_m;
wire  q1_apb3pslverr_m;
wire [15:0] q1_apb3paddr_m;
wire  q1_apb3clk_m;
wire q1_axisclk_m;
wire  q1_apb3penable_m;
wire  q1_apb3presetn_m;
wire  q1_apb3psel_m;
wire [31:0] q1_apb3pwdata_m;
wire  q1_apb3pwrite_m;
wire  q1_bgbypassb_m;
wire  q1_bgmonitorenb_m;
wire  q1_bgpdb_m;
wire  q1_bgrcalovrdenb_m;
wire [4:0] q1_bgrcalovrd_m;
wire  q1_scanclkb_m;
wire  q1_scancntrlin_m;
wire  q1_scanenb_m;
wire [3:0] q1_scanin_m;
wire  q1_scanrstb_m;
wire  q1_xpscanclk_m;
wire  q1_xpscanenb_m;
wire [15:0] q1_xpscanin_m;
wire  q1_xpscanmodeb_m;
wire  q1_xpscanrstb_m;
wire  q1_cssdrstb_m;
wire  q1_cssdstopclk_m;
wire  q1_edtupdateb_m;
wire  ch4_txoutclk_m;
wire  ch4_rxoutclk_m;
wire  ch4_bufgtce_m;
wire [3:0] ch4_bufgtcemask_m;
wire [11:0] ch4_bufgtdiv_m;
wire  ch4_bufgtrst_m;
wire [3:0] ch4_bufgtrstmask_m;
wire [31:0] ch4_dmonitorout_m;
wire  ch4_eyescandataerror_m;
wire  ch4_iloresetdone_m;
wire [15:0] ch4_pcsrsvdout_m;
wire [15:0] ch4_pinrsvdas_m;
wire  ch4_phyready_m;
wire  ch4_phystatus_m;
wire  ch4_resetexception_m;
wire [7:0] ch4_rx10gstat_m;
wire [2:0] ch4_rxbufstatus_m;
wire  ch4_rxbyteisaligned_m;
wire  ch4_rxbyterealign_m;
wire  ch4_rxcdrlock_m;
wire  ch4_rxcdrphdone_m;
wire  ch4_rxchanbondseq_m;
wire  ch4_rxchanisaligned_m;
wire  ch4_rxchanrealign_m;
wire [4:0] ch4_rxchbondo_m;
wire [1:0] ch4_rxclkcorcnt_m;
wire  ch4_rxcominitdet_m;
wire  ch4_rxcommadet_m;
wire  ch4_rxcomsasdet_m;
wire  ch4_rxcomwakedet_m;
wire [15:0] ch4_rxctrl0_m;
wire [15:0] ch4_rxctrl1_m;
wire [7:0] ch4_rxctrl2_m;
wire [7:0] ch4_rxctrl3_m;
wire [127:0] ch4_rxdata_m;
wire [7:0] ch4_rxdataextendrsvd_m;
wire [1:0] ch4_rxdatavalid_m;
wire  ch4_rxdccdone_m;
wire  ch4_rxdlyalignerr_m;
wire  ch4_rxdlyalignprog_m;
wire  ch4_rxelecidle_m;
wire  ch4_rxfinealigndone_m;
wire [5:0] ch4_rxheader_m;
wire [1:0] ch4_rxheadervalid_m;
wire  ch4_rxosintdone_m;
wire  ch4_rxosintstarted_m;
wire  ch4_rxosintstrobedone_m;
wire  ch4_rxosintstrobestarted_m;
wire  ch4_rxphaligndone_m;
wire  ch4_rxphalignerr_m;
wire  ch4_rxphdlyresetdone_m;
wire  ch4_rxphsetinitdone_m;
wire  ch4_rxphshift180done_m;
wire  ch4_rxpmaresetdone_m;
wire  ch4_rxprbserr_m;
wire  ch4_rxprbslocked_m;
wire  ch4_rxresetdone_m;
wire  ch4_rxsliderdy_m;
wire [1:0] ch4_rxstartofseq_m;
wire [2:0] ch4_rxstatus_m;
wire  ch4_rxsyncdone_m;
wire  ch4_rxvalid_m;


wire  ch4_tstclk0_m  ;
wire  ch4_tstclk1_m  ;
wire  ch5_tstclk0_m  ;
wire  ch5_tstclk1_m  ;
wire  ch6_tstclk0_m  ;
wire  ch6_tstclk1_m  ;
wire  ch7_tstclk0_m  ;
wire  ch7_tstclk1_m  ;





wire  ch4_tx10gstat_m;
wire [1:0] ch4_txbufstatus_m;
wire  ch4_txcomfinish_m;
wire  ch4_txdccdone_m;
wire  ch4_txdlyalignerr_m;
wire  ch4_txdlyalignprog_m;
wire  ch4_txphaligndone_m;
wire  ch4_txphalignerr_m;
wire  ch4_txphalignoutrsvd_m;
wire  ch4_txphdlyresetdone_m;
wire  ch4_txphshift180done_m;
wire  ch4_txpmaresetdone_m;
wire  ch4_txresetdone_m;
wire  ch4_txsyncdone_m;
wire  ch4_cdrbmcdrreq_m;
wire  ch4_cdrfreqos_m;
wire  ch4_cdrincpctrl_m;
wire  ch4_cdrstepdir_m;
wire  ch4_cdrstepsq_m;
wire  ch4_cdrstepsx_m;
wire  ch4_clkrsvd0_m;
wire  ch4_clkrsvd1_m;
wire  ch4_cssdrstb_m;
wire  ch4_cssdstopclk_m;
wire  ch4_edtupdateb_m;
wire  ch4_dmonfiforeset_m;
wire  ch4_dmonitorclk_m;
wire  ch4_eyescanreset_m;
wire  ch4_eyescantrigger_m;
wire [15:0] ch4_gtrsvd_m;
wire  ch4_gtrxreset_m;
wire  ch4_gttxreset_m;
wire  ch4_hsdppcsreset_m;
wire  ch4_iloreset_m;
wire  ch4_iloresetmask_m;
wire [2:0] ch4_loopback_m;
wire  ch4_pcierstb_m;
wire [15:0] ch4_pcsrsvdin_m;
wire  ch4_phyesmadaptsave_m;
wire  ch4_rxcdrhold_m;
wire  ch4_rxcdrovrden_m;
wire  ch4_rxcdrreset_m;
wire [4:0] ch4_rxchbondi_m;
wire  ch4_rxdapicodeovrden_m;
wire  ch4_rxdapicodereset_m;
wire  ch4_rxdlyalignreq_m;
wire  ch4_rxeqtraining_m;
wire  ch4_rxgearboxslip_m;
wire  ch4_rxlatclk_m;
wire  ch4_rxlpmen_m;
wire  ch4_rxmldchaindone_m;
wire  ch4_rxmldchainreq_m;
wire  ch4_rxmlfinealignreq_m;
wire  ch4_rxoobreset_m;
wire [4:0] ch4_rxpcsresetmask_m;
wire [1:0] ch4_rxpd_m;
wire  ch4_rxphalignreq_m;
wire [1:0] ch4_rxphalignresetmask_m;
wire  ch4_rxphdlypd_m;
wire  ch4_rxphdlyreset_m;
wire  ch4_rxphsetinitreq_m;
wire  ch4_rxphshift180_m;
wire [6:0] ch4_rxpmaresetmask_m;
wire  ch4_rxpolarity_m;
wire  ch4_rxprbscntreset_m;
wire [3:0] ch4_rxprbssel_m;
wire  ch4_rxprogdivreset_m;
wire [7:0] ch4_rxrate_m;
wire [1:0] ch4_rxresetmode_m;
wire  ch4_rxslide_m;
wire  ch4_rxsyncallin_m;
wire  ch4_rxtermination_m;
wire  ch4_rxuserrdy_m;
wire  ch4_rxusrclk_m;
wire [19:0] ch4_tstin_m;
wire  ch4_txcominit_m;
wire  ch4_txcomsas_m;
wire  ch4_txcomwake_m;
wire [15:0] ch4_txctrl0_m;
wire [15:0] ch4_txctrl1_m;
wire [7:0] ch4_txctrl2_m;
wire  ch4_txdapicodeovrden_m;
wire  ch4_txdapicodereset_m;
wire [127:0] ch4_txdata_m;
wire [7:0] ch4_txdataextendrsvd_m;
wire [1:0] ch4_txdeemph_m;
wire  ch4_txdetectrx_m;
wire [4:0] ch4_txdiffctrl_m;
wire  ch4_txdlyalignreq_m;
wire  ch4_txelecidle_m;
wire [5:0] ch4_txheader_m;
wire  ch4_txinhibit_m;
wire  ch4_txlatclk_m;
wire [6:0] ch4_txmaincursor_m;
wire [2:0] ch4_txmargin_m;
wire  ch4_txmldchaindone_m;
wire  ch4_txmldchainreq_m;
wire  ch4_txoneszeros_m;
wire  ch4_txpausedelayalign_m;
wire  ch4_txpcsresetmask_m;
wire [1:0] ch4_txpd_m;
wire  ch4_txphalignreq_m;
wire [1:0] ch4_txphalignresetmask_m;
wire  ch4_txphdlypd_m;
wire  ch4_txphdlyreset_m;
wire  ch4_txphdlytstclk_m;
wire  ch4_txphsetinitreq_m;
wire  ch4_txphshift180_m;
wire  ch4_txpicodeovrden_m;
wire  ch4_txpicodereset_m;
wire  ch4_txpippmen_m;
wire [4:0] ch4_txpippmstepsize_m;
wire  ch4_txpisopd_m;
wire [2:0] ch4_txpmaresetmask_m;
wire  ch4_txpolarity_m;
wire [4:0] ch4_txpostcursor_m;
wire  ch4_txprbsforceerr_m;
wire [3:0] ch4_txprbssel_m;
wire [4:0] ch4_txprecursor_m;
wire  ch4_txprogdivreset_m;
wire [7:0] ch4_txrate_m;
wire [1:0] ch4_txresetmode_m;
wire [6:0] ch4_txsequence_m;
wire  ch4_txswing_m;
wire  ch4_txsyncallin_m;
wire  ch4_txuserrdy_m;
wire  ch4_txusrclk_m;
wire  ch4_scanclkb_m;
wire  ch4_scancntrlin_m;
wire  ch4_scanenb_m;
wire [3:0] ch4_scanin_m;
wire  ch4_scanrstb_m;

wire  ch5_bufgtce_m;
wire [3:0] ch5_bufgtcemask_m;
wire [11:0] ch5_bufgtdiv_m;
wire  ch5_bufgtrst_m;
wire [3:0] ch5_bufgtrstmask_m;
wire [31:0] ch5_dmonitorout_m;
wire  ch5_eyescandataerror_m;
wire  ch5_iloresetdone_m;
wire [15:0] ch5_pcsrsvdout_m;
wire [15:0] ch5_pinrsvdas_m;
wire  ch5_phyready_m;
wire  ch5_phystatus_m;
wire  ch5_resetexception_m;
wire [7:0] ch5_rx10gstat_m;
wire [2:0] ch5_rxbufstatus_m;
wire  ch5_rxbyteisaligned_m;
wire  ch5_rxbyterealign_m;
wire  ch5_rxcdrlock_m;
wire  ch5_rxcdrphdone_m;
wire  ch5_rxchanbondseq_m;
wire  ch5_rxchanisaligned_m;
wire  ch5_rxchanrealign_m;
wire [4:0] ch5_rxchbondo_m;
wire [1:0] ch5_rxclkcorcnt_m;
wire  ch5_rxcominitdet_m;
wire  ch5_rxcommadet_m;
wire  ch5_rxcomsasdet_m;
wire  ch5_rxcomwakedet_m;
wire [15:0] ch5_rxctrl0_m;
wire [15:0] ch5_rxctrl1_m;
wire [7:0] ch5_rxctrl2_m;
wire [7:0] ch5_rxctrl3_m;
wire [127:0] ch5_rxdata_m;
wire [7:0] ch5_rxdataextendrsvd_m;
wire [1:0] ch5_rxdatavalid_m;
wire  ch5_rxdccdone_m;
wire  ch5_rxdlyalignerr_m;
wire  ch5_rxdlyalignprog_m;
wire  ch5_rxelecidle_m;
wire  ch5_rxfinealigndone_m;
wire [5:0] ch5_rxheader_m;
wire [1:0] ch5_rxheadervalid_m;
wire  ch5_rxosintdone_m;
wire  ch5_rxosintstarted_m;
wire  ch5_rxosintstrobedone_m;
wire  ch5_rxosintstrobestarted_m;
wire  ch5_rxphaligndone_m;
wire  ch5_rxphalignerr_m;
wire  ch5_rxphdlyresetdone_m;
wire  ch5_rxphsetinitdone_m;
wire  ch5_rxphshift180done_m;
wire  ch5_rxpmaresetdone_m;
wire  ch5_rxprbserr_m;
wire  ch5_rxprbslocked_m;
wire  ch5_rxresetdone_m;
wire  ch5_rxsliderdy_m;
wire [1:0] ch5_rxstartofseq_m;
wire [2:0] ch5_rxstatus_m;
wire  ch5_rxsyncdone_m;
wire  ch5_rxvalid_m;
wire  ch5_tx10gstat_m;
wire [1:0] ch5_txbufstatus_m;
wire  ch5_txcomfinish_m;
wire  ch5_txdccdone_m;
wire  ch5_txdlyalignerr_m;
wire  ch5_txdlyalignprog_m;
wire  ch5_txphaligndone_m;
wire  ch5_txphalignerr_m;
wire  ch5_txphalignoutrsvd_m;
wire  ch5_txphdlyresetdone_m;
wire  ch5_txphshift180done_m;
wire  ch5_txpmaresetdone_m;
wire  ch5_txresetdone_m;
wire  ch5_txsyncdone_m;
wire  ch5_cdrbmcdrreq_m;
wire  ch5_cdrfreqos_m;
wire  ch5_cdrincpctrl_m;
wire  ch5_cdrstepdir_m;
wire  ch5_cdrstepsq_m;
wire  ch5_cdrstepsx_m;
wire  ch5_clkrsvd0_m;
wire  ch5_clkrsvd1_m;
wire  ch5_cssdrstb_m;
wire  ch5_cssdstopclk_m;
wire  ch5_edtupdateb_m;
wire  ch5_dmonfiforeset_m;
wire  ch5_dmonitorclk_m;
wire  ch5_eyescanreset_m;
wire  ch5_eyescantrigger_m;
wire [15:0] ch5_gtrsvd_m;
wire  ch5_gtrxreset_m;
wire  ch5_gttxreset_m;
wire  ch5_hsdppcsreset_m;
wire  ch5_iloreset_m;
wire  ch5_iloresetmask_m;
wire [2:0] ch5_loopback_m;
wire  ch5_pcierstb_m;
wire [15:0] ch5_pcsrsvdin_m;
wire  ch5_phyesmadaptsave_m;
wire  ch5_rxcdrhold_m;
wire  ch5_rxcdrovrden_m;
wire  ch5_rxcdrreset_m;
wire [4:0] ch5_rxchbondi_m;
wire  ch5_rxdapicodeovrden_m;
wire  ch5_rxdapicodereset_m;
wire  ch5_rxdlyalignreq_m;
wire  ch5_rxeqtraining_m;
wire  ch5_rxgearboxslip_m;
wire  ch5_rxlatclk_m;
wire  ch5_rxlpmen_m;
wire  ch5_rxmldchaindone_m;
wire  ch5_rxmldchainreq_m;
wire  ch5_rxmlfinealignreq_m;
wire  ch5_rxoobreset_m;
wire [4:0] ch5_rxpcsresetmask_m;
wire [1:0] ch5_rxpd_m;
wire  ch5_rxphalignreq_m;
wire [1:0] ch5_rxphalignresetmask_m;
wire  ch5_rxphdlypd_m;
wire  ch5_rxphdlyreset_m;
wire  ch5_rxphsetinitreq_m;
wire  ch5_rxphshift180_m;
wire [6:0] ch5_rxpmaresetmask_m;
wire  ch5_rxpolarity_m;
wire  ch5_rxprbscntreset_m;
wire [3:0] ch5_rxprbssel_m;
wire  ch5_rxprogdivreset_m;
wire [7:0] ch5_rxrate_m;
wire [1:0] ch5_rxresetmode_m;
wire  ch5_rxslide_m;
wire  ch5_rxsyncallin_m;
wire  ch5_rxtermination_m;
wire  ch5_rxuserrdy_m;
wire  ch5_rxusrclk_m;
wire [19:0] ch5_tstin_m;
wire  ch5_txcominit_m;
wire  ch5_txcomsas_m;
wire  ch5_txcomwake_m;
wire [15:0] ch5_txctrl0_m;
wire [15:0] ch5_txctrl1_m;
wire [7:0] ch5_txctrl2_m;
wire  ch5_txdapicodeovrden_m;
wire  ch5_txdapicodereset_m;
wire [127:0] ch5_txdata_m;
wire [7:0] ch5_txdataextendrsvd_m;
wire [1:0] ch5_txdeemph_m;
wire  ch5_txdetectrx_m;
wire [4:0] ch5_txdiffctrl_m;
wire  ch5_txdlyalignreq_m;
wire  ch5_txelecidle_m;
wire [5:0] ch5_txheader_m;
wire  ch5_txinhibit_m;
wire  ch5_txlatclk_m;
wire [6:0] ch5_txmaincursor_m;
wire [2:0] ch5_txmargin_m;
wire  ch5_txmldchaindone_m;
wire  ch5_txmldchainreq_m;
wire  ch5_txoneszeros_m;
wire  ch5_txpausedelayalign_m;
wire  ch5_txpcsresetmask_m;
wire [1:0] ch5_txpd_m;
wire  ch5_txphalignreq_m;
wire [1:0] ch5_txphalignresetmask_m;
wire  ch5_txphdlypd_m;
wire  ch5_txphdlyreset_m;
wire  ch5_txphdlytstclk_m;
wire  ch5_txphsetinitreq_m;
wire  ch5_txphshift180_m;
wire  ch5_txpicodeovrden_m;
wire  ch5_txpicodereset_m;
wire  ch5_txpippmen_m;
wire [4:0] ch5_txpippmstepsize_m;
wire  ch5_txpisopd_m;
wire [2:0] ch5_txpmaresetmask_m;
wire  ch5_txpolarity_m;
wire [4:0] ch5_txpostcursor_m;
wire  ch5_txprbsforceerr_m;
wire [3:0] ch5_txprbssel_m;
wire [4:0] ch5_txprecursor_m;
wire  ch5_txprogdivreset_m;
wire [7:0] ch5_txrate_m;
wire [1:0] ch5_txresetmode_m;
wire [6:0] ch5_txsequence_m;
wire  ch5_txswing_m;
wire  ch5_txsyncallin_m;
wire  ch5_txuserrdy_m;
wire  ch5_txusrclk_m;
wire  ch5_scanclkb_m;
wire  ch5_scancntrlin_m;
wire  ch5_scanenb_m;
wire [3:0] ch5_scanin_m;
wire  ch5_scanrstb_m;

wire  ch6_bufgtce_m;
wire [3:0] ch6_bufgtcemask_m;
wire [11:0] ch6_bufgtdiv_m;
wire  ch6_bufgtrst_m;
wire [3:0] ch6_bufgtrstmask_m;
wire [31:0] ch6_dmonitorout_m;
wire  ch6_eyescandataerror_m;
wire  ch6_iloresetdone_m;
wire [15:0] ch6_pcsrsvdout_m;
wire [15:0] ch6_pinrsvdas_m;
wire  ch6_phyready_m;
wire  ch6_phystatus_m;
wire  ch6_resetexception_m;
wire [7:0] ch6_rx10gstat_m;
wire [2:0] ch6_rxbufstatus_m;
wire  ch6_rxbyteisaligned_m;
wire  ch6_rxbyterealign_m;
wire  ch6_rxcdrlock_m;
wire  ch6_rxcdrphdone_m;
wire  ch6_rxchanbondseq_m;
wire  ch6_rxchanisaligned_m;
wire  ch6_rxchanrealign_m;
wire [4:0] ch6_rxchbondo_m;
wire [1:0] ch6_rxclkcorcnt_m;
wire  ch6_rxcominitdet_m;
wire  ch6_rxcommadet_m;
wire  ch6_rxcomsasdet_m;
wire  ch6_rxcomwakedet_m;
wire [15:0] ch6_rxctrl0_m;
wire [15:0] ch6_rxctrl1_m;
wire [7:0] ch6_rxctrl2_m;
wire [7:0] ch6_rxctrl3_m;
wire [127:0] ch6_rxdata_m;
wire [7:0] ch6_rxdataextendrsvd_m;
wire [1:0] ch6_rxdatavalid_m;
wire  ch6_rxdccdone_m;
wire  ch6_rxdlyalignerr_m;
wire  ch6_rxdlyalignprog_m;
wire  ch6_rxelecidle_m;
wire  ch6_rxfinealigndone_m;
wire [5:0] ch6_rxheader_m;
wire [1:0] ch6_rxheadervalid_m;
wire  ch6_rxosintdone_m;
wire  ch6_rxosintstarted_m;
wire  ch6_rxosintstrobedone_m;
wire  ch6_rxosintstrobestarted_m;
wire  ch6_rxphaligndone_m;
wire  ch6_rxphalignerr_m;
wire  ch6_rxphdlyresetdone_m;
wire  ch6_rxphsetinitdone_m;
wire  ch6_rxphshift180done_m;
wire  ch6_rxpmaresetdone_m;
wire  ch6_rxprbserr_m;
wire  ch6_rxprbslocked_m;
wire  ch6_rxresetdone_m;
wire  ch6_rxsliderdy_m;
wire [1:0] ch6_rxstartofseq_m;
wire [2:0] ch6_rxstatus_m;
wire  ch6_rxsyncdone_m;
wire  ch6_rxvalid_m;
wire  ch6_tx10gstat_m;
wire [1:0] ch6_txbufstatus_m;
wire  ch6_txcomfinish_m;
wire  ch6_txdccdone_m;
wire  ch6_txdlyalignerr_m;
wire  ch6_txdlyalignprog_m;
wire  ch6_txphaligndone_m;
wire  ch6_txphalignerr_m;
wire  ch6_txphalignoutrsvd_m;
wire  ch6_txphdlyresetdone_m;
wire  ch6_txphshift180done_m;
wire  ch6_txpmaresetdone_m;
wire  ch6_txresetdone_m;
wire  ch6_txsyncdone_m;
wire  ch6_cdrbmcdrreq_m;
wire  ch6_cdrfreqos_m;
wire  ch6_cdrincpctrl_m;
wire  ch6_cdrstepdir_m;
wire  ch6_cdrstepsq_m;
wire  ch6_cdrstepsx_m;
wire  ch6_clkrsvd0_m;
wire  ch6_clkrsvd1_m;
wire  ch6_cssdrstb_m;
wire  ch6_cssdstopclk_m;
wire  ch6_edtupdateb_m;
wire  ch6_dmonfiforeset_m;
wire  ch6_dmonitorclk_m;
wire  ch6_eyescanreset_m;
wire  ch6_eyescantrigger_m;
wire [15:0] ch6_gtrsvd_m;
wire  ch6_gtrxreset_m;
wire  ch6_gttxreset_m;
wire  ch6_hsdppcsreset_m;
wire  ch6_iloreset_m;
wire  ch6_iloresetmask_m;
wire [2:0] ch6_loopback_m;
wire  ch6_pcierstb_m;
wire [15:0] ch6_pcsrsvdin_m;
wire  ch6_phyesmadaptsave_m;
wire  ch6_rxcdrhold_m;
wire  ch6_rxcdrovrden_m;
wire  ch6_rxcdrreset_m;
wire [4:0] ch6_rxchbondi_m;
wire  ch6_rxdapicodeovrden_m;
wire  ch6_rxdapicodereset_m;
wire  ch6_rxdlyalignreq_m;
wire  ch6_rxeqtraining_m;
wire  ch6_rxgearboxslip_m;
wire  ch6_rxlatclk_m;
wire  ch6_rxlpmen_m;
wire  ch6_rxmldchaindone_m;
wire  ch6_rxmldchainreq_m;
wire  ch6_rxmlfinealignreq_m;
wire  ch6_rxoobreset_m;
wire [4:0] ch6_rxpcsresetmask_m;
wire [1:0] ch6_rxpd_m;
wire  ch6_rxphalignreq_m;
wire [1:0] ch6_rxphalignresetmask_m;
wire  ch6_rxphdlypd_m;
wire  ch6_rxphdlyreset_m;
wire  ch6_rxphsetinitreq_m;
wire  ch6_rxphshift180_m;
wire [6:0] ch6_rxpmaresetmask_m;
wire  ch6_rxpolarity_m;
wire  ch6_rxprbscntreset_m;
wire [3:0] ch6_rxprbssel_m;
wire  ch6_rxprogdivreset_m;
wire [7:0] ch6_rxrate_m;
wire [1:0] ch6_rxresetmode_m;
wire  ch6_rxslide_m;
wire  ch6_rxsyncallin_m;
wire  ch6_rxtermination_m;
wire  ch6_rxuserrdy_m;
wire  ch6_rxusrclk_m;
wire [19:0] ch6_tstin_m;
wire  ch6_txcominit_m;
wire  ch6_txcomsas_m;
wire  ch6_txcomwake_m;
wire [15:0] ch6_txctrl0_m;
wire [15:0] ch6_txctrl1_m;
wire [7:0] ch6_txctrl2_m;
wire  ch6_txdapicodeovrden_m;
wire  ch6_txdapicodereset_m;
wire [127:0] ch6_txdata_m;
wire [7:0] ch6_txdataextendrsvd_m;
wire [1:0] ch6_txdeemph_m;
wire  ch6_txdetectrx_m;
wire [4:0] ch6_txdiffctrl_m;
wire  ch6_txdlyalignreq_m;
wire  ch6_txelecidle_m;
wire [5:0] ch6_txheader_m;
wire  ch6_txinhibit_m;
wire  ch6_txlatclk_m;
wire [6:0] ch6_txmaincursor_m;
wire [2:0] ch6_txmargin_m;
wire  ch6_txmldchaindone_m;
wire  ch6_txmldchainreq_m;
wire  ch6_txoneszeros_m;
wire  ch6_txpausedelayalign_m;
wire  ch6_txpcsresetmask_m;
wire [1:0] ch6_txpd_m;
wire  ch6_txphalignreq_m;
wire [1:0] ch6_txphalignresetmask_m;
wire  ch6_txphdlypd_m;
wire  ch6_txphdlyreset_m;
wire  ch6_txphdlytstclk_m;
wire  ch6_txphsetinitreq_m;
wire  ch6_txphshift180_m;
wire  ch6_txpicodeovrden_m;
wire  ch6_txpicodereset_m;
wire  ch6_txpippmen_m;
wire [4:0] ch6_txpippmstepsize_m;
wire  ch6_txpisopd_m;
wire [2:0] ch6_txpmaresetmask_m;
wire  ch6_txpolarity_m;
wire [4:0] ch6_txpostcursor_m;
wire  ch6_txprbsforceerr_m;
wire [3:0] ch6_txprbssel_m;
wire [4:0] ch6_txprecursor_m;
wire  ch6_txprogdivreset_m;
wire [7:0] ch6_txrate_m;
wire [1:0] ch6_txresetmode_m;
wire [6:0] ch6_txsequence_m;
wire  ch6_txswing_m;
wire  ch6_txsyncallin_m;
wire  ch6_txuserrdy_m;
wire  ch6_txusrclk_m;
wire  ch6_scanclkb_m;
wire  ch6_scancntrlin_m;
wire  ch6_scanenb_m;
wire [3:0] ch6_scanin_m;
wire  ch6_scanrstb_m;

wire  ch7_bufgtce_m;
wire [3:0] ch7_bufgtcemask_m;
wire [11:0] ch7_bufgtdiv_m;
wire  ch7_bufgtrst_m;
wire [3:0] ch7_bufgtrstmask_m;
wire [31:0] ch7_dmonitorout_m;
wire  ch7_eyescandataerror_m;
wire  ch7_iloresetdone_m;
wire [15:0] ch7_pcsrsvdout_m;
wire [15:0] ch7_pinrsvdas_m;
wire  ch7_phyready_m;
wire  ch7_phystatus_m;
wire  ch7_resetexception_m;
wire [7:0] ch7_rx10gstat_m;
wire [2:0] ch7_rxbufstatus_m;
wire  ch7_rxbyteisaligned_m;
wire  ch7_rxbyterealign_m;
wire  ch7_rxcdrlock_m;
wire  ch7_rxcdrphdone_m;
wire  ch7_rxchanbondseq_m;
wire  ch7_rxchanisaligned_m;
wire  ch7_rxchanrealign_m;
wire [4:0] ch7_rxchbondo_m;
wire [1:0] ch7_rxclkcorcnt_m;
wire  ch7_rxcominitdet_m;
wire  ch7_rxcommadet_m;
wire  ch7_rxcomsasdet_m;
wire  ch7_rxcomwakedet_m;
wire [15:0] ch7_rxctrl0_m;
wire [15:0] ch7_rxctrl1_m;
wire [7:0] ch7_rxctrl2_m;
wire [7:0] ch7_rxctrl3_m;
wire [127:0] ch7_rxdata_m;
wire [7:0] ch7_rxdataextendrsvd_m;
wire [1:0] ch7_rxdatavalid_m;
wire  ch7_rxdccdone_m;
wire  ch7_rxdlyalignerr_m;
wire  ch7_rxdlyalignprog_m;
wire  ch7_rxelecidle_m;
wire  ch7_rxfinealigndone_m;
wire [5:0] ch7_rxheader_m;
wire [1:0] ch7_rxheadervalid_m;
wire  ch7_rxosintdone_m;
wire  ch7_rxosintstarted_m;
wire  ch7_rxosintstrobedone_m;
wire  ch7_rxosintstrobestarted_m;
wire  ch7_rxphaligndone_m;
wire  ch7_rxphalignerr_m;
wire  ch7_rxphdlyresetdone_m;
wire  ch7_rxphsetinitdone_m;
wire  ch7_rxphshift180done_m;
wire  ch7_rxpmaresetdone_m;
wire  ch7_rxprbserr_m;
wire  ch7_rxprbslocked_m;
wire  ch7_rxresetdone_m;
wire  ch7_rxsliderdy_m;
wire [1:0] ch7_rxstartofseq_m;
wire [2:0] ch7_rxstatus_m;
wire  ch7_rxsyncdone_m;
wire  ch7_rxvalid_m;
wire  ch7_tx10gstat_m;
wire [1:0] ch7_txbufstatus_m;
wire  ch7_txcomfinish_m;
wire  ch7_txdccdone_m;
wire  ch7_txdlyalignerr_m;
wire  ch7_txdlyalignprog_m;
wire  ch7_txphaligndone_m;
wire  ch7_txphalignerr_m;
wire  ch7_txphalignoutrsvd_m;
wire  ch7_txphdlyresetdone_m;
wire  ch7_txphshift180done_m;
wire  ch7_txpmaresetdone_m;
wire  ch7_txresetdone_m;
wire  ch7_txsyncdone_m;
wire  ch7_cdrbmcdrreq_m;
wire  ch7_cdrfreqos_m;
wire  ch7_cdrincpctrl_m;
wire  ch7_cdrstepdir_m;
wire  ch7_cdrstepsq_m;
wire  ch7_cdrstepsx_m;
wire  ch7_clkrsvd0_m;
wire  ch7_clkrsvd1_m;
wire  ch7_cssdrstb_m;
wire  ch7_cssdstopclk_m;
wire  ch7_edtupdateb_m;
wire  ch7_dmonfiforeset_m;
wire  ch7_dmonitorclk_m;
wire  ch7_eyescanreset_m;
wire  ch7_eyescantrigger_m;
wire [15:0] ch7_gtrsvd_m;
wire  ch7_gtrxreset_m;
wire  ch7_gttxreset_m;
wire  ch7_hsdppcsreset_m;
wire  ch7_iloreset_m;
wire  ch7_iloresetmask_m;
wire [2:0] ch7_loopback_m;
wire  ch7_pcierstb_m;
wire [15:0] ch7_pcsrsvdin_m;
wire  ch7_phyesmadaptsave_m;
wire  ch7_rxcdrhold_m;
wire  ch7_rxcdrovrden_m;
wire  ch7_rxcdrreset_m;
wire [4:0] ch7_rxchbondi_m;
wire  ch7_rxdapicodeovrden_m;
wire  ch7_rxdapicodereset_m;
wire  ch7_rxdlyalignreq_m;
wire  ch7_rxeqtraining_m;
wire  ch7_rxgearboxslip_m;
wire  ch7_rxlatclk_m;
wire  ch7_rxlpmen_m;
wire  ch7_rxmldchaindone_m;
wire  ch7_rxmldchainreq_m;
wire  ch7_rxmlfinealignreq_m;
wire  ch7_rxoobreset_m;
wire [4:0] ch7_rxpcsresetmask_m;
wire [1:0] ch7_rxpd_m;
wire  ch7_rxphalignreq_m;
wire [1:0] ch7_rxphalignresetmask_m;
wire  ch7_rxphdlypd_m;
wire  ch7_rxphdlyreset_m;
wire  ch7_rxphsetinitreq_m;
wire  ch7_rxphshift180_m;
wire [6:0] ch7_rxpmaresetmask_m;
wire  ch7_rxpolarity_m;
wire  ch7_rxprbscntreset_m;
wire [3:0] ch7_rxprbssel_m;
wire  ch7_rxprogdivreset_m;
wire [7:0] ch7_rxrate_m;
wire [1:0] ch7_rxresetmode_m;
wire  ch7_rxslide_m;
wire  ch7_rxsyncallin_m;
wire  ch7_rxtermination_m;
wire  ch7_rxuserrdy_m;
wire  ch7_rxusrclk_m;
wire [19:0] ch7_tstin_m;
wire  ch7_txcominit_m;
wire  ch7_txcomsas_m;
wire  ch7_txcomwake_m;
wire [15:0] ch7_txctrl0_m;
wire [15:0] ch7_txctrl1_m;
wire [7:0] ch7_txctrl2_m;
wire  ch7_txdapicodeovrden_m;
wire  ch7_txdapicodereset_m;
wire [127:0] ch7_txdata_m;
wire [7:0] ch7_txdataextendrsvd_m;
wire [1:0] ch7_txdeemph_m;
wire  ch7_txdetectrx_m;
wire [4:0] ch7_txdiffctrl_m;
wire  ch7_txdlyalignreq_m;
wire  ch7_txelecidle_m;
wire [5:0] ch7_txheader_m;
wire  ch7_txinhibit_m;
wire  ch7_txlatclk_m;
wire [6:0] ch7_txmaincursor_m;
wire [2:0] ch7_txmargin_m;
wire  ch7_txmldchaindone_m;
wire  ch7_txmldchainreq_m;
wire  ch7_txoneszeros_m;
wire  ch7_txpausedelayalign_m;
wire  ch7_txpcsresetmask_m;
wire [1:0] ch7_txpd_m;
wire  ch7_txphalignreq_m;
wire [1:0] ch7_txphalignresetmask_m;
wire  ch7_txphdlypd_m;
wire  ch7_txphdlyreset_m;
wire  ch7_txphdlytstclk_m;
wire  ch7_txphsetinitreq_m;
wire  ch7_txphshift180_m;
wire  ch7_txpicodeovrden_m;
wire  ch7_txpicodereset_m;
wire  ch7_txpippmen_m;
wire [4:0] ch7_txpippmstepsize_m;
wire  ch7_txpisopd_m;
wire [2:0] ch7_txpmaresetmask_m;
wire  ch7_txpolarity_m;
wire [4:0] ch7_txpostcursor_m;
wire  ch7_txprbsforceerr_m;
wire [3:0] ch7_txprbssel_m;
wire [4:0] ch7_txprecursor_m;
wire  ch7_txprogdivreset_m;
wire [7:0] ch7_txrate_m;
wire [1:0] ch7_txresetmode_m;
wire [6:0] ch7_txsequence_m;
wire  ch7_txswing_m;
wire  ch7_txsyncallin_m;
wire  ch7_txuserrdy_m;
wire  ch7_txusrclk_m;
wire  ch7_scanclkb_m;
wire  ch7_scancntrlin_m;
wire  ch7_scanenb_m;
wire [3:0] ch7_scanin_m;
wire  ch7_scanrstb_m;

wire  q1_correcterr_m;
wire [31:0] q1_ctrlrsvdout_m;
wire [15:0] q1_debugtracetdata_m;
wire  q1_debugtracetvalid_m;
wire  q1_uncorrecterr_m;
wire  q1_xpipe_bufgtce_m;
wire [15:0] q1_gpo_m;
wire  q1_gtpowergood_m;
wire  q1_hsclk0_lcpllfbclklost_m;
wire  q1_hsclk0_lcplllock_m;
wire  q1_hsclk0_lcpllrefclklost_m;
wire  q1_hsclk0_lcpllrefclkmonitor_m;
wire [7:0] q1_hsclk0_lcpllrsvdout_m;
wire  q1_hsclk0_rpllfbclklost_m;
wire  q1_hsclk0_rplllock_m;
wire  q1_hsclk0_rpllrefclklost_m;
wire  q1_hsclk0_rpllrefclkmonitor_m;
wire [7:0] q1_hsclk0_rpllrsvdout_m;
wire  q1_hsclk1_lcpllfbclklost_m;
wire  q1_hsclk1_lcplllock_m;
wire  q1_hsclk1_lcpllrefclklost_m;
wire  q1_hsclk1_lcpllrefclkmonitor_m;

wire [7:0] q1_hsclk1_lcpllrsvdout_m;
wire  q1_hsclk1_rpllfbclklost_m;
wire  q1_hsclk1_rplllock_m;
wire  q1_hsclk1_rpllrefclklost_m;
wire  q1_hsclk1_rpllrefclkmonitor_m;
wire [7:0] q1_hsclk1_rpllrsvdout_m;
wire [15:0] q1_ctrlrsvdin0_m;
wire [13:0] q1_ctrlrsvdin1_m;

wire  q1_debugtraceclk_m;
wire  q1_debugtracetready_m;
wire [15:0] q1_gpi_m;
wire  q1_hsclk0_lcpllclkrsvd0_m;
wire  q1_hsclk0_lcpllclkrsvd1_m;
wire [7:0] q1_hsclk0_lcpllfbdiv_m;
wire  q1_hsclk0_lcpllpd_m;
wire [2:0] q1_hsclk0_lcpllrefclksel_m;
wire  q1_hsclk0_lcpllreset_m;
wire  q1_hsclk0_lcpllresetbypassmode_m;
wire [1:0] q1_hsclk0_lcpllresetmask_m;
wire [7:0] q1_hsclk0_lcpllrsvd0_m;
wire [7:0] q1_hsclk0_lcpllrsvd1_m;
wire [25:0] q1_hsclk0_lcpllsdmdata_m;
wire  q1_hsclk0_lcpllsdmtoggle_m;
wire  q1_hsclk0_rpllclkrsvd0_m;
wire  q1_hsclk0_rpllclkrsvd1_m;
wire [7:0] q1_hsclk0_rpllfbdiv_m;
wire  q1_hsclk0_rpllpd_m;
wire [2:0] q1_hsclk0_rpllrefclksel_m;
wire  q1_hsclk0_rpllreset_m;
wire  q1_hsclk0_rpllresetbypassmode_m;
wire [1:0] q1_hsclk0_rpllresetmask_m;
wire [7:0] q1_hsclk0_rpllrsvd0_m;
wire [7:0] q1_hsclk0_rpllrsvd1_m;
wire [25:0] q1_hsclk0_rpllsdmdata_m;
wire  q1_hsclk0_rpllsdmtoggle_m;
wire  q1_hsclk1_lcpllclkrsvd0_m;
wire  q1_hsclk1_lcpllclkrsvd1_m;
wire [7:0] q1_hsclk1_lcpllfbdiv_m;
wire  q1_hsclk1_lcpllpd_m;
wire [2:0] q1_hsclk1_lcpllrefclksel_m;
wire  q1_hsclk1_lcpllreset_m;
wire  q1_hsclk1_lcpllresetbypassmode_m;
wire [1:0] q1_hsclk1_lcpllresetmask_m;
wire [7:0] q1_hsclk1_lcpllrsvd0_m;
wire [7:0] q1_hsclk1_lcpllrsvd1_m;
wire [25:0] q1_hsclk1_lcpllsdmdata_m;
wire  q1_hsclk1_lcpllsdmtoggle_m;
wire  q1_hsclk1_rpllclkrsvd0_m;
wire  q1_hsclk1_rpllclkrsvd1_m;
wire [7:0] q1_hsclk1_rpllfbdiv_m;
wire  q1_hsclk1_rpllpd_m;
wire [2:0] q1_hsclk1_rpllrefclksel_m;
wire  q1_hsclk1_rpllreset_m;
wire  q1_hsclk1_rpllresetbypassmode_m;
wire [1:0] q1_hsclk1_rpllresetmask_m;
wire [7:0] q1_hsclk1_rpllrsvd0_m;
wire [7:0] q1_hsclk1_rpllrsvd1_m;
wire [25:0] q1_hsclk1_rpllsdmdata_m;
wire  q1_hsclk1_rpllsdmtoggle_m;
wire  s3_axis_tready_m;
wire [31:0] s3_axis_tdata_m;
wire  s3_axis_tlast_m;
wire  s3_axis_tvalid_m;
wire  s4_axis_tready_m;
wire [31:0] s4_axis_tdata_m;
wire  s4_axis_tlast_m;
wire  s4_axis_tvalid_m;
wire  s5_axis_tready_m;
wire [31:0] s5_axis_tdata_m;
wire  s5_axis_tlast_m;
wire  s5_axis_tvalid_m;
wire  q1_rxmarginreqack_m;
wire [3:0] q1_rxmarginrescmd_m;
wire [1:0] q1_rxmarginreslanenum_m;
wire [7:0] q1_rxmarginrespayld_m;
wire  q1_rxmarginresreq_m;
wire  m3_axis_tready_m;
wire  m4_axis_tready_m;
wire  m5_axis_tready_m;
wire  q1_trigackin0_m;
wire  q1_trigout0_m;
wire  q1_ubinterrupt_m;
wire  q1_ubtxuart_m;
wire  ch4_mstrxreset_m;
wire  ch4_msttxreset_m;
wire  ch5_mstrxreset_m;
wire  ch5_msttxreset_m;
wire  ch6_mstrxreset_m;
wire  ch6_msttxreset_m;
wire  ch7_mstrxreset_m;
wire  ch7_msttxreset_m;

wire  ch4_mstrxresetdone_m;
wire  ch4_msttxresetdone_m;
wire  ch5_mstrxresetdone_m;
wire  ch5_msttxresetdone_m;
wire  ch6_mstrxresetdone_m;
wire  ch6_msttxresetdone_m;
wire  ch7_mstrxresetdone_m;
wire  ch7_msttxresetdone_m;
wire  q1_pcielinkreachtarget_m;
wire [5:0] q1_pcieltssm_m;
wire  q1_rcalenb_m;
wire  q1_refclk0_clktestsig_m;
wire  q1_refclk1_clktestsig_m;
wire  q1_refclk0_gtrefclkpd_m;
wire  q1_refclk1_gtrefclkpd_m;
wire [3:0] q1_rxmarginreqcmd_m;
wire [1:0] q1_rxmarginreqlanenum_m;
wire [7:0] q1_rxmarginreqpayld_m;
wire  q1_rxmarginreqreq_m;
wire  q1_rxmarginresack_m;
wire [31:0] m3_axis_tdata_m;
wire  m3_axis_tlast_m;
wire  m3_axis_tvalid_m;
wire [31:0] m4_axis_tdata_m;
wire  m4_axis_tlast_m;
wire  m4_axis_tvalid_m;
wire [31:0] m5_axis_tdata_m;
wire  m5_axis_tlast_m;
wire  m5_axis_tvalid_m;
wire  q1_trigackout0_m;
wire  q1_trigin0_m;
wire  q1_ubenable_m;
wire [11:0] q1_ubintr_m;
wire  q1_ubiolmbrst_m;
wire  q1_ubmbrst_m;
wire  q1_ubrxuart_m;
wire  q1_refclk0_gtrefclkpdint ;
wire  q1_refclk1_gtrefclkpdint ;
