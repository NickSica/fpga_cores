`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
V82h/mp8FbHcv3//3zVZ5VW10Mue/LSt5dvjsUkiSGtG5WaH8H9Fv7j37k+xy+3/pQvfXcpqBF/k
iaz4/vETUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n4WSOWV3uUjyMD/l4IGcKD1bHONRRplCKgax9lu4YRYlORLHEpckVBvOD9geZHtnlLIjTLNUcuHS
rc4oO2K5x66eEf5+m+hNzaPYWCrVKWQI7/tyX0imMAsD4JQXzU2CP3ATsQoldRyYOQZmggmbIMiB
stLQ3uoRuVc4t0kXI7U=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zgo3FUzRcS1G0FRTCr4C/JBs44dp3dv5CUvkYU2vM2fDyGtu9ekJcjDXnFGi3Qx2X0BV1gEyWxsJ
xqQkFlu/f/1mutspkUjOMtKZNCgPGDHkGfwBEPN/xT22fOBwQJUR+Oj5KSeDWe2U4t5UJ4XXcGMb
ZV9syPFreDWYOTWkkl85cAKcf/WXC6oz+tOUowqV4nSLA1PaSrK4ohf8oaOGNVX+4Ji/w6ViTIJJ
OqmPJQ151npm7Kbt4RW80tp1OmABkNI+o6h4rwtTS1IHzM6bJ1Krrp0V+2aEmmqoZkuKINjX5Pw3
P4Vi6iUmJI0uMpdsCPr3MEC8HH4v95WCnjh0Qg==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A45QQ9IEoKpoNXpmniz3AuFZmGAAZIhtA2hP4/pi+Iwurx8nPI4ZkKpYXPnn4DfH42bSsec35aiS
Ve+A8f1Q00bmFgtclspinRe4YgFesk40ftn1mzy6g6sLCNXhUm/IIjCSNk+ie6jVQS7STfOdio+z
cvSm8QQePoJjzlJz/jkNhsD110PhDAevJWb+C5fforY6kT0k7ZmJmE7btahod6wU3o7t2HM6+XGU
DDNZ5E+RLS+IiJYVCOwsdqQFDuRaWwS0k8Mk4UuDiVWtU0+QLFZ/8UGJhy2ZDSYlL/8TrrsWcD/1
Vku2N+fkWCj38RSMWEEe5TmUHSSzP7uBI6QwVQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b+wEsHDGMmVXUM545W/2toIjDItLsHFsIOyFDid8Fv6KhzBePVZlc9t2c1LfdAa6UEpdqcx5kgIr
+oVEglJG3R/fb6dRp2mvlu6+x0AYh7FK0My5t84q7uKZ6EPBxHnDds9FLGQdMDUFv8E10WtGrG31
lkto5q+L5WLAzYgiD3//MgdbP+aqLc/75XWIRhw/PfRn4OqyBU7xSBeoK9TDxBwOscUv0cQ+dauJ
dUQ0W2ZCXwF6cP5c47k76Ikfu69J0/IO+FTLKMkjAB7Wzsyqbpl6RMVdJ/iYscNROh1xxo2k+52w
4l9VnVKN7wTWZdW75B3V/MsNTrKb2I6dBdveDg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Uyn/owx08GdB/M0CwlYM5XwpK1DLRGgNdNGvCa53fvz5ftb1LM2R7yhWTTXlm8iqXlg1S70wvPmw
WVO2ZNZ0csmDdQcX4HNMiokrI2gpR08Dk8n3nzdOhqyFyh79/eVJzQItyKMQmJZNCvFfww0mtX5K
FbNe2x6ria5jEBEBp3U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J8WwILioFJtk4e6vNsFHYZhWTjvAMbsqHcnvhYKYzsY6fpaoYuWnjTNNNxS6JYZj7bKOFgPjdnBA
rKaGPLghV6UU9fx6UcBVLjNOj95AU3CZPEjWGC/GqjGRPxOkhGtDka91PZuOBRTBqJT8F+5qIgQR
vO7WJHaKezpaUm2zbeC7+ShM5p4Wm9L4dzJ1OuUGZNm39p9FbORAZNzAWa35wpfJ6PPOgATFMi7Z
sN0Hg00oxMFCKSg1bxvN3p4iC3rVT+wV6yuzOecq97B7Fu+tfvP+shqnUhodTpF0WYfGWHeK9ocM
Mg7nt62XJybi4Tm5rgYGMIIM0i67934etK5Aig==

`pragma protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AF8EDKLpUnsf5U27caIfzjHsL1dKCT4FvrlOxjBwD3ZJ9vsXwbWO+EJTOJOFymKnoSSFnuslr7C8
ZCAbkJJLJrLXJwfvC9hiPRksxuYzuxWrtwsjJd+5KWtue3gL5kHClD8Tbo/V+Dnr3gvKzMRNdFRz
i+4p8dC6/32xR0/NITJMYT1uOYu0oBFDHGLR02Wn4PqghcTR3gQMVeL0RsDhJibeNnf4Q0NsKqCF
7OscDpis6r9ZAFao+mdpLGI93rreTlZvJBUPh2RcpqOjL/8IUv0iM922KOCZ6j1LtvD0igXehvHa
5hOx0DDcMjOoejqJiwIqLij0FB13lDBsu+fjWw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 34048)
`pragma protect data_block
BMP9G5RAk03qFRu5UmzfhEwWXVNssrcytF3IPfT2D1Y7zMepdmoJXiO60J9qg8C88NA9LyV7Y7GW
/BkcJir+xcyyrAUmxPTsXNJqIpYv/2xiZOu0LvfgxeSZMklTV3gSYEVIqR6TBQptZc6tmB8AoQrR
zyWNOVO2HCDIZVd7//y7GA3kvPi3Qj+A06GgKfPILeSZlmayQW+4oEHX8i+eb1pvAPfqyGT7LGPg
DAWMso9ERRTCHVBGnERh9ic4VEhmVFh/k6zjE24YBes2m+N2ShOQVs+PV3fgFN9ag1zs9IGu+msC
agBNaDcuNFgz3Az691GXwakgdGlw4cMM5iVJPcdj6Nif91wpgXzliXm0/BzwvtLNLmzHMbdvg3oM
Eg0IzKZntGc8w/P2KRFMeY2XsnREkokxrCF9pyofaRFz8p3G3SeBUcEqegsCpCS382fv8BjaBcah
PfVC14p9hf82JmZAkFDS01VzRbc2VuOlQwVwtequBwY9LWLbyVoPfGSr0xB1Ly0gGY2NyafWlqh7
LaWGJLJYiFBgSlVVOtr2+T2vaVY/OwZS5Fk15PA44uUQrmJ7sZfPiEZRet8wq0g313AkV+tGrBEW
6a3ChPbenuVystFMc4LOuspoj7+jyRBBBmZEqua3VP4f9vWBYO+y11lt0W33ZXx+TAqz7vTaPM3p
Rt3Ry2ELCc7UtQ1smt7bDNePugiiHKLZmrb4UFy+yIx4/j+7iIHTiXyQfqM3zbNqdGFjWtEbgBKf
rJmBC3xw50FjVkiT7lIq+rsIgYGH+dtM/kF39ZlFXehDIBLdjecdKnqLJxjtHUXDeG+jpUsKTqHs
WcWtookLuVMMzsyhtx8N1LpmGyI+RHOv+o6glNpNu5LwBlegN45yz3XvOU8mguwfDu6jBgrWsoAc
Kb4vuhtk6DXeUrjnLfp88JkXuRDXeeQ3O3Hgr0XePW8OSJUOFuANc+2haXwrPhuB7/qRBzHSRgLh
Ct5ZRGzqpP2/Ra4VP5c6LQrQ4OJDcGLMxFYFjaTZRNujWfnJ1lUOngO/LW+cIfHrJvLe5m1/fCYl
5H4rfZPZOYpxa9g0tJVSCml4QKoBJQRrKrSV1jpW5/27aw1rUNv8syefxd2d3f8tRadAtBLFaBAx
cEr1noC+fmO80MDsUL4f8JWTNmQmLLLuFr50dIE/KwaO/sK5AkYtkz7mt5dGuOD+L7kURpAGhaBj
vffMmMMps/1a0Cx3f1t5H5qJ7ZWAnFz1E2cQPEvxAfhDnSHkIVCM6t6gRGhbaF8O6k9w7dXHWkx0
+obGkIsDJkpfMoo9k009MDWPF9lrKz6YhJS0qoRnTO6uFFsudK0a58kJpnxWbei1CUO9A4wtHhdn
yxndm1/ZAKJWqFEWKfcRyVNKAKI+NcMF05eylSUbc4YHwqir8isHJxnQzf1W//ou88KIChgH3JPQ
AZP0Xr6yQxvBKQorjSlfQJqyRuYg4sRdcDZ4arlnkFUBBzpWj4tVfTH+DU/eGEo1d4fS1OA3oLPJ
x5IVx7uU9hnMgnrS5CeTHYZ0+b9X2TXKnuKGFjrPTWQhM0vvcHjvhtkUZLjpwNGv0e/gSZY8/nAK
d2lRP6vdeyBzCd+0Usy+ArSo8KfuA0r+MVzSMM7V5rlKlj5RRnomqrMGr2CFwKy+EW53wuv4yN/u
57UZLDVpsKeP4ihVA5N7kXGv37hDf+vwugNVkn5icAXeRMOdy7Q0+TdEyMUwGpYxa5ymCP3XaEw8
KMZijlbkbUNdXw8GjAA0FFGrSw08OOgyYU8cBsxfwriO6oqEcZsz7WyxyxD/ex4Ov0cFxmpTJGXB
fMwzao53TMUYOd4jrKWAjDAtsplha+n118jWwrktXvgs0adjCdsjfMqbRefSq+RwkPjZPfts2YlS
1plKUP41dN2kUGDyu97vvE7DBjENzt813CNGIbRkBX4Voa+0ndcBRhsr2taneVW/9dho/PFGpNNp
x9hla1OzNp5OH8Swun2LErZDi/FW2PAgqG2NxSNtY15IQ0GgfpfGhtkD5mcFKyRdy7mS6Y/G+LXS
9/5SDg3PrqnMmaoPY5kT8s5wbZ3fiC5YEliwxZ6/6BxuVOVdvI1LZ2ixvC4nAEVMF1u8Xd/CmEw7
YYXyeMHjiYej8DwyR/JvFfVZXgxK/kJHJoiZ1w06CX/JXEpafUcQanMIyI/5Y8nrG8uAEAkVNhLf
SExmhV1EGs2Xdg5IbuVytzo5lVfQDNUMnV3rxyREOT17a7Lj2xycx9iXDIoivC6WkhMMcaheNch8
P5nruaaZyrwPUpgMK0NWB7WqA9GbTlPJXtWl2W1Kq1uD8MmpJKbY1QAkutab2gNtZy7t1Pkv3en8
hlIWDK/OQnhSfExtwRwJCCZ+yb/v0MMbukzFqg5vumn8U8YHcwfnYxcZ6dKCuKrob7lTAUbaBH2E
qajcNHBvZ3sVUza5N6v9sspFS8OIGtI2d5ml/IddOd/3wORpFSMkwcVkKxFOaSigoG4U6PyiRgmT
qweRuOIkqsv3pDtSNnXy3BymJ2ItlvUnDa9uRQrphdjjYngCLDjjplreg7G/VR27rB3GqGrKsftJ
gr7LgwJAKUJYMrtIaJpqesLl+QJfRMSZNNmmP0veEFOl6dkfAXjh0WRWqJHx8Bp5kmHx/EysDQ2j
rK8+03/jueFN79msmd2OsMOvv7y0B6UNvwlq3BtuoPWCrPfDXdvusj+/pEUeeK2/xwVa+Qx0z7ZV
Qp0lSHSiryOb8k7B/9r1DP/bhXk2omS1hZ7qnQg4G03KqeKuaEM9pgAg7QWEzOHV/dYN1giK9y6d
NGSpChFFLa3AwwWVdQL9eDHRwKzwow1LM8Vb91sbNnkCSh57q/HTuNc/z7h2qcSFr28oJYyLY4WP
Pxg5NHoPnsFmyDob5WpyQ8M3kWf9p9I3RXPT0O0tw4DbwFo0ZhfRZCfjn7Uq/WY1+ct05lVgU4mc
u9oq1yRbwQk8q2miW7SqsdsVB3vuVRrPpUJ00ulW8v5RDuxCT3uu+0vqhUqNXTahokdi6EqFnIeH
zu4PRrFd6Vzhg+idmV5+VJh4CqwpPeVLTvh3L3lXVZRXPGhV9S6cvWmemMG84MfToSLURahSAb4T
nVQTt1xjp34SJXB9McNCHmYnK3ImjgfDFLGpMrPyJp2M2PyG209XgR7LU2QmFQqFCv4Q5J+yM5MF
+CHA2h+7D1bO8Am//0LLNFILjU89TMYtdTWJynBcNKpvvJHYIEBHyFe1Omq04+HxDk8rg9d3H9zc
IssPpvSiDQTUD/Ur+8ocvw8Sx9JC2n/zkEjWoygAb+ocGUMzIve522FaBHOaIIlCS6dwfa/V6wNF
oe4r+LjoxRZ0WqQMIearPb3xZl4SiLSN0jZMDlDGm1NCpGVj9EXjEpXg2Tx/kmzqZFRsXnwykmWH
gg1ASqK69aizEoicfZ7saM/FBc7pq+kk6ooUxLQmG0B1aVitLRUBnhHAt+xflRkucwGLr4uAwvsX
ErebjfFah9VCSS4/9Nj1GLpEjbtyIDKg/LCzFZ+cAk4tP1ygL6j+PbeJ1JRmYqFynqNSA6WeDwcL
nopooJLbmz2PL+7l5qSW6G8K4ndgsZWxxk+PiCQfOsI1SahUnQQOQ349LhZuxBBfjHUrnO6MougZ
ZcMMFp0fNemCU7drlGgiaBnYN/eZS2FltM3GygTMFeFK2fE4Hq6geTTJs5KxfHJ+pX9fcXm2Zpwi
vHJHmEy6RF4sbIvq10pMm5X9/yAd9n54Dwo4VQ+sdHg2rAdWPrbvp65dS3Ahrs74NLxh1RgcD16k
8NTi4HhuASSv6fhMedY1+eA+3GfpXfCM2K+ClhllUBdzBFVl2e5itU/0sdGZU29ShtJshYekqrE/
40hkB6vxhtfabyaM3cLVknu6QbHkh9108SkCH3kFCzda/1O/bmW5gBwXdfQmCvPvbtddiVEKqB4v
I2Q6uaw7fRYRKK7KOx2BjZMeTtPBHgVvbzo9nkrXpUQJ7yfYlut1RbI7LvuUEVj4u7gT3DxQLqov
z4mQ0R5ryPFD9BA4t3BabahTvBvXJq0LSVmobCbPqKUeQBCZxcjifwKkoKTt9uWaB/vYPIEo8RLC
PBaCdWoXPSHWsRXnzNerKuKX35Rytbp9lLDg76nnds650wUXF6GEVB8dm0dzbtNOfmacEGHf8Hx2
sicpxeSurlXbLdcwZTwC/+kEJGByuCyo7rqGAyrvj1o8ES4aKfUh48QyOu7vjSPhxvuS6ymnC4Is
dwlgIl5PHeB29u4hBFL79rDyxutj0fRx/W9Qfs3onAilzAEvTKL+9vTBTTjZPye+3Cx9bsRIciy6
FJXPeyoE/qKESQl3EnMEwlOU1vWXCbf2+p4s6Haujqtv9fZ9NnfKjzNRP0sjRX6qMxplCaMzvleV
nXknte0chkaIDW885FjYx+OcRXHbB9uO4MUD1ZePyzAVAtP3OB9tY+IL0qIQvNyLabO/k3/chN7f
oN2aiG/XcAQ44MUw/dQSTO67l3+zhKRgImiw8RtwQ5EqAX4Dlvqwkdbfbxkq1HXbduxJuIWCX8+/
4ABRCb4XWfvujVhzdPDgGwI4k0BjN1g4gIX22NT0hKrGXMGA2WAt7qAYipDXCDfG0/vlJiFtc9F3
7kH+VXcw/fZjlRH0HOErX7wXPE4FfebJoaAo/WEn1r+/0Ksn9xN5CNDqLk476IN0IOnf4AUo5DeE
d/GP7fLv306/zWexY4clR0oMwf6gve2WPtkZ0GqL27/6ukaqsZqbY4Hx9Rp/aIsUD7+7WRWsh22f
8p6IZYzAPmGnA6okq5u5XVJcLmJpOaJk6+HDTnjDVaJEVa5YOsEkYrbIEdA2GtkZRzdwgM/K0jcz
eXyteH1hisjtLfSbZpZE6huRUtwEUO2Ywe6KWyTpnS5Lh8pU65mgiLHWZAt0UtEkHOSqgMVgeCl2
7kzKiBEigEQnSOjk9CbiVvTeskaBjxwSI0UBgCf3XbpdCFFDqiVIrSrFmySADonvi7n1owmD7Gxz
ICjKvezSvyyr4wU8ggo5kfi3cK/iW4V8HOP/aNz0lA0swSFlA2TS3qM4XHiDJD9eOtdvJX1ucHt8
1dXcVs/buSb4uauc61qybgXtruYI2FxOtAxdFq2FSLvN8Vod6A+6w+2oMvtLWcar3pYdFwGL54Yk
XDDfLFMrgoDzauNZX7+8wMLkt/HtnGlAMq7SuAPnhYv/bqdgN33drEZSvb7+xotghcDCCjVPEFYc
1H0G4fA8ZmuIzX9LgMRQ7ZZnqYLhyQACawpWrf7bdP4FBPUSD9+VleacQKbvMKobZFc6ELphzx6g
rCjee6miibcIXPNZVVMPsDG/9N3sBCLr9dlrkSFKndTF96BujJwyXQmeOe48kiO0kruRUFBEnGAK
7BTzagBxDd4xYWIYR6G/ofHyXWC9yBoe2/Lb+cUODIAcpGqpP+xQvO9IYoB8EZtgHlgD5rDrRsrx
Gka1zcE831dyAoLD3WctiyooxDaqPN+LG0GqsXkflegk4k1wsy4gAjd+udyiQ5TVOgbyh5mOuKSX
pHkbbM+ooNO2hg2kYmPF0X0qEjjOYp2snPVjC9Uons9LhGGS0hI2AC/ZZBfYyVTo9Dl5isq+ICQI
GtvIQWnSJyHTaQooA8g7WDM1/lT4g7AqS9T2TU4wqZzVDazU2JdTUiiXue26vjQMYDZJFUKKg42f
QTkfMGn49DCtUKd/trLTkAsm+Np6i4uluklTL8m7j95lsj1H1fm9JUX1NxHP3ig3VE+kpkXgJe+M
PFTLKJA1GzCaN8VLe8xnSAQa4xJcTxQ7GWBwf0BqcZgE6XJY8wtYfbUQQ3mbHa+tpVAsN5gqVAek
rd4o9eGfvNpN1k1NT/aDFQGxs5jCNXge2LQC24MwilBt0A8gd5k/5oKf/qA4qLr6JZvoZ51Dh21i
fXDJyaO81DbgSRsNmtEU3AXJTxZQi9TwFKIhiaZBss/48x7nfBYY0lRr8tg+XaJSSUyfADq8fdT1
Mzd12qmsU18/0lPc6mSwMz4TNYbESo+7dZtWA+B3t0bgoQ/VYGTiWby765TMttaBC68JS3AWyvfi
usu5Tfzqlm0Q4Df5eX72dNhp7OUr/J0V6qf/70Gwdggy8lpvTPHB8kLOW4gk14eLQsmszYgTaf9t
jWSjEccmm0/n/uHFP79fhnNSkzYOFAlOnk4bhlam+k6uJcKi6xpdN0N3mHfiZz0GQoksRxqXedT3
IEdr7eLnNAyon/rBZQNjc/rZAVJhvdFu4olAda/s10xMTk40W4os34A3nRGEHwfFLLc3LOdeczQf
abrSjsNBheiwdsvcXRfi1fk2qhyk3ux5JC8oVp7MaGni+aeC/+Dds4ghLTzq+c+j2Jx2m27omDX0
lU5LjWNgiun63nPys5v+EwfOstnbmNrFr52c+3lJ0G2vaFH6zPTheuYiRQR4BjbqXb8p/9g7JHNw
Z9lRMHdxmWx/G1KQ6vvxkHISabZOFiFeQrNX/utqPh7v8TU8GewP1rS/aBkf9IrCA31yAn1C/l17
zZkOWNhsLis1ESpGz9CV/PaJSH5kwQFvVCyYHetP2kYb/NGiMPWCxpuD79dScDR5tevLyyZfgRd1
sBLTJJtxa7Cip6sr++JDKb2fDb8Mwx4+GB9IbYQsAfqivbN88JL72haCNVRMMFCsv4xESsWoiyr4
mCDTzHQZYZPmUcUzlu7A75vbyk9VHBRTExdpvB3b9GHSy5WBSGaf0rGwDsErAXR1JUGD8kH5qRvb
ugnoq73/Y/rbcasB3S2tQOCmNdOL1FUBn8RCifneFweZ8B2wM6h13ezI/ifAW3CW/NGhBDcYm5t/
rLX2/SebZS176swF+dQihNBSa/dMm1DCF5tjW3dWghotk729ilbjPuppLpjsgd36rpungaa1O750
CmoEPiozAUeliKIqBkwkFewuNfp22a0rxjvv2k7aBDVHobJC9aUzrpA4/MGzAzKMaOePwMVvzWRq
CAVN7zzTkg3VHH8Dl+V85toqbGttSEUGA/xgl2Pbyh7RUHAy3e0Y48jXG82q8UC9+HBjzWuXNiJV
CiGHDelsqzp8v9NR0enfH3yOx06b9G8bSJushp1otuzO31c+tpkMrOL3sI9q0z9KxU0F0py2RPLm
1dd1O6O0iRs6K2fUQhpQvSrk8HHRBVb6LoJFD8N5lm67QtfW9WYHijRuv34ajOo0pmyjLalhzR7Z
Q7rrs+hECNUpUzq1oC/5UoqquOMPZzk0176CrVvBzg9hh6erb/AuhFYs0TWo04Lqv8r/FL2y3jdl
jDhqWIcVhMAjmPoU6dLM0+TDiGQEv0R/+7R5MUxYZXZOkLguAfGcjL2kNbnN5SeYVTE6snQImK1M
GjOw0ZAYDDQCDrhV1V+4TXoMhHB1Mm0xXTaYlwdKNtoTD2kp0TEYUJD0UmHIO1nOI9GYAF8vigHg
pnM70FS4m+QZNUXyQxi0ITvNbEC/6RHr8BJx8SX5YmUngapFMJGlYRtYuTTy1mBCNaqydU/90xI6
obj2ZHoGSHfzIsecAJsX1ZK/egkAY67aT8HmS4gL83hA5Za9U2DPfYGyvhNxnPmNPN5zWJsXogtW
qYY7UMr34bvGwVPWJT4f9VQYSHQ7zi+OKqO2HnAz+l9q6hegrHfuz3rAB1bxNbX3BoZZ4LD2A4Mo
mGrTJclAkPRIPSW7GFgEEoqgzASr6l+KmmM5c91w2o4Uei+4eFb4A0NR+cAgHRLYRFeOBVLOtpeX
EWElkhyFN5DrCIRUr3ZR6L3LCtdXPYoXn2KpiQP1JHDdt08nFWTFZNx/tW7uhVlqTthzIv4SOjvw
pInUwtwaNBKwguZDAMzUXYvPadspFc5y8fPsQ/G7hz2rDitWb87FAtfd1GABpcffXhozeD9KvBRl
6n5yCI+KnHVHjAGxzVnChghSjdDN3prFy9BzRXcoZjU5xu5qs96jFua5a2lyT12yHtVs4qOejh9I
DoU4WbdEVFpOMc/Jp3kL8HWhXs+U6av3EFfF7Kkmjl4twF3uVyiD7/VgPKJhZuewYybH5AmhNtrW
gwpv/2G+1+kV+poNEin28EzGzrdiuX/EV1oi0ULX9mhD5735bXp9SoD64g4Wd6P/HsfIUQEodHRY
jMSJPUUHg4XXyGfgNqLT9Q/PMY0JhuWXem73Ni+wQ5NyC7URq6H+rPDJN2FErsoJ/HbCWPI36jcL
92AvkdM1HZ7/QIAW6QgdmSnTmlBVsXJ1j10PoaB1jrSTxXlciCgY6eHDboDyee/g5BoZFbK8RetF
hSqJGt3udd9zDrCrvdDapb7Ly3+zZszHdN0Lug1O6ZWRUpcFhTuyHlOYXbNVsFfDfNjKDGwWjBLq
H4nJA401uDCdfMWnHebqOCVdNPbeyjXlz437i4BvpsFEmwkiIMty8MSbAb5oB9G7GAzsZY0/JMEY
oknEs/5BSdwlSmiSYPkPp66LtPJvlCjfc9F1qb/Xl/8gnNEoozCkX5I6gVb/zIVRqIY+nsE2YXD9
RL5jUyp7srJDhPi+LRotRoX4az3Lcn5l4HjFBLp3QAAAdAGTAwGgIVcl5fIrUKfYpUWcRaiLC5zd
N2Lc9JJZ2bh6GY2rvguU8XOAjKSj8wwzh5U8JbhsftPzfqYVvYWEpeMg6b/hi/Zn1S/b1AwLaTbD
SCFj0kddGZWLq99IMXBd5gO+Jevsj1tNqC4a3VFiu1CvuMY2u4FzVnxolKBq1Pxw7nfe4raqgf+h
+iT+WuOMU3vivEbIVVLZ4/r2xotLRzj9pulcBRMWqQm42PBc8EzgvjE8Syl6vD5o/IrrfToBDc2f
jJqe9OSEgWFnQf1pHIquooB4eS9MsApB/RuW/i3I8foEAhw7K1K1p9pS/4BqJuzKCdHz+0/SGyAS
3lmia+Syos3/NvTlcj5iq3gkkuyoUfm6tOqagX0g58g3LbQF1/1hK/8uupX9+qrGAasH20Dko7v3
4M8J2J/Ytl2rwh9ydp5RRQwH1L01HjpIi70csrRywLKtdv5pISvCYO1HQENiKQ7bWA2b9TRcnEgk
zsLeE/LlKCuq8vXQWUEG9MGsk7HCeYIn+z6SOm6aqHg8btT58k5N/L7Z1hu/JxKEzbEDsOmfxAMb
QbM4oSoBnMd1J5Zes4oG/ESdpnb74sszlnr7RIQ50NTovJOSjzAL4djIoc83Mq7SEEN85yxQ+pH3
UWQjWLlJXksrJf6Y8Z9CyoOpjGuOIxYRDGP80CKpsYc9K4MP4h0//4XqBLqy0HX3kFmvMJXO7fo4
dcvJWOv2W8YkXMGE7PhDizqvIQh+7HG+MdohRQNCg6uUTC/lV3bBEdyzSfAH0AZasGUYNW0nDBzq
xtLjKAc8T7TSNtoRRcDMOyntB1X4jJcMME8oA35MphXucBgYMup0FN+5OwoXA0kqEI8OuTLaWzgl
XRO5OIbhKwNwR1iiInhySOeMJGDT1A3gHcD9avW1fz+z6t5idRKnfKvw/C+dgHhwfIbZ8CdRHtcU
mAlR9mEZ12zUH93lm08rrzMaXnLVQkkq1t68JdQ+1wEoqHhQTKqOBVikRewhax22Gw6aIGOXMdsc
mGT9dZhhwKZorxajplR3w188Yy3m+ZU84Xf5VIEXzrn9XFn2G/jsDU3/K/e2Omvx2zRi3WGNjh1n
84fQvtoiscAnlTINxtglxBXgsLwLfDXA8UfdHZRVqMV7N8e55AWKsFGgIbyeUhQyBPZBI/r5l4Iv
Gey1oqvl1/mePpiaGJg4ve9trJdBeZWlGy5xQUx9IweQD48mseqWhhCLQTuPrbTm+xOuH/JlkIM1
Q0D2+fxq2yEgTNCZ+hR9KXVyv0XMQbSfy2v7pb+wdRPuH1TzTUN81M8m/zheM7mBZYvPTATDtU4G
ef7AUPJMvDpLR9KvBmtd/AvfO2lugsQ5yRIlUbnyydo8o8Osor6B8oub+mhiP5xEl0S+Kc40/MvK
a/eeBkwfjPPqpB86bIpy+Y17HY121LmecQkOXndhxHpdYlKdIy5bU4qKskPXhmqFQpXdW86Xw56n
PBxffa/h3AV2GACylAloXzZBt3/PjVXBqd8OGEF5qLwy9HrHTaacGW1paty5FrOkQn0rMOKLTkrO
fplg2VaoiRB6Jzvmz6cqnffMdkNAIXcc4zGiPD38c8mL3bBNTAP/fdQi8zJU8NtpLEykGz0LPRg+
0p4IMXo/s9A5q0/1NJrMUZcX5lYliqItQBRIKFT6AY5xYfYUi66Us3stWgrpEdU33tSfVissY8BQ
Rr+PZhExhcXxEioQEDdr+9d4r0ukSZft5thNPSNity/Jevo0wk2XkbKbM6eQbD/iLkmucBYZ7r17
4a9XBXQ9vA0pJ3qz2QpNm1s7bcrGbk5umXdxWkBHN7wJQNHe6ZDi83NVMFQZNuWe9jT99Osj+NxL
7FYA0dRH70T+qc+mUWnLtyxho2k5cMUTmo360aBDsKNnBT+N6KFC0hvwquIfApOQrOhVid9D7Ig+
fAjqzvW6mpXFmgUy+0IoOPcBLIGz/dKVI6dXN5JqoNZ/rYFoYTldlup+UQ9y/i4ia8f2I/w+ijZh
sHc7k8OiJUOEoQ7cqU+52xAKsRw2CDk+U3ccJueZHdMhtNunhkYrx4fWX3jVC/wukuxrpRRXfQwX
/EbECC84AXweXQUlPk3X9QQOplAwSvOs7fd/4flsTbNL/tVBhzPlDh/l/N25GoFISzW/yB1bunKS
gDIKYFeHEeMd6J3TO0tRjsXWgFctyPMmjjmfew2mk0OCXwjR7sGf9hnmHvzbOBN4quiRsXhW0eum
PEEEjFlPuB7SYQwWTo8WX60cvtW00A1uoQBxwdV5FwML+3vZpEtlVZTYiwhrOCt9eXjrWZX/HH86
YUtv7f5NAEVtyXRCkAobrGO3bptKgNyHHOMC14F7dYDi346Zx2EtDF57Xy1Zlsus7ghZGv0tUoD3
I7QeT0buJK+aVQ3h3CPw1riRF/PLAFx40dpBGM4FACuCzj4pjI7FdkGpjn6GSl69/FT8p1jnjDsh
IAiHiE2id32s3tKCSVlY95/SlHi/6MgLdPkjNymgrFO1+YbEVN4OwPWFSsR49LCBlDA1E4Rp+zIP
wUrhhvaHMYEIXcT4q6a+3gbESMiXcHepNpA7Pb7uKrCBEVF6xUuouOLMaWXO+ZCYDDZCoJ8UmKwO
ASE5KcEAIZnHni4zPKRwwO7C7LWgheZPSUnYv6ouV8OuUDVV3CRuVtEEaQkTuLdBiK9rHbf+XIsv
WbscKuHvMgYGVigqcnoRYiPXahMZsfYZE3qD9CGF6jO0AeHW0nG035E8XgWe9xFEoS4F/Pf/Ww54
gnakgQociTTXkBghXE16trz4LpT3s1ilhMN9lIgksjknI4jd8s3BYS5t5nX40HRfBnbtQjpHLIL0
2oxndbrixUgz6DW1Rvvgup/RZlRSsyL5Mf7Y7GA3zYcZbVTdO/ZlJl5+yJLlx7B+Bdnuk+okXgx3
nTtkg57eHn2enpX7GPvuDZoluUOX02Qkj+i9Z4UCbr3V5xLnfue18xRDgNboK0LQt84ZJfoVnUXt
gowCKgCmRMZ5HAW15S4+n/+soz5NzmOsVuFq+KtIAiEWlm9uxbOydB9OUqsHvaCRqm7tCimI1ZwX
heFlUK9zd1sqE6G6bVP3xN8GssRMPaL8TlqLiSbHMeRKyq+7EXbfbhhvAyuDG1s+6AVyMWJlPPwU
V5W+Dni3BqpNHjiKlURQyn7YyZfpnXVe9rP7HvB4WknXRhcQmX2QK4NRA05rtm+imuSxk5pHDhDP
UzuuJlLMyh5zwxzOU6M71eSajNLCbaHEnUSQqXHngeGbNZadNOU+Qr8SKYdjyCy1SguT2YruVtUb
V50ZM+qHQFqcZQ3Eu6RQywOiPUT1wP9UvXdJT0qmBtzELHxk8ucsxzkotL5/baP+Bm9Z6qieK7Gq
552cpfa0X9aIJwLwOkIij3dsSEbuSXCkuyw7jWKmNE4nMOn4RL6qTKylFGu2DVZDGIpcytJPY/Ts
NaXLvaRX3VksaAElKOB95cG7ptzU4Cnv9gqBeIlublthTGt8zVHf+Yrc9VORa3g8JicgtzKZ557P
SUSmt4xKqNsodOhLBL9DQlNsooPQLLXlHfo4o09Mko6ytOcPqciz54UonSnPFSYBKRxfVGMPIXsp
icHjW4ZrY2V/1rYF+kTtbz0OW4U7b4/pMK4R6uQs10fHKv4qjwCfyXlCVa/HH5lOdpxppSk4bCgd
XghdkeUr5dD7H0dqDNm/BN6SxXgpSMMqEwUQu14/wn3UzDIDfT6gEu7oVIV/czswGqbn3fy8L459
+VvLOtZ0om2mGkZzYlP0HHdB6+inFqswv7nImJc2sUF1ZeHb+C53ZedV7umc5cA/xiPFcE6e2G9a
PG0qgAyHIuOSbM3j7yGwOEDyta12qhGDmEv1ENpkoM8JFKz2ybL5JGHGGNnRqotDqNyyhXmuw85u
VkafvlnDw59Fsu6qc78ATHYl3ep3dIzAbQFBUHQhd/Jp64umsZjiMDqrMR5xZ9n2ORTTTB8Kkhyb
aVEVuPil7zlKBJAwZh5kQlduuvf5uOaBvZ7acKkyYFAAYAmi5ITKgiyDV4EPo51R31svKIJGQoG8
eIJ74/ANrKKaqWpvVFQMID/n8zGuzkKhb0SxBugcdKPoDC0FatRYQ0LG6RnESkedc15rcsMgRHTI
7s6aoA1acCi1AoYeWWilzIN6J1/GlQGPmSHT19W8u6N+YLfN2dToIs9fU/ql+6stEoTUXM+BP/yC
0ghkja3o/fGIRXPdrcFMre13sAvBAumEqPEvb6ArXiZg6K/o842OyrynMec8N0lc0DycCQCaKoqz
OGcBO1c+r6HxjL+7iFIprT1V1vlE3b7sIAHXb6u7qJ9ndySQsPJMeK7p3JqI7cms10TeKPj9pCAJ
4RHHQvrQuuiCRO3XikKUL9TUDht4tr6VAehctzD50lu3xSnvzwk019BAe0Thn04cn2OnNTDoX9pk
FUd7xo9WE0GU8McUEa3eaCeQD0Hj0Q2dlqx+fSoQdlqbVQFlozdtOhcpgeEqFhQ9Q/vMvvNzgya2
cYVKJGAcktcyMxQEtSA9VhgPk2tYy1KQrY/MnVNq6VEZA2KWeb5Eq6KfvavAwLJ5WW9bRVO08B+i
rudNU+gVJfMLXxZo6xMVY0jjJaLn1xT1qBdOl59uEXstUXf4pPViRUe/jiFG7Xedjv3X4nDPutaR
3aPFump/43lHQDI3qfD6FV17iahIST125LFy/cwXDA/ClVfsnEopIu+1xt09pBU/oI+kqo6qwSI3
xcN/xYPyhmiEN0r46ydb0oTeaH6zbDgSZDKTbz6LOh6HijX4XddaAAfE7gfaHL+Y20JZ+FdZhuku
hq4bIWpoRX14scQ1S4D5She0GoMTzIBfJddEgjVRZfVIHeoTjJ6nZW11N/2D/gnkEA8rWktP09na
H4BAQxAlKj/RN+Zitk8SQO4gRXRPN9W4w1o/B5b+Zz7JSBdecKCO56MNfgqFVZH3gm4vA+DmAqqg
zkxfFfusV4X2lpXdye3vH7+lxGsk10/rLIbyLLYumGWURBU6fKRa1lgvrWPJQYcrz8xRWeGIFVo2
tad42V/AFuamNgdUJw8IKbdD7z7si9ZRYarMVyIe8Zdn4K4wsgFykypVaqGuQ5CjrcQTmq/2516n
4Qj+7ClCSswUP9ERYro7/iOf6Ahv8+CJ+9yOuJtVBhxhEDWstHpOxTZ2l2vJ8RYepTm/KxprYJL2
DeCHFJ/2UhfQFm+SyLjc9ic+NibvEJMb3ykj8rFNs1jAshCyJJS2IX3yVS0hIe4WA7ixgA8cMgpE
LklzWrp/leOCiuqxzBeVmO+TG1HLY52fX0EdIkwgtT/9cWFvbmtM7sVAoie2UI+3aiH21H94soqk
4ii38gKDH3qlJ3MGzGKaOc3RUER1PGqQZMKqZvu3sKP6e16qhcgfPtriKe3qMR/HE3N143GwO/Pp
uiocCOoBXrxLdwpNvoba2/PDdZQtf5cdNtEpUt6bPJPNGrsXkhcKLjc5CYBH2l5zlNhOFcNwjFvW
5AtlG579GSGfwZCawJVwlEpnDEuxfAXlyh8Wqt69WuwSG2DLzeQUOh/NnLt//lW4dLY5KtGLjgHN
QmXUM00cA83u6WWHm1zn2OYAWUG3hU5zNhYudYvCHA2yXyVDOlvHB2Qu144iFyK8Dmq23REH07lz
Au8HoWQfhmCLUGVqHIVYGW7/Rhe2S04DecOgk5XX18TvpyJWOdSz2eXeLy3e8wHhMAMIBwgWxDiP
KC65sS/E2Qu7uS5QqdWvAjFich/SSoYQE2Byd576NA/mdxXoKmtc0+nxmTH36HC+GoYqWgk1b59h
brmFLYBslOmD7lWXwvMwpfBx1XuplyHTJd7JBrPHhZ7G//MBI5dNnURRQbxXL0xJBtoCeQVVb8hW
vbag8eVYLNNOhE7+AEQtWaadP0KlCcadJJE1+rm4ruWw3FIeftxJmFs1JT+4qgY52QRzEGZv+Haq
1qnnG/qywH0HX1nt7H10866UjFCtuUwegaq8mgcufA51AwA+QfRyIKBbGWuaWG8RGZvqWgjlzt79
LeX+x/UtJxJ0rYc0C9Yco9DMsHk3itBnMXHx+OkFsRAogmIgbw83///Im/sGYgUllzPHRsur1yS/
U5kJy+nq5v/yPmR7N9yIcvohaJ/4gmmg3uDREYl/047LH3t89FulQQx0z0evw1aYvoxzcRUc0pc6
bwP41V5QU5Gj6PgIk1bhvbJOXE88xw9tb2PALBj2vwK75Q3xhtE4KVQ4Knp6GIpecApvQvx8wugY
tu5Jj9RncHifna9pfwMOPCC8Y8a31h1rOShh/ddOzGUpxL4aBm/fTcT9zJ/7/StLnYAIdtmvG5j7
qLHOCgGBL5pHglZhtBDtIcIMF4hHQgCWThg2Ww5IvF+TAyOWC4X5psGHr6vCTsOUd3YfwZvlSlAM
L5Yvu38tYzjhLB/yAec/wl5eCTT4RYy6PWCN//1hanw8vzNXNOlWHq6qsD3NmE0CUCg+YbTMNDkI
1kDV+q6aQ8Ka3/h0FFjig/160AHLwZzeVmuWSSg+xeH0bWHgS0O6U3W19sAjCImRA4WXiD9EMpT+
LT6ZE3a4dsM/U3CB5XOuoirP/HwoR2CxFoN1o4afz/94H1HHuBQuLMNOPyPC2y6FvnqPwHiC2HyA
OxIEc1KXJJAFRcaI60V4TTvLh0GHbHysh8nWuOJ04M6Ml54tifsEfRjDTEkJqhKFIvriPB//m1Xm
mneCcgVo2OVBVEXuuXxw7q2sZPBPnb3c5FwcDwbI0IyuVGD5GoHo5UjQsavVrmUm4TbRIzRzkWDS
KSS0c5D4klNLOItAC/eX/P3ZEilt0idSU9fik1HBmXsHFG9hIJLM0JxDA5HvFF4wsUVzqvuVuclE
q5UNodutdSAbYhszyprUMRapDEGx2k1Dgo68BBb1oGDrrEmSRPLvzkebfyWYC7KEOUxn5+KdsZ5r
4t1YvtqquzRd4RMOsUx6KAtmqn+YrF6U560hYDcSgbS3JG0QubsHA2RXzOv1LsuKOr/TIu/i3U0E
99+jSKNru5nA7SFvQtKost2N1EITekZSf8fH/Dezx3oovd7PNdmTFq+ZbyJyi0NxcRZt88rAPEw/
IHlTdlEdtBiWXS++SJmtYNRt5ZxqMNVl3f2CLWQ2zS7e4+tuETsV5EXHsEkbu0Efoo10SPxAUJ2o
hPuDOTFoXwVMtVfa/eHOKzQZ1mw5X0vfq1+iOQt9ncrv4IPyJOudgtvmwXLHeqf2ncRRzamNHQNq
xXUR7MgkA4nqNLrTNBGHVIRS1E3wkR/xOYxo85WdrmAN4AjAr/dekNRIGNOAIIDEmZfphAIwCSEn
9N11B9ZCOl0v/b2/3EdJzJI+ahYzzCL9h5dEwEeMseBBRpWDf8olJOjBjHAQTGDBGlY5W48FVPbL
pkgeI7g9kd5EOF86xDjLnGw/3nIzuF0LMjGbxUldbXEdfdDqRDACHbh8qwKfblX281IWWVhSF4zx
YudhMmNhFfl51qVSCeEantWVPH/ReKSjWixkHM0zq45+rJeviqnRU48xqYwqrp79/pZPHrWmfeai
7ptDByNnlZWVmtFyrm1M91J1kznVPHjqms6oIxdjCrhzFuzSFGcZkWkbQwaeBXjwv7wnDXJQdiZb
3m4mElbWZ1Z1HJTZCU3OFPVQLT54x4i+f4hifpgtvGFG3hkKWPF2VcLYsbv9n/fRvn3a8wmqJxq9
wj4sOtBGm2z4yb6YF9e8DO0KmO9lTShBKl7pcNXUVb9lXcOA3Xw+YBijlJ5v5L+rjQWXPRs5cMrk
e+gyrkVoWwWcviSWZQx+s6ApAzuOMzNtwvxL0/bKjisX4neyLu5QBrxeZl6rhf4eaVQGipP2lFXY
sDuSJNwDjxcW0jOtkdK/xnHyNwx5yK3n0n5gXejyjxtYmCsUqoaucir6PBl137zlmPI7MVAZgXHK
+uOWOMZw3jgcEZ2eej/EqRYWwKFYcVBDSnzeZQmAHWJqWLmOahxDkTcRDiXOupwMsr0UQIGn7tDr
9nECJ6pvfuJS7Jl2jtx8wWGbSqZOb0yTEFYxICe8AN9alD09apq9+l7slR5upgHhqJpuPQv5qPYU
YP6J0Ad272CvjGdEdGfe4V5xzEvJIJ+oUnbDN510/qpV4e7JrtiasktXsdL/h6VTWYD2zOo0nT81
V6QJ9022oJCyYhiXd+oKG/BxYW5SfG/yk1xqzqXN3XDouykZEL7ynVASsZLeVX3POA7PkcnetoMt
0RF2JA2Wpl0w1QG7581xoxYeOYbFfrnHS11nq81kWt1YaGQXaHNjbSv+cSOPm11Nx2HQ2mBg1Xm9
DExynP+0hxdDx50iO3+Un7g887Gz92E5DF83u39CwGew5mrE95XEP68g003w69ow0St6EKT3zzgb
UQ2+5Y1Yiktzly8ZQvrCAzmXXhWdyBNaCQI7WtOAixQdlibuhnsoJ0n+9s5R86twNDBS5FBDjEpl
333+J74db4EO6kmq+RewSDh/GExyQQ/yAUZWdwssdxMFEc6mam043FIyls8Cj6GY/tu7ylFcXdvM
OeemliJhxRG76MR99PMkxDFJB1DxYa7FybdAJ5lksJZGAuMR1pJHurlS5nbJhPgeG4qmxVY+zVnu
Y1/T+jrxKPO/RS1S6WhHvh58YSR+3EY5ATX0RmTZEf6sn2BJErvcIjsoZ9s7596KIVj5icuAP2uN
ODNzwLBk/srFgxkCQ/fbscRT8P2T8xFJj9EBAa7tEOBAzDYdMViO9mrT4bQfnZguFSDUQNrhnrt/
BTwnRgH2+Wz1KKtlaIGmK042bM3vDDZKJDuGD1p/ONPGcvljaePmIVkta9vTmj9lztDfDaYUFW3P
8PWd87dpdhMepvYjqkFze1/CIP3yFqfAQ1yqfdd63ovyx0PhONTSy3dOv2V9GOJJrDelSlaF0+02
6JyF63C0rP5vha8lLKn+epDciQcKyTZgQYV2zjDE/OQkx2hB5e6Aud+b16qq38TOiQ5ukxfqEpVs
0YACPQS3jka9k6hJsdNODBKDYuBTYoeAbiZYjdz7Q06sPpNAVrtZehI8KwrcLdgcW+okxVT2x/pA
dCBQmQa0BPlWOIt6SVeb+GSEc2a136nyqZQWLsk7C+VD/3JyduTYz2VN6sldR/tpy6NYn0zFQi/d
+OhLl5GVm1mCBn7BIFrInKAEuHl86/zF4EPZBqBNj3aSl5VYGdiB5ePxq5/mAwux+KeYxWHJ8txY
/vJulMiaStXkfxducXafT+RORxa33ngx1jYZw+JrKCudJGcNtiU4QkuARVzsBuEHGPAXZcG6o2AI
ztNLlSf2/bL4P/1z83an918X+a8ZV7CA39jzTca5oDVSYqZ+wiTLCuwwlsbNFtaG4VVtG5xYrx9W
hvURof1nbZi2s79C9u/8KgBoKUPSvmQf6GzhDPpmmfQWXgoQQMkjGo0SjLIL8UfcsbGkSmR1UROf
yye4v/gVF1LIPbJ4rgF0of5qextuZe7s9uGiKi230BNKutsvoUwRYKOKy7lT47BmvgWCPHZwhODz
+x2xLvosW8RvGJEApoqt+XWug9eEvhiT7mTBOQK2TjjM6K2d9eCfHMWKUGBicfpHeMi0TXlssmgR
+sebJDCBy29gbVrK2s2HfrqYvRI0OUdGFQyct7odnwGyH4+C4+mZOmTpZ9xE0SNRsdlTN15yh+uz
rcKRzVosTwzOT34YO0wHRzUI+0pbgkvftH1qzV3eJevNx97jFsXx0lgV+ubRWcdOcYgQT9D7Hekx
WTpw9HNAEYwgCKB3pO8Iv/nCjyJ5OPwhIQpCQCrUlHajrR4jfKlLZkXtU9B7q6CmcVgeCNVWR9Lt
HqVJ6A0iNlT11hHILdVmgLRYSkaYpJE1HzQHNb2QqM7my3I8sdy0MDrBY6GRgoDn/lsYXG4xD48e
1mM0RdfOvKaBauoIsjL6JUg3d+GmiGxtwwPhwkxgQhIGLeaD6FJEmtssZnd1Df5itCoR1Mvj6WQv
nnQlQWwCsk+vmld5P1wjxltTRXOSCnvfW8q7Ona2rZPHORGHH6bZ2p/TWZ0VTNTaQ3ad8wpN1+dd
VjVBUUN8KXf3+YeZwAMLtRYr6GJgfqAq0qBIonWPwnJCxGI0Nno/A7ybF70zAZADFl3HIzFXoAeP
OcFAoPAg/cLnA+c0Z8a2m3DIhCyfk/xoCQP9dIkMm//hvOKsdXWaWr6TYoOedN53V8wWPqHVDyXa
FUg3y6DkHGtVqQiRiXTR1tlJTy44igeuGfwZCGnqH9ZqK4Vgh0Zb/twMlAC+tcNXKGch59xEli3T
EnBWy1QEfVUViDuahfC45XHI4DoxqlTiitfnPXDohlATzuUNzz7ljr/XxQ28WVcNLuIEOJvzm2A3
Sx/FKoWHFHBw4/cebMLDgJMr5A3QTTIoHiB8Ehr3V/O+gp6p7yLr1wlUMTK32kR1aiyS9khlDZ2q
ziIcTPLWGBuIXSvYIUCdrbN6JFEGPA6wC/SLWRrEJvH97vWRQZokILUItkSMh/6RNxdtAlAiQrrs
16oxll3unYFdjIRQgBcrYkstbah+k4ESvZ4y3qLhxkllYqD6LZu4WLNQJbayhFo4Ve9vuC3uw5gT
SravPYz4asPC9eXjomRx/JZnbTPwlrHTOKYu57wTjFj9SlHxZL3zxl2czJ5pNOAQhtoK/Q0k1UB+
wm49dQc9JiaKnRDccx3Q6paaUn1byI0dXvLZq9ax59jkuavH7ZL5c0su6+Fu5bPpojenq8jGFUK1
aAccrVORAmu+MwbmCUv5GftCjho9a9rtRyTdYBse7tOGR5RVBZ1dR9wDjWXS3dtPLTdT+aFOOSlr
L03ovqnKlW3oQuu1Gi+Kt8v5TyoKsbNMRJeNhI4ioq9KhxWTPCmrLDcXgwN7cVHs0tFcxDya70S9
lMa/u4GdxyJcKGmclIwqxbObwN9cCGObFYBdd9UhDT7sNmlhRCary7ReK/sQemJs1tfogfZzwvdB
ph3+VpxLRZ/9Bt3AkwqTE2J74n0GD+GxjPZ2kA0MBSrpiYxtp2BQpF+bKRmKBVFUlAHAOz3KYtpo
ZfmNiyZVy3qoI22kDPBYXDouPkHAf5WXkmkAHU99gdr5n+PfDrcWGA27r0gFr9cg1oX87T6n6WFJ
D1fnQtLH+BgZv+Yxt/kcVIfg/UouIx1BI2WHbyCXAzs20fd8X/WKTxrI/4O65wDbnTYHr1GttjWt
P3OQqa7sH/OWsP39Dh7yD4r8kCZy872/SRlPoHZ5C57gKtOI7XNebtKw68W9X4nx/d3b1BqJBC4l
amRKuFpqvDr/jD+ofQvPtgR6SrsKYcttiN21ALuiUQvb4RKypL2pD7PmINV7vvxeX2lxVwg7bw0G
NKlMOqXHIVUB0lDAgR9CzoMjjekIjIKo62lPfpkKIbF4cNbmcvXSn//yBne2kC+h586tf2oMfySm
NX6f6rvRjm64852YXAMhs9kk5PlFHIk70E7xWx+5yKeHqCfNcinDpBVZmkEcIMjoWS9a+qqMtehp
dVF7cJt76tUOVh4pQ8Bik2eWjxovUhWDKBQ0PhD6e7AmJjhtijPdpklT+T756+848URs7taZnOZj
JqoP4u6LGOyWOeNEfeE2JX6IGT1tUIqgGrZ31Yudq0m2wJm4iwHKJ7jifWYyWpAJbV/o0Fv/YzZ3
lU9deHAnoKjS9hxEXNfQS4nZYqEH1YKpQH9tSYTowF31pbzQuuNXMr3YS3/csXAleVGPklUKTnH/
KrTi9HLpP8+iVwbbrd5TeJ+zP64R3IROXLI95hySSE6MfofQnCipp1zEx9hGNYevIqTIO5bW9jdU
V9WXgppoAEKPcA5inshVKvMflh8u4B916fYE5TDeZdoVKB25GFNByK1HwfqpGmdX2pbqhEmTnUK6
wUILKaHE8qtcFp2ckF6zjPtHdnxspMyaOH6NeufXGEaIaOGnGcjUM4G1LjDQx7ynWJjzDGmI324R
IT4zeE037o/YIjvq5HxlI/wwAOyjf+DRbKb9YbIJTtztMMuocn+swP6IhHkNNiEJlMrg/8wfqspu
FMcTxb8q1+TBx8WkmsWh8NlVwb7pyyx+NDvi3tixzNCUUWbsp7d/1D/3dpQvi/+ZgnR8XKXcpn+c
MqAG6QAF1QpuF2cX09G/HjCfEaH4En9Yq9cNtLyUZRQIafyKT4MfPD7VWhl+GCZfvSRzYcUoUTD4
2B0IDyy7ExDWT0rrHWEMLNcb2rYUjmtaZ8zaa6701V/JcpebPodwQl/74zshw+n5hqAUADw7Psu9
33amGlw0fzKLfO/KeyqBI7SI43QXnYo735rnnJ3G/qvDTM/EOVnQenJ9G8A0Q/qIywYMapeSB7On
XoGN1ESHRauoxlKZ92p4RI9Bl/0EyxUbSjrgDl1TDoehzWs3h/p3lm71ms9UWUFa6uw+Cp2Oee/G
id+scvVQYfj41bD1jgbYWmoPUoPke5oDR9KWEXgWSFN4NGRLSAww6/xizSuCpXsKtFm4DvTB65C0
p4gTFAmni++cWpb1bUzijhFqWDTTYRoZ5QdY9y+L3fBJSpjPVw/Aj0UQfWCIs/wT5V7SC9GqYgbU
xDdLQuWLqiByR5tl0vx84Yew9Baa65Y8WppPo7Ns/E0O8RpAN/e9rBSjI93MGOJvUu/zFGgnpYoI
yLj5/vZ05RxlkSt3LLSNbOmg5LB2cLFrHqcPpkGxsxtrrBxKcPHncd+F23dbbbvyjSVl1cMLc9cB
jnZyQ9usX4nmlt6a4+pWCCv7ujKdtJ3OL/RuT5rL/g3+ZGopjbICeQpXanU9M/Shwpce9VYunBsK
w+kmtDgsAD8cB9zy+1NifIEG2Vbc2EqQOukK2U14DzSUbXG/mq+Msxm8wILJDBjAdgOi/SK6Gvvy
aHdon1RZWYkUFsa0zRn8T3jDptWSR7NLWu0WV0PmPYzv29MqtYGaxso954+V8X78JKS/2s5A0K3P
TUVrWSX37GBdOzcQoDP9ty4QiocB2niiJcwukal/e2yhrzRm1SLorTUaTV+ogMC2X4xowmIyBf9w
kvT//ykIV3xaBxEjwuBwOW3iHtcc2hHTG4i6+IqxfKdg1qN10S81Jk40N1TgvAkLizabR3zdFmlO
S9PO66vnNTuY40+y2AFGN8UswerEVb23wvE/TOFeavMteY6VZUQJQahxa6ls2oUHQRzqvaiugmt7
tGwn0M0m4KWeaPSe+o1Df6yi63tcrOfTz+GsmG6DiZZX11gzf7bacGsMDngBSSpcsJ/Z/fIIXuLl
94rqDy98TpPjJR0zBJtyPOtguUfI0avNY1ru8lSV6TnFREbQOj6IgqoYr0FciAb5/y0XcHtai15r
XnRJ8l+Xzts9VgLQ0INuvP4iBUNp5+C17cyMzV++ZHKu3yBI4JXMNXg6Z4syLwUoMLJ9v+afJ4tx
68xVpyBxBzVd1VJJnT+nVtuVqiHHrNE4DoYHHR4pGKij1jkdh/eEPrHtY/xno/w1zSljICZ3g4ny
t05KvdfXo0glRyG6jGvZDz0yESDQZuUmg3zN3GdnXGf/wZG7KF+CfDENA58fBpy/o9/LcKfQC8M8
loZjgmztXIGdzojf5oTsRmbuAvxnzIcRDHjKzaL4kZ4GeIsqQ1DII5BqX/mQHDqwupttTOpC7D+u
b1GxUBhoaI7ajokb/Q0rSiV9rP4Y19a5RBdaTW7dmwbKw7aoME2z1Rl/Oe4tmgcJZ2HFMxFRsT9b
m6Jsnhdupila8Zi+fMAnKO3ywclplc7eWy3h8xkzwLU6xdK4Bv3ATK8YrgWtHfgAMAfmy12Kq/Fs
UlwxxPGLw5HYFSa1t0Iu1nC+1CEo72KF0uTkXrB0BW4RlWRgQ/WVFQqLd+lVI1o3hUCduhBZlPH4
7WEAIjmXl7Zp94J0spNyussySV8coxQFF18JmWIjxD7CYRq8v8umhhy04P6x6D9PembFNlVGsn2c
5a8RjPZHeUh+8s963eUcHxEnf36nq6hVN0WWT9zJuMW623bV4UhGCPOPwUCKHkzzRTH1EKVqJ+Mw
nRgVoHK3N4IRvohBSuPENqcK7Pta5b9kwUh9phOsDGhjHMScDJTQXfY1X3YURs7/5SZU7bVVTsqq
LQbkA3+w+94q4K+HNQ8kJSW7a5UYSo9eEh8TIa39/uH6I3KkDpuhHSSphlt9d1YeJXpYZgxVpg79
pKciqDpwPtwrjiGnEhSLq1aXnctVAeR9ysqGA0wGuNfh4uclcP0HarC+uVBFgLy5Qgujw9Hxvz14
PEUbORzLr9Pj6J4yyePRSSU2xJn5AP3ldJEjUYZNOSTKZO3PyFdLYrZoQAYM2CCTpAj5UWrzGaiC
Ri1U2IBqisI6Fq+Eu6h0CWdva8E5A9bg7+ZHoIomgZmy84/8MpVY1ymCUSzG8LnILuUtbWv0i3WZ
+QMy+tIHIoR8RSfEr25d7fQjyziEHvPa/9RAfwiRp2gzQmlErZCXcb9ukuZLQJQi5PlL3kjF3PWD
kYR+qAYaehnk+JE7GMa/wQb6tl9zJzUQotM8By0UFGV5B/6SASdtYF9+s8VPtLurgsR+NvDvlFI2
eCYd5KKJH9RYkVWscdf5BSeq356DOUMxYZRT3Xmliz826l6Nz1IT6SvkyKVx1ySR0iMGaTy8n5xI
DGNl3veU75JsyyFQjBuS0uSKzL6//oPm9koJC+fxJ37GA624yppN5FvN7T3lblVWDpatin3EzhhV
Xukh0k8vrnfhQOT08lWbEl3a3KrOKguiIzCVxcHh+TyI8v+UFHoFdhRgMCLndM44iKTuEpnO+59F
VF0GeyaehwRVsIymtguUg6Scm7KelbnhPxAazQ+AdmpRr3o5uxWgHOpNxrmeEOWd3AYxKXatzDiP
IcefcaFl7cqgfKONgomJCWIkgDcU5yhXCuDjSClaR2VwlVqCRjD4KmLAHRo/8alvcqyQlzQyYXQd
iDqP6zE8HmjwnDHgqk6+Mt5BJRvh/UwLxF8/bV3h3aGx6lpH9+7l7hZQF6AYxK8eHw5DS4W091xO
QvOB7Ji2PmsFpDoPDAnHH2aZLFXGC+gAM8Hxkkz6Dtc9K9dpLxq5KKvfAymaKcq2/RbwNxscCTay
iW9gbrG077WGOydWMMmFtNt/W0/CibjaruX2clH7Zl0Ew84GXX0J29A/Y7Udr9lEag4v6rp7Z+At
nBG3cy9hHfLwqAO0a4xQEKWQZ7cOS5iNOeLBbNPWB5mZ9G3rI0NYb/bVAAFUa+mxi1AU34/Rt8mm
7E7Q0rCp5ECaMQPjSjUHoWeTP7SP9vv4fvm4Twmmr7xWEj5GK8vaimJZXsS7Rtt/EJ1K15I4TKN5
lpfLpt2U09r5aACZCPI3Od6eQKZWvdO+eq45KlvVZCP3Axsn6Z8SSwwXo16XWf4SbkfDTH4868kO
ql5Mm2BxG5qwM3RiG/rsQd8yEAQQO1JNFdKwSsV4j7LU55VVVQQ7aMUH7opjXAS4uv+uUTdmD/EL
o9FiURYgEizCYDuBxSYanSQVB1smvlEHt8V/97Pz2nS+6m3zw3PN4hvRH9IhYaQ2DJHlnZWsj6xn
+gm5Twg04ECwTafUcWr8FJssH54pCP2tpc18qAccBEjA3ipYHarrJVfUyOSnpODe6wWBG1OIxkwn
bsqRFFyxjJjAFnn7nzgOu9+eitrnILCavXYowDCxzyKsxkY/sVnfpT0FuIvaAI4kOi2p6FdPnP9w
aHAFK5V1HhfweMj1wPgk+nk8xgvNNNHqXejcxNp1CDcEmMxLEtPuW/irbcncGe7zheQz5MWvUvM7
yZTPymHLYxywRadV78+R6N2HeQVdSeMfrQQ2iaYsYbmhi7LsfOc7PWGF8olPzAEWuo69rmPqQYFh
vYjzT1CCfSrlzlgHrdY//KeeWPNMhGjL9D4730WdBt1JUmlGZ3Y4xABQ8PC02zYhF1lpjoKHSEUH
3iXBUHOAk6e4HNP4VxLXbPd0n54NKXHxOH9cMsTPW5BCpxsHQp/XVMuY2eOB1/C8t2twk2QHynkb
drVt7W+g6MW/HT3XNs/pmzIHHk4+rQcFUuMzUZPMxL2TPHVGDStpVYDzp+8DTlWmT2ljl8eKyaZ2
qdB8ojvXeDkk96Iy0hvn15H0Em3zaXlut+jTEu7wAIf/quIGfzsyCKOLOgfN4ZjDJTlsUU9EOYXb
SkZAs1BHgawAdvvj8B7FO0w5oXuD1PFRVAhtHxJEob/b7Z5MH5TjAjobwvMGso/SVUdqYIF+3d97
jljV0yxsueCkqRqUJr2m8uic1IrH0pNN41cKfxv6afe6wIx5rk+t1Gtf3hP16GJGMkCW2KBOiWh4
vfBCeRtz/tIfBfWhe4dIXV8MUH+t1DCg6W38Yq+bo0nI1m+b/uqUqXq7ToD1jzmdEJkyJenA9q9v
F6NoJ7QkK+1NPkmN6T3yxQZO3rhc8fwaL/dCrDTdLz19tcMfkrQpfV62oB46miuHwE0E4btpRbTr
jWU7lJVXVNUJkQ7aJrUJawFxliql1rJ8qAGPME/NCcolSSWozlYemEfoAryvPw61Npm+mC/Zpf1k
35H5iOF3dOsBNZPaHAvQT4KCxZd1btuQRkayXvvjWP1QV9hAs6WR2TfAPh3Jv0d+McXdpypzh7+M
f6TZEn36waqEbB4ivxzx9+/qPO9b3KNeN2pWzWAZxgRD5epdYJiaMjN9ChgpVaCKC+Rl/2vGMTTM
7883RJI262eudZSHRb5GmFmJnEDuloxtuO16QVDyDtiu2k4e6U1SrxXcLsTbf8VXGBwPE8Xt2mWR
k2hdcMMZf9mpSCgmvMO7aR0R2S5HrCBzCt3icHHIcwQPxlZxOnXgp6VZQWqYADJpyMu2KWO1iFtC
93qMZI8cmPqskuFgwm2bvgOe0ceKCdstR2j2gqHKmxl/Hrwwyj3YU6+nJUk+D1oVBJXT3Nn9MVdN
uQpo9KLN6s5Mn6rI0b6Nq51FO9fskwZB85VRp88jwpzh6KFkizd8+RmWm6d6a/u24pCWk0fyXwtP
ghtYWWiQLYuPP5JYIojzGndz0Ke2rW6Jy+6dOURWZYt/Rq8ICOpjeZ3/rzriYHAKKejHG17Lh19/
M4NCCmcoXsSzQUmIukqvlpA9tGmhHzcPmxhw/yyiLG2j2U2S3L/FH6BvyKoCK/yUUse9c+2jd1aw
vPGBJVP9+6mwg2xMPmNFIwH0MG0YIGmxiKrJof70f2E97sBLMjjhc58uqOeoL8DTZSG3LFlIaEaJ
JHRoHW5++Dpd5hCz8LIGO7Lg/0na7gKmBZTQFx0V5p7BHIq6MsKrBM3UbunwIR5/bj9vhQIASVaS
LXIbMvYtfKS7VUqluGvB39lBpm5s0Wn/sf9OCvRpVBshsCRMdNIQEiXbzAGJMH5n8L3bQNw28uab
40Qr1aRnQeZvm+zaEvPbj3oXdshhsifoXf0nXa0PTsVTjeywcmQqLLAeeUt3rHZjaLV6088kzdtV
LaN7QeLA1RIhVlGQ/GtL0EZ6bz/2dXUTrHwobkbzcVs/7cYpwM0o9BwdjXEuLMQ2HVEzsim0LKp7
JT10DC0WpHrE5mSblPyYxELh3OHNZBRjV6H6gKv2uPRlGZll1fDYzno93cYQ2LcvRIHNTsQMvJBW
E0YjwOP9tmclfLzn23zPIlx1VMQky1iugkvCivYwbhf0tSRy15vkykclirj9dJGOYSUN9PGRzbP3
vO4CzVmynDtGSGx5ZYj4MGvxMWwLz24SZ89CYzxLnjpNOFj73VoOUs/EROjM0iZ3YnVgSjbyE6BA
WjcgoC3EcypxF+rBMU1MDHUYWOeGYV7fD4n2rtFbt9nTS9HNVTewyc0PgoFTtJAFVcxk3oX5CNto
9fZcmW0iRmNVhThZyLZPa66W/05agyU3gR9orIloXSL7wF34+wrltH7qtlYKlzls6a5+HCjGpFOM
CcdVF3sBrLb3giWWLVJrPX+x5tczcpwfuhnQca5VFaBXFWvwgrccnFHrMv4EPo8SURV53ihkrj8X
SNjGM5r0G4RvzRMBiswxokAGoG1KGz0yqDjRAt/4VKa29lnx5zfPBU/9lbcHTHyJA0TNVBSURd5k
l9pQDrOlA9mLg5XRTbFgYWWwxMbMUHdhjeGmmXon4RBzO8pHd0bQ4EsVbHGnHMoZAm7b3LKFX5X/
j0YYj2OnTYoShlbwTy7Qwnq7pBHIt7j5b+2leRjIkPy46aVqgM9ViU3UChJwtgboILjRMewJXUlV
42FHL5iBNRYDHAMShcwEpQaXBSaIi7kTBCCNHaTuynXiAM1MLWHH/8FZvgAiGpqOBTMtb06ucZJS
xvkRHL+6yspG1WLOdIw8nA598JmnscoQ25XQNLbTyRpJw/nvPfkF6x5upg1ns6E2xtpWKrKCNFn9
yNZwX8xsPWIbnuTomMO/NkHqXz5zKbBHUAwin6YkkxE2knDWHHx49Ro0r3u0HaBtLBI9aVG49Vxh
Js3L0R7oD/qUoXDFK1dqoQqOUUbgQUsjhT5v/jJiEv+IISDlyBSJmwTpgm7P/rlcM8o6xg9+EzH5
jaFmMzRYkgYKIYs7enhRwZJ+uvTOiOBLLXCH+wBS9+p4lilV1/vIIn7X9RzeSenb8tDtFV2XdhTS
zLfollYU/BFTmraEK4hwF36mmViXiUGCorSv7+hs/rHvgaANrBzKJYiWL/DDs8msYvyQDykPayon
OWP9PSCnxh87+684mOCuMoCGxp1FCIuKyBvBLLSdfkvi5c88PAIzMXPaTVO+f2XX3QqQ1pdtON1a
vkbHvGSFgZgW51Xw2tGXZvdXJt0BjXKY7wzet1NI/ODDFZqZ8a7XQC0x2Wzu+szIDFV+Y05ao3vH
DtkSSbWzJ+ejKxhVYT32ThBf/viPgU87zKiJVrCyun+kI3G0GFqdtrA0iDi5BuoIVH9LKTLFIzOq
k3PK/qqMzOGR/6qWco6C3GGr8yLGqiqr/qzQ5oBSHEWBOYtmS9R8I00nM4P5HPOUcrEXzf0fO+cc
JkHKXevesYWPuGB/UniMWX4J4AI5p17CZjntSiTQUJlUP2M9K0MlwdoxVHKYAjbfpjMQpsbH7dzz
S81Swk3Un1OtjqAybGA/obpnD0WV8mnF06DxbtFxdZ1xtFQKPbNEE3/3smh/X0+gxQiqxBW406zP
DWkN2fCnp1CuwTn3sbALFV1614rNlWd7DUBGbQbeYuJguUvUPspX9wL8MQ9oLG2WwIVaPjRDQtyz
pcC79GDwGi7PicROqMv7YXvC1KJBM5PmLejAtTX/Dve9RpHJA89GrRZE9GAwycFXTQM2tATgpdBL
FgE16IpwiI3vBiqwY7rG33QmbaUygUNx3gVJClNQC05wvQYjZNozrtqZ/+tM0f55wJpL6Qn2nEDT
wAnIvin72Y+Hqdl7nCFaUHBjRyQIZk8BRPKSvEI7CiJPiXAxJfXUErvPkTuFVoohtSOQy8haEvyT
ZhcPffLwo0N0VbqukNTGy1xo24eqESVXoXXsf6WoyeiVuvgSpm0DGOcfQssveV711440oevvOk4z
Zd8r9Z0TzzCJPoodxvuT6GvSurMU6p8y9YXBMVqIwS3DBxbgpPZM2BwtN3ZdA+btq/CDjuT6pXDu
xySXswMGFBc2uXzVGq7jol9UL7VR+4tnFFRQJAA+Spc92OMSlw8SAWMTSund6Z906pzz897Vwq8Y
tjAwOqaliW+yxRfqc97lFXD/abSxnmeCRPUcsihqq0r1qPnb8eDJPT8iE+5H1ZC5oU5cCqc18RUw
EhQZo3HnIs68agZY7Zvn8rEZiGCUsi26y39M096qtad9oBkxAX3EV4CzHLxZFc2cD1X++vmOo6th
hlrfCHadgE6vVxhNyWo8JbRROcMPUIUlGDjN4YdDkq7v42vkHJs56G26hnxndvueyDbiEm6JaRtw
lXdzsdjNNCHvxYf8v6CCwuOugrD4yJbO5M+Fz1kb6nyrmxI1DR4cZZ2XzVlEthD7oi8CL4qp5Qc/
tsPhxNGJVjwtrGOHtFaHLipbuuXl4HzRJrTzoE6oZ5afFRMuUjl8hrI+Y4p9dBBjzIF7qczxUzq8
+lsAHhacPxC1n6DBAMzar+iovGuRIluGeSdBKPDtbGnz4kEa0k1wiu07+nvWcxde3vsJ+3SWeXFQ
qEUiumUYehysZKT36aA/Zp/cGaJH8j9WE/B4d21v/R73IwazJToAz71kLYZoymLyKGuxmFFv2E1b
gxbVxxi6saET9kfgrkWuM5FFoNEfQn6LJJdSZdt8AX0IZndvsoU2eEBZAyG1G1JnTJBrsHvOJhZe
enO58xVLlWmfuZwGpAfuwT57mGZMEF2lUycxqVSSgN0PX5p9eoa66nsCF9VGDI7q9NPlfe1kLNZG
z3KqoXAkeSwE2987CuZxMN2+e2I8XENrLOW448+4OJm8xd+wHnBaJFzaHsaUKuOkU8FnjjTqtYMc
mbluK9iA+4iAZm3Q6Q2hWukF6dtG9aMMVf+gu0cPRfy74yXfjXjFdIWl/rFsQsLx43DTLkA2Rw5M
WVc5lwGLdio+hrIKa8dB5fRGhoYf7ggqd8TM4xCxFcYonKmMuQf/oyPsoMDJck4f8ujPPPZDqfT3
CIog7is7ChCqgC5L+XnPAAG7AeYua1alYp+T936xjUhZxEjHnGDSZvkqDNwzqRYC3mDUSXsQLN8+
2Cq35RXOqsitAzy5Q4AyKrCFZnxPHeyA0QYXDFHAY5wBWVga8oVT9cYnIWdguKuoE5NtbMdW9YeC
sN/L3UjNiwBfIlW4E/SMEWgmPUaJ8GKkQLgnHzmo1qTNc+s1M/kf2I8/L7pfR29adbdjh6kHFufF
fL6eZEflqYaV8EVPAvnqKJie96ZfIY5/IrBRt+plfBOq+e7rNd9esxWboPaEiP0o134vxoT8NKav
i7UZMfFmG2peUdRNDswNBRP+CYq7nCXUlFQMU5FL0OG5tcbg+5WmY5rnvDyvvkcytSGHdrk2TZR9
KN+YQR/vS2IuyexUU0a8yFKO5DE/Byo+VraiWrZCcBO488nfOtdEBpHZPMyNx2dEQ+Dky6iQcRTD
6uFp2XFQ1LgiI/AEQtNKCAvzuBsljAcibepGR4pUOmo3BMvW9lcLQ0pg69+e6Lel9m9agaUaOVDU
l9oaTjnJxOVXDW88C623pE1qzqQOdFs8Z3LmOxXpepQA+agrLXg75alOB8Js29HAxXofJpyoILGd
kBgwqWCqtRmsi+e/1jk/eU/eDx6E0hGucisGO5Q25dpSAmX0X5wSOPxjQPeG4ESnXJW1fukf+WYt
yb/r5C5DiiHqb6kHC6XgcMB0UAj9CVIZFTFZGubM1aNPfB+1ztJICHpceSh06C7h3aZtSKbEF2zX
iCB3cWnIA0oy5op4m1MDlXyS1ZHnKc+8T3FeTw067LLUR9OTiGFtH2xZrCaTTc2LNJ2ca1CxoHEB
WlNwa/HQz9BSuJ8zlPEWTxEGBraJ4Xf4kwtqPW0+kiYeJU8lJTrDWK13Gfr5A+rW09uF1gfbuIrd
WQVjmUCUbVeTW+Hut/AoUYlHBhCDyoDhhjNjgxTTjZjCna4vblg9LtsYairUv0+WjBkAC6a6ZCcA
sPrt1bmdQ227fcp47Zt0snN0FFnddJF0JoPXnSZ/1ALrU6UeQ0kHDj6PTsQLWNJVTfot0cPh/x94
rrffZOGJULfVPOyLXmxHh4Bc1WH4sfApWyOxMhwcbUT7kYIOniCtdDbYOARdqKQ5+EyD+muQC4UI
cfBZLoVlx8B65nnVM9Ny1i4cR8BrKCGXWAgssC5iQI1VKmLaxgetBhntAe5xMc7tbpM2r8wvhr+Z
PDFOnEnMftZaLkxw1vIDIAPHeFU0VIMYZg+adzjNw9AsUg/C1okaoi7cEvzhM19kNjkjMZWy2mFV
JD3gAHIF8R5TEKoC+HU1xORP1PQJEXkSBGkc0PaPUoGq8sQzTJVWGj2+ts63kSeVMzQJLQvKfWJJ
KQ3n0FJkg8sUydvDEXvd7lCzl73dfLQHi5+w3Snkfbjp6UoKhR7hwvuwwozKIxcTQbqsOAlDWA9U
vfADoa596jA5J+Rlun++GR07F52+wK8rnCaS389aqR9t+KK097+HiTvgRmlQBIuVDD/j6vCswghA
o7fHsEhVUB1zUyOFMB61SE0CKL50QIUzWJULMQr1MY18FPSdvgYwwumrwXWGg2PmZ9HL6EzNhsLV
9Z/9NVwCsLH17GkbPeHveBeMpccRMM9XnYXa4ZVVUCShqszmB6OQDbrAULDHonQgSPjyiA+DoXBQ
KA5Ea5PWNpGCX+DD6P/koNe+9CvjT65RLhzXDgc20JqO/1XxF/HqqqZ9W44S4c/mdOJcQpjte0gu
N2czgiIrc3yaHEx3arxYG2iI0IkOB5Sa/+T38cQcgr7FOGfNN1+gXtO6rd2GOwICUoWuCUbkJ35J
vzpzBVLFohn3/42Plcj4oJH+u/RxLl7/krRh7Oe940g6+FROt6NGPO/IIk5CFlhig03cmi2UIVvM
aEEOj16AItTsIpCMCnWMDi9osBsjBTrKhZ5bjKdKb16m/2ynH1iWca6Ri/sDZOo/9uZ9XjHbY1Ra
dbLoP70PS22Qx5yUDghwrvkNOV5lDhRX+MTLXUM7dEl4l/1jh4u/4UrccoNtsE6lW7qENTEnk8Cq
0wcFFRCuEV1vKfQqobVI+v8BTxjDumj4nYdgGumz6ggMzRofIQFvlhO3DiGIDZwJNdxS/h7d4ax4
MjAdhyjaPI6WYwvTPtPnB78pVqn7ftRuk0//hSrBmQQ+JjBARjCbfF4L91ftssDndzCm8bD4CKR5
Ar1uIZltbzz0R3Rs0/B/4AjZTZ5eBlqykBXep+1fXqUbdFnFqi9DD85KjGin7ib3C1HImb329sLX
n4U6dk3KWfTGjTgUDph6cbM0kckl4mKgwCSAE+9SRYXM7N9daf6YrITYuhuhXY9JZzP86mGQeedu
IUypaOLUOSrL548UZycvX3YknCMpXQ+qCMHf3nMGtKHR5LLh9gTjBW+nkt6tygv3hDJ8krP+L1gA
FXFF6GtyhNOLoTvxMBQAP1zt5oy7uCFcRyeickspdMAiuA6IGzgK/ewVCX8NZLF5jLkR79w9d+M8
REdijX95oDIk4SeJSq8PtWpQIcmHSmurtVWKzwqOTyYX3KxQUGfbR9dwdxX4Z0FIc1TK+vcxaD3G
miso9yoxr2plj4pjipe7X7CQYLDYPSQxhkaQ4nHt2dJedR/RasMhSdmJDzCouW81j5tlZOzTmjvV
QQfj/BenGjSMddAfCf1GJWvnOwMQJFyZbiHzBsYU/6iSgpKmT6U8gqbY9r66OODTffRZkdyCz40/
OMRNP8gRrQKtQrKN7jGw+zv1sI8dlxhIT6Y7Bc68339DF5NAhIL6WGebVO2iVCRj1ik/dRuvqvl8
EtSpltcSGa7FRTVOgj+7s5g1q/kHXiZdcZqoCvG1l7qo9IGr7sdGRHRhwmdLOzpAHRKUk+IMAE3u
8CYavszwWSw9c6XVrJ2f9F0XD1XVXSr8BVc+cdlwkO8ACdlaheGvKsckzM4dXKVtF6QKMpESdQ2v
IDll/ve4CMuI/v7ZCGC77KMhqZGkhCVJ8Ie1nwLGDVFjnJDc7s/kjgCkjuws/fJczTjUIxtVuuBe
Ooml5OYtPEGQFgbq7JYeukXBclRuCIeBNt+e/L8dm3Pcg1vyBHywGVYK2XRF6wmXCYgtcFmz5R7Q
2SdBHNZ2umFpVpXgltm6OUznoxm6YleGvu42g3pyJQnV9uXW+domoEEEVfIuutA0mevesX2VzzrH
kqEf9xtnb2e+I1TNqeQ0oOGo58xCrTNtSyEp0D+/Lro/piF64Z4fE8oBNrm1KjiPJrtSaNyvR4JS
rSsI5cYK3fLPT9z9MJMknfGZGDaVX4e5lRVajTJtmReYoiubw6wzOY6JyMlfjs1fwjBVbEDQSKpg
5HiPHJvbXrIm0qlAK8qRFv58Nm0dmpqeOWeBeBX7PvLs5k25mOQsubVto7aZUXsHknY7Dz0MalFf
g1b8HqVTzcv8NOvcw7sceKGoO96k7VW0kXh1VEnkNyTRPImFLrauCqlFO/bnEnMwrocyZduFLldL
Hcunft4i8VIbOC4tO62YaKJMAFP5cnw78R7yEqTq9pSFtiYNvegSn0yuNfsbNeLCq3jznGvxazpG
aiZVIFG6iBLcJ4ATz6Uxjk+EBbVDZEFie4hWh6tDkxONatOSf/vdg2J9fPgtDRLj0X4Rgp7Vtk2D
4YkBt3T0nljSSALEX83Mh/1I6+Cw1GTLl6PtNAN5qykQ2yAd7nZ7Ca3FUt0PEWqYZ5+GRnWucHLv
9n/GiZzyACFpGTj5mWJDkknoEwJroWX3jzLpURHQ6Uv3jKSx6wzCHLiZjRIuvDg6Me7Yz4kbanMO
K2uI301aDTcj4AG1HPLiDCC75/nA0hnZKyur6KoA+gih40cZKDkR+C1eML4jwI6EiN/t9WQJLqK7
TzLtWFtl0WM7tFg86gpYoNtoMnR3ETUQAH52uY0hIuHAGI43CfT1gcDTykqc8qn0GPSm6ExTAlk+
zLogB8tYpmYsX1gJW4XVoTEyvrOK9by+7VI/VVPtVGWydB9mGs1lWltNO07gnBSpD65cAXkXPObL
qI2mrxMI/SSGOHRBCSIOupOgtHa89rMLtqp8n/bN6y6IjdpuI9XtCA7oyeN4ORjZbgMKWYl2cFXi
RCUO4a0ujvBmDmkVCCAR325pg+C5xRXVbs4sS8L9xLle9dIw4a2Er+y56xJMajRufl6UxaQEkmBh
SljeovL0Tv9EDlkknGD+txLCG+IsNIUZq5FnP5LKrXOm80KCg8xacWWz/Q67eimOp46zvwdKFVkg
JhLL+sALV5UPjF1phhCjxSbFYcqy2BkwsLmvlFKfFZxnbMywIzE3UGvwSg03KaJXPgxDQQevaxbj
WBRCFcjZHoWPBEneTDJkCflboLAZAyrn9ujfDXA5iRa5TAw825ap3lrT0P1sYhKHZS/CPGmH5pkk
j+sQaziMLKPFeemJOgieePr7WutFK9b18pM7obiUu0yw+PAEv2TgTV8SNZiP+s8Ms0HQXfpM0upP
g2iCi9kk/9EuSfyJYBj0Fjb2rkvVvp/oOSSv4UfOtKrVWhj1vOdC/qt3ak4+j8RGJ9h7CPAoQY51
WwG8R+CLkXNgpgLN6XBTcdghl6KxrW6mBjn6+/TPl1PPPDxF0mkWjhNMaXuAcv6+UOUnbilgSkb5
yTuyWXmIQgjW6lT0GBu88wSVnu0LeSc2yr2QzF/4690z7Mj6Ch50xl2OFCmSdMypHUQUShOILzF0
TYhwLKgIHNZxt6EJM6X8VF0yxQfUwiWbXKEbXB7M4Z4vzpvx1AHFajntwTW4iTmIJTu74EPFdf9C
/QCIoXWhCC99ixLc0h0uAy5YhHktIh7qO7yYhiC6aP9CVp3OF5T5H5S8OSjLlx4lHy6aSnmISsRw
RhUUzcB2MlMeBs3SH0bOYT5bn1pYq1c/z6FP8Hexxa+Zx1ANFdf5NXu56k/edlksX+k+ezN5vuhx
nDgyPige1vJ7+jCu4wliy55sb6jFMoUFUz4WVAfwQ3giWJ4TgZmAp48maVkEOH9oNj9NiaKWWW39
Ck+Vyuub1jfelYCwN86E9VTKXLf7bhYbQj5lCbI4XPr2d/5GDhFuUUL48f+SruawQgXcwkNjQ4w9
7xyLqFQvL1pSAoHo0hGJOp8fsJOjVcrGMFLsRqqt51eWPkJaq1nkHdVA1qfbTwfWZxlRxP7ID6PO
ixok9jDCwHK/rngP7hqO+wwbTEwY2/hVWC7Z6wJAL3rafp362aTTPabYtjwJSBU33fgdYKeMc3nL
51+vkEOclP+OWMq8+dTwDaPAWqqxeBW6qrJbjSeseMWXv6LQyFGtXsOYPFIzMz1JqBeRGrYiiZmQ
dO8u0e+ov79kBwuJdTeTREi/LnG2yj3kWqLvGVt4aIJMwh5M96QFAsyWqp9xYln91blbJ9QA13HO
19t4a6/LnGRwoh/sdYFPmMYFdLRfHUEp1htymt4kxGv2ZqK0EpVYkb+Pmd5bpP7B3Vx3r4LR7fU3
uVa0vIoedi+74/LMPZkbJHaS1dL7d7S00dzqnSQRNOjcJL4UbAuj7x7t9DDNuAZcuAxY1RjnuYaO
h83sMGj6LCdIKOZcagacHKalPrYHI9iPiu362kjS+Y7rMBRf5eQ9HNnB70QEDTFEWFx+nc7J4Efn
zw0f0ytvd5obEVETQbOWyZRjBSn5lmwXVu4WjeRfCU3drJYRtVmMWS1BwKchZsVtkRO+vJ4BxW+d
Tr7TP4WgV5ayon1lnISSEBE83dWGDV2XAe5tqscwQMKW16ChmRv7lpbwoDRX4bmiTjnQjWtdN/Ql
W7iBJNAfoU4zTU/yqBN+ZmXHoCHtaWWKVejhpDZxR/Wev8Uyx+jAFqkJmwCvBXjAG8lV7O+1opic
TEcocr5QLj5pwQDZUaQy6vKB/VZs7zQlyf+9EH+2AnRxj+qIIiTYKUBJwQKNOmmw5X9hpzKSNfNs
UYOMGuuCU6ttsc2M6CynNVsz/zmTOOqvvV6VF9DLwl3Z4hsuLLr2uIWLocVEchR/ipcRocma8dYb
rgEG/cbQU31eqcghPpeFqZqi70c6FHTtq6Du4F5xn3jh1Rp/wC6qlzR8lQFa+sroIb6Tqk+g80uY
SeLTru679J/WziR3ATOlsfywrmrUT6jgXIl2imzzwzdsfcgB5ukSfVT+uQsqDnMMtzF9VbJq1jG6
BPdGGNamSrMtebHxhegHr+agvey33wyGCp6ujrj69LrqEyLLrKI5NDsMSpKUUCMNWBbpT92JkjQD
OWsZtiKJDi0N33dDJMTTBlMrumkAr60jX0lmR+4TOy5n1YbdK1fAYvLRZyIyfh33jRz+p1xis+yO
1HzuquRAYzcQGA7Yez0e79/pl8q9PGnNxwGVepIFYwcUEQtuAYhpA2K1V05u8Cn8+cjstHjYdiag
cnC5BQzwLpEMlk9QHU6rFonyeHJnnPAx61ifFXYXXYpRNR7AHHSTRuHtzE8Aen1sX1emIc+JasmT
aO684jhihtPOmOOvFoJByiX3seWhKQyXdse4It1dtvo4UloZ/bz83vWXFw+eEJX3FB90suchkyIE
YBbBWBMv6rtgFCwvCmZVmZrhmsa2VbFym7eF9bgv2e+QeDpFFyVdtCfrkJUsVK+3Mu8ZlHnP0P2a
PXRIg0ni+nWZUDXCscoDYAgc/ehXMCkMfAH9dc9kd6bgAJFa/nD9x0ezETaFT6kEzry2X9kOIplh
Tc/koTTjnFH8vUuuY2a68pa02L9/Gzm49ZlbF/eqOmUFJB/g8PRCcVx/j+iIlLX/E5ZHyaWRCZ4a
qtbQEWMxSheFpC9JYtmz3P6YEhchDVhYXmCcqV5RGpvhZd9npvpi1en4wFM6Q5UmzMinJl00k3e2
wHwm47fDArCu05yCrNXsYCkdChDq+vkJF/a5BXl+OQ0695mbX4dSwLvigq7gxnrCddGKlbISu3a4
w13sIhNBhMNiQsWqX2PeQIEMuxbSYdDZQmUtTbvobaIn8O0X5DfqoXY9YYJnNWiEaglQOnqt490r
UnQSpGGkCLfePhPw5q9bEIPjb6Xold/0kvr37PvpabvKadqJ8Q04mppXl8jiXNp0HjCz4rJdiGvP
MUwicHckJlAH0uKLuVBXGZ1kynzSWUQ6nDQpYDC4Bou7s2NmVlrYYRRbbeOXxXXtQfMCHdLNoAAT
5N0CYCGvS+LsOZcw53CAK/k9eXeRhjJ0EG8uF/MtSGYL0vmqkCp9xzE2G3FHNNuRInxfijjgkOHR
U6vACvMwZUSlCHAgpqUjOlj6hEugOVmb8IKE2GoDEmCvTYVRDtb79YmJkcVccx86DyXS2M0JNhCS
s2fIBrXPr2B1yHiGg456xNkHXrXRp0NzD/naHmhxcmKi9HWWf8S0LeHhUpTffENHoJVoOToSClij
x+7b4GZUGLblLjyQ3XSu3oZgUJ5mDY7Kc3TX9vUW+KnBooCT5bVTuUGBfYRmzZrOOpQ02/WXU9TY
CjVFaaLkDia6su+6RTJP2gPLWYRsaTEg7EGj29lm3m/FRD60LKQw/cH86WVQCtzJaILxp/92xbwH
ashANtE6GxAgIbypYayc8jaBtRGc0T8n+JSY1gZqlO29BDuUO3jVhxHm4I7/6C9or6em88LT5Cgh
ptaKC2HIvKkOXD0iAHIJqA+cWDFsG55mBQs2zPI8H5uxPNgcszx+VBlBEYrRcvAspxs53mwcFGwx
XaUrTuLUYWNijBCQUToYsohIkX6gmlOlywXu1yltuPC/6q4KHV1yKt1B/WT1tAraUwQRNYwrSeJb
xpNf1Z5EE1JFbS3lZVe2iE7sAgVVbtRBRJ/eZBUgh90WjWFMbYsiBtOBFOtYXofTUZjkq2PVq4Hh
Ll/4e7FTnIA5avoYh1OOAbG96+ACp9csMU7PzWTOX1BypF2a069x7V/RfZSQKdBl3YpcKZb1HKHW
WHzgO0MgaMqQ34K4Tzt5cm2BVnIv0qJxgUj/llx6EB5XVxJQ5Sxiueb0Oo2KJrPNtJbS7x2EKoh3
jncsiqXTKHZgsQf9TldOi4BltssFrSdRtNp63hbZ6N2S5qACAIkIG4M8qJT4c4Nd7UIP7pA0pCeZ
aFzQXtc1SlPZb03AEmJvSDpUKLmzpwVyVF6lRBgQ//cPOFlu2ZuC9NUcTrnkj0y8tAudP9qgF5dm
xUFg/DmpKrFME3+WRRJ+DZzXd1PrmqKA3mFUWLbGsPmaCp9swZh31gPF7n1n0VE+IYFX6lm9JUoY
YEsjfoAokf0/82eEKVcCDHdaOBvwyp25XElkLlyuykVRXrR2qGMZa/Is+KRCy2SP1O33/x1ZXvJe
DMCaIG1e0b9wMsMoADJQ2glnBAWlCgcVOVw+8Qr9TVcZ0dY2e5w176QUD35apTHCfRfA+gV89pQQ
3xbewc48zDMK/2nC9PnBwkurEG3M0OAGiJdFJIBeL4MmyuSGzKqmN2sSLF+oUbuioU3nnfzVoxiX
y5D5ydd2ugwloBjiFeE0+8bgeANWKUIuCEoa3cmqDmtNDdYAQrGJnlJogpOym7/hjeqFZLOKYoUw
DBEebEMoidK6b5wBFNJtqMmFHvGjS/35XVt8Brg5welu2cDIF29NRAzMva9Lrijr8QgSkD6I8e7z
pci/HRfKHEmjFdcIwDr6U6KWo6GpiaMxfXUyCvSeGRJxKQHYI4B47RHQV+DUfWUU/SIb5R1GiW69
pFjg/xVQdsdpM9hN9PS2Yy9tjKQSrANhOVYPqYY9PsXN0kaLiiSbLBpOt1M3u0jVICEzPwPxl0BM
u+Q4TIXMRTwnjSCWETVEMt1GWYJGoCFcphOVjlmdlYcZ4zMTlNe/n3B0+G29QRL6yvtB49pBMAD+
ZojYBbajiB+8YEmXukEDrywBa/7aLd22ImuUj0UJCpQ0LGKkBk07Aov4SpOAx+Kw9aD8kUhsKLAK
pymFSKtLmfi+LQ6f7sIQs+kd+BYlz/3vjtpusUpixQ8PoNytD3Mhk9MzxSElAtImAN89Lz6cHXZ+
9GhSPnozp1O0v2tTKHejGcW2N1/EYpr6HObn0NGiSxv00O4FUl2T3XVrWoI8aeTqXmvRdBv9WXrt
WHC/VUN2GhKiCuMzUUf6Te26hUVgn2SR7/HCuzVniISIfANvLtEpUV7dnJ+owOZCn7l5+wcSWwro
11xh/KYj1xeMqfMu4mZqThVUZM+g5yx0U3QsZIJatzSvS+bVoouNxkxRVRU9xDpMwrVfF0hCikTZ
uQSSVkrwHuZbP5fY6f488NKSfsTKwWq/9roJ6uAc2coqLcfKR+R3tv7AOFbe2Mdzz/2BksSffqsP
7JMSzUKwN1LWZeCwjSNEVtFrAiIXEyq5+gxt3uGU6MwLhRnMoMmKtEtsFqC/ueZoLpGYfd7lpa9I
7d7+/23DXHMaQJNnxuVyx6QQSgmqzdOqE5fNjc+y1wnmnn3SDkraBh6DphqPlh3I/keKkrg6mhmC
YxS6GatCqlH4zKM/4KlfG7ArfbDhmTAeUgv7dP6IRUEiUJ68nYCXepm6boosUU3APKr99efk08uO
W6ofpPPUnLW4/JcxK9ZDcItBJrwr1bz2nWVf32l6MOhFBfi3QZAC+Wmg8pRaHOa78XI6MTYF6AfK
1nmNDckG7TDujbunUNGVD0qpVoQFWVw5bhdwmwBa4IdsuS/2tgxRHtwzUGaN/qs3NI88sB+nCNGe
jUeDH1rab0FpTNvEiL3hiwdsMabjskJaz0jNRube2GnU+4d37lX7qIJ4KkV/27RyfVp4QQ6Tw2bU
plqBW4iX3f4KQ/agFh3R2igQh8rDZU82jl5igOLRKPhfPb294H391WJddUcj6Y1ODSqQSvIfGyDw
af2Lm9cDDdIVONGuXpuiaWfTV8H4gUZpDu2T9OKWOUBCyfTc2h2oXg+m8nXtvFpQUNK23PUGLo9B
SX71biFwWhZK2y2VoC7RN1DwP07MIxocpFmCQ5OOsfgHIVMAAy7kJ6jP3Um+8gBrXittTPojAlak
isSLR6eB1JAJYDMlG6xALXsAdooEJCWlWzSE1BajFx+iFrKZ7s6ZgdK6Xucgot8oXE2JhDZW9iUs
7M5etUlBZeTSSTocuUJEuzA9u4tmX9n34MbA8pDPSRQPvba/DGnhqFKZe2ayj2JXEfFgGNaYjMqy
ONn7tlI1XKSWug8OFyQRf/griLIHWakJyd85jHuJAvbOL/a85CiVZAVMSCHJaaR+bXcm0H5B+Yrf
/vmQDd+qaWAWAaOsxYf2AF+YIfYiiNz5IyUFJYp77ZRt1Eu9DgypoKtieIQ2QvirinLtbIUi8MV/
c/6znn+Mm7nLWHWKOcW/6gVcbuaemUBKviM/1nD4tUDG8pbHzRLXWELmcTtnHaDheHJvDigf7GWC
8Sniv+fS9dXSqfMUxwn8oPUa0aBIFAAtDAlIbY6WjxzZJ+oMvSCn1fWm/FPfnCsr9t6LumQTD9kI
6XpSD6z7BOV+3+ItTzFAVDf9gXEvFB2v6K0gvzJMyvPZnPJmiBuv1TtoqLROgFl0Ou32l9Dp+u7o
gNZolS+2z2SvnQ8j+oUCf4Rp8PmjUSFOI0/p+XRx39R2WfFwJLJ8sAw9Bi6dZb4D2OvFEMm1JcTf
KgPkDRFEzCORnWLdsY5IyPgQqM0H76rEokQ+ynR8DDCe5QHylko5OglPvQ26JTIeWh0FOaJQWVDN
DSe+JoAASk/4cxlYqpuDKgbM637qggfvhFGbH78+6igZC5/lGwLScqL1sMgyi7En00KToNxlIeCV
aCgeVoIMH8nIESjmZxY/YP3VkT9imz6oyVoU+xxAv0nlNTLIeQEhzVrzGaVDKlh8inFcOu+/lOkA
UoP7V3rxcke0aQBnyP4h7oE8+ghiDXHmBy7I6+Z873+8fLFd1735EOyMoHBda8fFBs4duaIjMXd3
5AM4MJXLrNz/s5ElMXYyxYj+KwP57H7iLkpP/IVHv1o0fliydLN69G46UDciCIe1eN4T7PDeAEgS
jYdnj4xF8Ld/CUss1E1ltaCK1icyAvTTZfDEiq5KJWHPENlYTEi7IqUIxgITAyTg9IoVZXvNbxwr
N5qAi5Rkk7xkvQlF2lLRyGoFuCYmjKOLZKVHZS4RrOC53tnMkSGa8Jd+Hi6zprp0fVMpRLQS9NXs
KhVsPdzpZQoaY4pPR176l2e8+OXMmEJ7/78eZtZS9fKks3Af7Q3777PYSqhpr1SYz2Z5kFO3gtpu
1P/CUGoUr7T8KJk4VF5lmsUzVE5mJz3utNRsNtmyzR1FOAbky9/G35sC2Ku13fsf43gRGSg2fxBI
iQS4sPPauB0AIH7jcfsO1iVQSWgnSlbfmW5cYJ/zxMHos30Ya35v6OH7qpR4W91dHGBXUjM47bvq
RItxGgbcZC+/tKvwhrOS8oUHb2abCczeGrirBMwRc+cson5P/2BRfGbEmpevvr8N1Epg40RGgyNH
LrO3OqOI8YM8ry6+pdF8atXhXvShMmcIyLksZ3KtgtWxYIJyOQMKcNYj34lfT8pFf6UTGLR72Axf
U0ytVVigGT0e1j7CipoHzJTCHp3/vIh2N+rmaStkBoExG+ki88m+yPVbXcO0iPjzmTDBo1QOC/ZA
bsoBYlebrRowDLAHdDhRbL62ncvv6qUAWP0TEId5xhg66/+nx4pELkW0jAVFw0OA62kRDeJLBb7+
G4Vq2Kxciqb4eSuPDQmB1C3GgCJ2knFPsgGsCcl1TJchrhpDVMMOc5YnzgaNfTY6vxNYFBrdR009
OK4Zi4qFT9iWQEeXWXFBCf7sEYgMrX9RHYJ8PFv0aNzKBbNbJdMvkFjxTZgIzOMuXV7Tx49hDfgJ
OINUBzPskGs4r1cXCoG195X+rEV3641LdV3QGSUKIx6PMMrksKtKspZxXW7qeMJh8oEDt7aMnRqB
IxOR3EBxnCD7abLEOC08ysVPJhzIkhparkgmGFO7lbZ8BqjryIJTADVA3GuxfLIe5Gc8etWye3yv
5aI/vjamaseMkVUTWPkkLokPTEXhDEGkxSQNNJCo/HQqs9WZQARH4nzxsdBfRKY5PuKyvMC19UwL
xW9KV/5ROkELdd9f5+sZQIUp4l99x00Kmf+4RUxdZ5FA/vkA4JYYN93mw028xlVCv2lvgRJ1ov9z
bGyeN7KAKjYGoUCR/lTicr5K4eLWgfNoni012mLjGgFcknJP84SoNBKPIKRxY2CfXffrmHKGMfkv
duYWiFmVanmGjPQzoviPLOpFZxluD8p9Zc3yZt0R8XcYNJwjRt1ThacKbcOTjsYeBc50KNWFRNDF
d9pQ+nh2UoARV7bCOfIFvTa9vBxC2yANku4PS4NPFNw45+9KYzyGzuM79RBHj0XOuoMQ6uQSXMkD
KAnDEp7lH1i/SiiTD6NujyawmJxV7RC2/V1QCG9Xdj5702ZF5cGzzoyP1GZuY6hDMCQAzfP8yQ93
ib0qreYZATy7826x9lR6q17ztbUh4hlipUTJQcKSyB+3Z5Iijr/pI1ylrRtKmUtAM6IPzm/nZD6r
3bGASqaFGc+TtzbtmpZpizFe4ljM7nqnb9qjJfNl/50hJNpBcI4PJNMPxfZ/YONY6AC1ruxSOHVj
MXYAA0zvWl+mxi+gwhrkelveNYHhYGvtHnMlcYrP2Vkjvagq/57NoeHRnJssRhMwZHoqAC7xP7y5
jVKnXcQECahIWmfasfUBt7QR8ts5CvNdPTaVb/4hDiNck9dcQjmJgpmBRkeL2U/IZMOf9rEIIB4x
U56eBq6Sd910hqs/FTiqmIdgojCYJDuc8N2k2ixsOy1NvpgnZdT/wai1PQJbHtspDxWO3HgiF1xQ
+wFVNU/6Dx3X3IPMb7LezWc7t4x7Emw307HFI7VUmz2aOxu1VVmNc5nxCSLU2aUNhM/BUse/ylWr
8QSs0+zWBL2CBQVblKGt8QOo7ZeiEP/j9282BpsXI9H7yTmBXdULMQjQl1tCNKu6Q4rBGk+MtD4p
Ld8S1ca2PKiIc1dXWAzNlCDzwEC/j+RWc83vqANQIDvSa1427bKkiMi3zINrOtX8WpxWlttv3ZRX
25y5XsxN5GtIj1xNs4SYUtFkviF4lYXIweEZyfhkgmrVS0fSBBW0I78TT4C4QMqtq2HBdXmSW9x+
kScAS338h9OUld2W1eA93zo/r4T1CPtFHcA65nv6OcJGyw2CK/VsAnldOtbbEFDuYGSyrQXRKtGS
6vNrdQe4UVWtU7+kkRKS1Mmwq7+aR/f36cbfkZMAQ6tGnbF8j0UcLx9JEO1qrf6CNW6BOMRMiaOE
ZRkfnLxp/AVwIL+bvmg2Q50uWx6JNKn0dw/i8pUBAJva9mM9Fdoonhi0nsGc8eBxHuDwPNOiTmWE
kDcyCahrtfXPLNo98xqQ68dGksx1PXW+bBOKgjhmULeoMRJZdvHpgbZMUh3dYTgGws9G+QRBaR3O
C4PLhqzbHsqPLZbBz0B3a6cPA6I69i2uh4LG6b9YkShfdTrPl8aL0ic2628tacjGQUADKqLW56Jq
JtNGZaAPRELgm9qLbKkQzJ6dYkwUFGzXCITFZZixvZdgOzjx7oAhXiUkMWor4Nnj1RefbA8NI5bh
jGFNJXFO43ikHpnnNSOazL3mIDGdW1UptAbY1f98PcM9se8Hc12E1c2npFlw7qI2hvSWbkdUyTrS
uqau8je0O97f4AuSaJk21Ze2Mxy/2unqxppdepjvdfJUcyDaYA1kkeXMbs0aM3V3XZwL24YpMuRK
NquWDHhj+wyBwHPhkaNGpH5b4DJZCaM/rFrXzK7Cfq1QgLrFp5jcJU+f0l3d3DwLY+ZmO/O3eUkr
Xt3MKFNvbRzh/mOa7hLptKjhCt1yKx129zel+xRoxiTrhXZd5U7KYs+5tpmlJFd6hLZ7XmBJnJYi
6Mqg8Jm5WDuouX2sWO7AJGzrUmqTe6srtjYplnicmwu3H88rxrwFEbpfEJtWxanviobLDP0Y1xxl
8vX2Kh5gbVAVnzr+pxIwKI7A+EY3AFjDYVhoI5UuxI4xXBfItkZOSH4BPUM3UfiLDPm0jg0eVlRj
0hrT1AXF+Nep9bqyVXSnerWqVxCQ8yBETrU5xsUIYKbvlJE2RRQKNtLtoUOobPpsTcReIvtZjpjM
aYjYzxzToe4vGlme162srzvNRZumNnOOJ7M5oe+KU4hGVfFUsUfkGKycGZsIDBO528SMXtAvEL/7
BMuPOISdRLb7VcmuRo99rqFHQ3Whu90XMro3+7ODI9jYSZ7vIcbCQrmcyvuEyOrm4hi1vo/ateJd
Gg7nxD2Xu5ybSSOuM5Om/xu86JzDD0ij0QZOSXJQHSJW2L7aPrM7Fc0uEKGt9pqmlTouxjFX5lRZ
3Qd6vPirF5iKliYaw92NRkueTkos4KSx/Nglk+NkPs074wpy6P/uR7L8zKOmlsK3z/2u50j+JZR3
StbXok03+j0PSW2IVS8IN5lq94FLfTok80LmOHBHVaougLUje6LH94V9W9z1lUZacfy96mg8xctL
d2tvQ8MMhwnDV4irDyY9qjk6kK3b005cT5JZwYrcPHTn5gJt/JREJjeCbsV5K/fx/UpH2F/gtHUy
fSRH/WALJatzlYPl+pukEaf/4gL6XTLXgv4zoGb/p6MpNDVkGvMSf9dszWVvkrg5ZsjmB5kF/ETA
IoXY8jmDS5UvoLpQbDJqmd4Ntw6J3bnF3P/O+3oUsKFYLKJdb4i8csrsaEAvsg3T3wDt6aQej25j
T9VxljP4nd0BFI/FpUPevz8KHkYQ/+LuJWFH+z1y7O7xbIObJBJuE0XJFvLjCl/3hjJIqhMc15U3
JyyQKFVnhLSGclWsEMru6Hjzixpl4hWYkA2uXwq7DDl0yFrpak4zpK7BMaiJXLOaRJiLGUrF41XF
19AKXsUgliIozSIEMZDVNd0AlFNREzz8wzp/kOFrzHS75briWolulXQYu02FiHX5jRvsOzEp9uLA
rdpRScnY6pFnWk3rsfNAEehBcXyOJHEud9b+A8Un49cP9Tf8Qq6nteLuFVA37o0nFjtwb44EuzkL
yBQVxiGMKqL4gG6Q4LGceu91ydcKQChiuxO+iBx/w25MAzL94zKznZCOTBrvH4BOr1mIX1keVGuS
g75l2h4nCbZQtWBEys8jZKbhN6eckd1dX6Wuwp6FlCpcH00tALqCYY+QYc/6RMBEsLMjZW3oVBc2
XywpJp1HT+X2qxFwlSWMGbc9mD2Rt3j8kDxrkNEcGpCvTmLEE4uJYeFAwc5hqAJTpmyByUN1ZTGI
B/16RDVI1pHtcpHteLd3nQ4POvP874yO0sx1OIZvEyRAXE4kP0Z+BcBG/XsqnRvPhzapzMRl67qE
TmP68wpaeYDPI+Q3sW5yTQiCY2xR1SL3dwxgFA8R+rtB8rZB/BsyJPyYU+vZYVlh/XqcxNhdFJCz
/RYNiNcqrpv25sJkEgOKn08+uFZNG+Y09+69rqwQa/+OXkZr1E5xcz9vDuyMViorte0MB6WsLQxk
lGJX0FIukpK9z+XdBQamJT1/n9026ALQC2WMXAby7Uy1cxZ2wCtLxlgzcwx/Y77JGp8FN7Z2w0GK
gz7JQLeRMzQT9NAZsg3efDA3cHDcVvJe7pKiNLOeaNYQ/gJuD1SMFWcQKjSz0O5n6kKExOXRjHqu
GSt+Af97Q2YnQwhyk3imBcF8r4QWiIPmJAC3WnIVNbXPJ5CsSRtLb35XfrADtsefmfE/CAxGfwjQ
SHCUXkt9VKsoUa1Oes80zFKhjbKn2Yl3OtJpynXRkC37L51w4ZvjWr/rT2DewBQ5D47z7QRhmFiO
9z4dI8o0Wgua0eFrYrZS0pb8BjYyDmGxPcY5Btr68hrRdkbR3Qplp8koNFus6smDRd54wRGjD/CK
AkpEqPJAuRGjpYX0qJj92UpVTZw9rUQ7m1cG/thDWyq63eDOp7wUfa6gTsTm7IUzgghc/tk3nZTO
3iFD6HrYcW4+AjxzPsv7n8u+YIhxegS9lg+3fa0uGhXZsJLXNQ2gDIISFPDpI0f9J57OLDYCnVd3
Q0kFmruge6v1woL2vH6JHh2bWCfYd5V7OBxqeXFQbqBq0H6azmF9WHKzn1f3nJPmF1uslOyEtV5x
N7z8p0Yq79z5b0akagQL84+0rCeWmAp91ra/4/v0OxraBvbq6c/y6DDcqvPgAdz2NA27A9jERCJL
J4sT7kHfpbz6eXDyetwndyMfI6XmfKw3tUZDE3nXP/SJNVHO7kRvGxBq0dhCY+EK2WvHiVLOJTeS
mzSm5cu3JHXSUuuVIz+h0UM+Dd9tD1j1oIPS02tqzJM6IyksNckLolvABC2v9qIUZWisvHA2CJiW
l1Ap1w+USHGR+9XM9r4JFYN8QQ==
`pragma protect end_protected
