          "REG_HIGH_ID0_P01"      : u_nps_reg.REG_HIGH_ID0_P01  = value;
          "REG_HIGH_ID0_P23"      : u_nps_reg.REG_HIGH_ID0_P23  = value;
          "REG_HIGH_ID1_P01"      : u_nps_reg.REG_HIGH_ID1_P01  = value;
          "REG_HIGH_ID1_P23"      : u_nps_reg.REG_HIGH_ID1_P23  = value;
          "REG_HIGH_ID2_P01"      : u_nps_reg.REG_HIGH_ID2_P01  = value;
          "REG_HIGH_ID2_P23"      : u_nps_reg.REG_HIGH_ID2_P23  = value;
          "REG_HIGH_ID3_P01"      : u_nps_reg.REG_HIGH_ID3_P01  = value;
          "REG_HIGH_ID3_P23"      : u_nps_reg.REG_HIGH_ID3_P23  = value;
          "REG_HIGH_ID4_P01"      : u_nps_reg.REG_HIGH_ID4_P01  = value;
          "REG_HIGH_ID4_P23"      : u_nps_reg.REG_HIGH_ID4_P23  = value;
          "REG_HIGH_ID5_P01"      : u_nps_reg.REG_HIGH_ID5_P01  = value;
          "REG_HIGH_ID5_P23"      : u_nps_reg.REG_HIGH_ID5_P23  = value;
          "REG_HIGH_ID6_P01"      : u_nps_reg.REG_HIGH_ID6_P01  = value;
          "REG_HIGH_ID6_P23"      : u_nps_reg.REG_HIGH_ID6_P23  = value;
          "REG_HIGH_ID7_P01"      : u_nps_reg.REG_HIGH_ID7_P01  = value;
          "REG_HIGH_ID7_P23"      : u_nps_reg.REG_HIGH_ID7_P23  = value;
          "REG_HIGH_ID8_P01"      : u_nps_reg.REG_HIGH_ID8_P01  = value;
          "REG_HIGH_ID8_P23"      : u_nps_reg.REG_HIGH_ID8_P23  = value;
          "REG_HIGH_ID9_P01"      : u_nps_reg.REG_HIGH_ID9_P01  = value;
          "REG_HIGH_ID9_P23"      : u_nps_reg.REG_HIGH_ID9_P23  = value;
          "REG_HIGH_ID10_P01"     : u_nps_reg.REG_HIGH_ID10_P01 = value;
          "REG_HIGH_ID10_P23"     : u_nps_reg.REG_HIGH_ID10_P23 = value;
          "REG_HIGH_ID11_P01"     : u_nps_reg.REG_HIGH_ID11_P01 = value;
          "REG_HIGH_ID11_P23"     : u_nps_reg.REG_HIGH_ID11_P23 = value;
          "REG_HIGH_ID12_P01"     : u_nps_reg.REG_HIGH_ID12_P01 = value;
          "REG_HIGH_ID12_P23"     : u_nps_reg.REG_HIGH_ID12_P23 = value;
          "REG_HIGH_ID13_P01"     : u_nps_reg.REG_HIGH_ID13_P01 = value;
          "REG_HIGH_ID13_P23"     : u_nps_reg.REG_HIGH_ID13_P23 = value;
          "REG_HIGH_ID14_P01"     : u_nps_reg.REG_HIGH_ID14_P01 = value;
          "REG_HIGH_ID14_P23"     : u_nps_reg.REG_HIGH_ID14_P23 = value;
          "REG_HIGH_ID15_P01"     : u_nps_reg.REG_HIGH_ID15_P01 = value;
          "REG_HIGH_ID15_P23"     : u_nps_reg.REG_HIGH_ID15_P23 = value;
          "REG_HIGH_ID16_P01"     : u_nps_reg.REG_HIGH_ID16_P01 = value;
          "REG_HIGH_ID16_P23"     : u_nps_reg.REG_HIGH_ID16_P23 = value;
          "REG_HIGH_ID17_P01"     : u_nps_reg.REG_HIGH_ID17_P01 = value;
          "REG_HIGH_ID17_P23"     : u_nps_reg.REG_HIGH_ID17_P23 = value;
          "REG_HIGH_ID18_P01"     : u_nps_reg.REG_HIGH_ID18_P01 = value;
          "REG_HIGH_ID18_P23"     : u_nps_reg.REG_HIGH_ID18_P23 = value;
          "REG_HIGH_ID19_P01"     : u_nps_reg.REG_HIGH_ID19_P01 = value;
          "REG_HIGH_ID19_P23"     : u_nps_reg.REG_HIGH_ID19_P23 = value;
          "REG_HIGH_ID20_P01"     : u_nps_reg.REG_HIGH_ID20_P01 = value;
          "REG_HIGH_ID20_P23"     : u_nps_reg.REG_HIGH_ID20_P23 = value;
          "REG_HIGH_ID21_P01"     : u_nps_reg.REG_HIGH_ID21_P01 = value;
          "REG_HIGH_ID21_P23"     : u_nps_reg.REG_HIGH_ID21_P23 = value;
          "REG_HIGH_ID22_P01"     : u_nps_reg.REG_HIGH_ID22_P01 = value;
          "REG_HIGH_ID22_P23"     : u_nps_reg.REG_HIGH_ID22_P23 = value;
          "REG_HIGH_ID23_P01"     : u_nps_reg.REG_HIGH_ID23_P01 = value;
          "REG_HIGH_ID23_P23"     : u_nps_reg.REG_HIGH_ID23_P23 = value;
          "REG_HIGH_ID24_P01"     : u_nps_reg.REG_HIGH_ID24_P01 = value;
          "REG_HIGH_ID24_P23"     : u_nps_reg.REG_HIGH_ID24_P23 = value;
          "REG_HIGH_ID25_P01"     : u_nps_reg.REG_HIGH_ID25_P01 = value;
          "REG_HIGH_ID25_P23"     : u_nps_reg.REG_HIGH_ID25_P23 = value;
          "REG_HIGH_ID26_P01"     : u_nps_reg.REG_HIGH_ID26_P01 = value;
          "REG_HIGH_ID26_P23"     : u_nps_reg.REG_HIGH_ID26_P23 = value;
          "REG_HIGH_ID27_P01"     : u_nps_reg.REG_HIGH_ID27_P01 = value;
          "REG_HIGH_ID27_P23"     : u_nps_reg.REG_HIGH_ID27_P23 = value;
          "REG_HIGH_ID28_P01"     : u_nps_reg.REG_HIGH_ID28_P01 = value;
          "REG_HIGH_ID28_P23"     : u_nps_reg.REG_HIGH_ID28_P23 = value;
          "REG_HIGH_ID29_P01"     : u_nps_reg.REG_HIGH_ID29_P01 = value;
          "REG_HIGH_ID29_P23"     : u_nps_reg.REG_HIGH_ID29_P23 = value;
          "REG_HIGH_ID30_P01"     : u_nps_reg.REG_HIGH_ID30_P01 = value;
          "REG_HIGH_ID30_P23"     : u_nps_reg.REG_HIGH_ID30_P23 = value;
          "REG_HIGH_ID31_P01"     : u_nps_reg.REG_HIGH_ID31_P01 = value;
          "REG_HIGH_ID31_P23"     : u_nps_reg.REG_HIGH_ID31_P23 = value;
          "REG_HIGH_ID32_P01"     : u_nps_reg.REG_HIGH_ID32_P01 = value;
          "REG_HIGH_ID32_P23"     : u_nps_reg.REG_HIGH_ID32_P23 = value;
          "REG_HIGH_ID33_P01"     : u_nps_reg.REG_HIGH_ID33_P01 = value;
          "REG_HIGH_ID33_P23"     : u_nps_reg.REG_HIGH_ID33_P23 = value;
          "REG_HIGH_ID34_P01"     : u_nps_reg.REG_HIGH_ID34_P01 = value;
          "REG_HIGH_ID34_P23"     : u_nps_reg.REG_HIGH_ID34_P23 = value;
          "REG_HIGH_ID35_P01"     : u_nps_reg.REG_HIGH_ID35_P01 = value;
          "REG_HIGH_ID35_P23"     : u_nps_reg.REG_HIGH_ID35_P23 = value;
          "REG_HIGH_ID36_P01"     : u_nps_reg.REG_HIGH_ID36_P01 = value;
          "REG_HIGH_ID36_P23"     : u_nps_reg.REG_HIGH_ID36_P23 = value;
          "REG_HIGH_ID37_P01"     : u_nps_reg.REG_HIGH_ID37_P01 = value;
          "REG_HIGH_ID37_P23"     : u_nps_reg.REG_HIGH_ID37_P23 = value;
          "REG_HIGH_ID38_P01"     : u_nps_reg.REG_HIGH_ID38_P01 = value;
          "REG_HIGH_ID38_P23"     : u_nps_reg.REG_HIGH_ID38_P23 = value;
          "REG_HIGH_ID39_P01"     : u_nps_reg.REG_HIGH_ID39_P01 = value;
          "REG_HIGH_ID39_P23"     : u_nps_reg.REG_HIGH_ID39_P23 = value;
          "REG_HIGH_ID40_P01"     : u_nps_reg.REG_HIGH_ID40_P01 = value;
          "REG_HIGH_ID40_P23"     : u_nps_reg.REG_HIGH_ID40_P23 = value;
          "REG_HIGH_ID41_P01"     : u_nps_reg.REG_HIGH_ID41_P01 = value;
          "REG_HIGH_ID41_P23"     : u_nps_reg.REG_HIGH_ID41_P23 = value;
          "REG_HIGH_ID42_P01"     : u_nps_reg.REG_HIGH_ID42_P01 = value;
          "REG_HIGH_ID42_P23"     : u_nps_reg.REG_HIGH_ID42_P23 = value;
          "REG_HIGH_ID43_P01"     : u_nps_reg.REG_HIGH_ID43_P01 = value;
          "REG_HIGH_ID43_P23"     : u_nps_reg.REG_HIGH_ID43_P23 = value;
          "REG_HIGH_ID44_P01"     : u_nps_reg.REG_HIGH_ID44_P01 = value;
          "REG_HIGH_ID44_P23"     : u_nps_reg.REG_HIGH_ID44_P23 = value;
          "REG_HIGH_ID45_P01"     : u_nps_reg.REG_HIGH_ID45_P01 = value;
          "REG_HIGH_ID45_P23"     : u_nps_reg.REG_HIGH_ID45_P23 = value;
          "REG_HIGH_ID46_P01"     : u_nps_reg.REG_HIGH_ID46_P01 = value;
          "REG_HIGH_ID46_P23"     : u_nps_reg.REG_HIGH_ID46_P23 = value;
          "REG_HIGH_ID47_P01"     : u_nps_reg.REG_HIGH_ID47_P01 = value;
          "REG_HIGH_ID47_P23"     : u_nps_reg.REG_HIGH_ID47_P23 = value;
          "REG_HIGH_ID48_P01"     : u_nps_reg.REG_HIGH_ID48_P01 = value;
          "REG_HIGH_ID48_P23"     : u_nps_reg.REG_HIGH_ID48_P23 = value;
          "REG_HIGH_ID49_P01"     : u_nps_reg.REG_HIGH_ID49_P01 = value;
          "REG_HIGH_ID49_P23"     : u_nps_reg.REG_HIGH_ID49_P23 = value;
          "REG_HIGH_ID50_P01"     : u_nps_reg.REG_HIGH_ID50_P01 = value;
          "REG_HIGH_ID50_P23"     : u_nps_reg.REG_HIGH_ID50_P23 = value;
          "REG_HIGH_ID51_P01"     : u_nps_reg.REG_HIGH_ID51_P01 = value;
          "REG_HIGH_ID51_P23"     : u_nps_reg.REG_HIGH_ID51_P23 = value;
          "REG_HIGH_ID52_P01"     : u_nps_reg.REG_HIGH_ID52_P01 = value;
          "REG_HIGH_ID52_P23"     : u_nps_reg.REG_HIGH_ID52_P23 = value;
          "REG_HIGH_ID53_P01"     : u_nps_reg.REG_HIGH_ID53_P01 = value;
          "REG_HIGH_ID53_P23"     : u_nps_reg.REG_HIGH_ID53_P23 = value;
          "REG_HIGH_ID54_P01"     : u_nps_reg.REG_HIGH_ID54_P01 = value;
          "REG_HIGH_ID54_P23"     : u_nps_reg.REG_HIGH_ID54_P23 = value;
          "REG_HIGH_ID55_P01"     : u_nps_reg.REG_HIGH_ID55_P01 = value;
          "REG_HIGH_ID55_P23"     : u_nps_reg.REG_HIGH_ID55_P23 = value;
          "REG_HIGH_ID56_P01"     : u_nps_reg.REG_HIGH_ID56_P01 = value;
          "REG_HIGH_ID56_P23"     : u_nps_reg.REG_HIGH_ID56_P23 = value;
          "REG_HIGH_ID57_P01"     : u_nps_reg.REG_HIGH_ID57_P01 = value;
          "REG_HIGH_ID57_P23"     : u_nps_reg.REG_HIGH_ID57_P23 = value;
          "REG_HIGH_ID58_P01"     : u_nps_reg.REG_HIGH_ID58_P01 = value;
          "REG_HIGH_ID58_P23"     : u_nps_reg.REG_HIGH_ID58_P23 = value;
          "REG_HIGH_ID59_P01"     : u_nps_reg.REG_HIGH_ID59_P01 = value;
          "REG_HIGH_ID59_P23"     : u_nps_reg.REG_HIGH_ID59_P23 = value;
          "REG_HIGH_ID60_P01"     : u_nps_reg.REG_HIGH_ID60_P01 = value;
          "REG_HIGH_ID60_P23"     : u_nps_reg.REG_HIGH_ID60_P23 = value;
          "REG_HIGH_ID61_P01"     : u_nps_reg.REG_HIGH_ID61_P01 = value;
          "REG_HIGH_ID61_P23"     : u_nps_reg.REG_HIGH_ID61_P23 = value;
          "REG_HIGH_ID62_P01"     : u_nps_reg.REG_HIGH_ID62_P01 = value;
          "REG_HIGH_ID62_P23"     : u_nps_reg.REG_HIGH_ID62_P23 = value;
          "REG_HIGH_ID63_P01"     : u_nps_reg.REG_HIGH_ID63_P01 = value;
          "REG_HIGH_ID63_P23"     : u_nps_reg.REG_HIGH_ID63_P23 = value;
          "REG_ID"            : u_nps_reg.REG_ID        = value;
          "REG_LOW_ID0_P01"       : u_nps_reg.REG_LOW_ID0_P01   = value;
          "REG_LOW_ID0_P23"       : u_nps_reg.REG_LOW_ID0_P23   = value;
          "REG_LOW_ID1_P01"       : u_nps_reg.REG_LOW_ID1_P01   = value;
          "REG_LOW_ID1_P23"       : u_nps_reg.REG_LOW_ID1_P23   = value;
          "REG_LOW_ID2_P01"       : u_nps_reg.REG_LOW_ID2_P01   = value;
          "REG_LOW_ID2_P23"       : u_nps_reg.REG_LOW_ID2_P23   = value;
          "REG_LOW_ID3_P01"       : u_nps_reg.REG_LOW_ID3_P01   = value;
          "REG_LOW_ID3_P23"       : u_nps_reg.REG_LOW_ID3_P23   = value;
          "REG_LOW_ID4_P01"       : u_nps_reg.REG_LOW_ID4_P01   = value;
          "REG_LOW_ID4_P23"       : u_nps_reg.REG_LOW_ID4_P23   = value;
          "REG_LOW_ID5_P01"       : u_nps_reg.REG_LOW_ID5_P01   = value;
          "REG_LOW_ID5_P23"       : u_nps_reg.REG_LOW_ID5_P23   = value;
          "REG_LOW_ID6_P01"       : u_nps_reg.REG_LOW_ID6_P01   = value;
          "REG_LOW_ID6_P23"       : u_nps_reg.REG_LOW_ID6_P23   = value;
          "REG_LOW_ID7_P01"       : u_nps_reg.REG_LOW_ID7_P01   = value;
          "REG_LOW_ID7_P23"       : u_nps_reg.REG_LOW_ID7_P23   = value;
          "REG_LOW_ID8_P01"       : u_nps_reg.REG_LOW_ID8_P01   = value;
          "REG_LOW_ID8_P23"       : u_nps_reg.REG_LOW_ID8_P23   = value;
          "REG_LOW_ID9_P01"       : u_nps_reg.REG_LOW_ID9_P01   = value;
          "REG_LOW_ID9_P23"       : u_nps_reg.REG_LOW_ID9_P23   = value;
          "REG_LOW_ID10_P01"      : u_nps_reg.REG_LOW_ID10_P01  = value;
          "REG_LOW_ID10_P23"      : u_nps_reg.REG_LOW_ID10_P23  = value;
          "REG_LOW_ID11_P01"      : u_nps_reg.REG_LOW_ID11_P01  = value;
          "REG_LOW_ID11_P23"      : u_nps_reg.REG_LOW_ID11_P23  = value;
          "REG_LOW_ID12_P01"      : u_nps_reg.REG_LOW_ID12_P01  = value;
          "REG_LOW_ID12_P23"      : u_nps_reg.REG_LOW_ID12_P23  = value;
          "REG_LOW_ID13_P01"      : u_nps_reg.REG_LOW_ID13_P01  = value;
          "REG_LOW_ID13_P23"      : u_nps_reg.REG_LOW_ID13_P23  = value;
          "REG_LOW_ID14_P01"      : u_nps_reg.REG_LOW_ID14_P01  = value;
          "REG_LOW_ID14_P23"      : u_nps_reg.REG_LOW_ID14_P23  = value;
          "REG_LOW_ID15_P01"      : u_nps_reg.REG_LOW_ID15_P01  = value;
          "REG_LOW_ID15_P23"      : u_nps_reg.REG_LOW_ID15_P23  = value;
          "REG_MID_ID0_P01"       : u_nps_reg.REG_MID_ID0_P01   = value;
          "REG_MID_ID0_P23"       : u_nps_reg.REG_MID_ID0_P23   = value;
          "REG_MID_ID1_P01"       : u_nps_reg.REG_MID_ID1_P01   = value;
          "REG_MID_ID1_P23"       : u_nps_reg.REG_MID_ID1_P23   = value;
          "REG_MID_ID2_P01"       : u_nps_reg.REG_MID_ID2_P01   = value;
          "REG_MID_ID2_P23"       : u_nps_reg.REG_MID_ID2_P23   = value;
          "REG_MID_ID3_P01"       : u_nps_reg.REG_MID_ID3_P01   = value;
          "REG_MID_ID3_P23"       : u_nps_reg.REG_MID_ID3_P23   = value;
          "REG_NOC_CTL"       : u_nps_reg.REG_NOC_CTL       = value;
          "REG_P00_P1_0_VCA_TOKEN"        : u_nps_reg.REG_P00_P1_0_VCA_TOKEN    = value;
          "REG_P00_P1_1_VCA_TOKEN"        : u_nps_reg.REG_P00_P1_1_VCA_TOKEN    = value;
          "REG_P01_P2_0_VCA_TOKEN"        : u_nps_reg.REG_P01_P2_0_VCA_TOKEN    = value;
          "REG_P01_P2_1_VCA_TOKEN"        : u_nps_reg.REG_P01_P2_1_VCA_TOKEN    = value;
          "REG_P02_P3_0_VCA_TOKEN"        : u_nps_reg.REG_P02_P3_0_VCA_TOKEN    = value;
          "REG_P02_P3_1_VCA_TOKEN"        : u_nps_reg.REG_P02_P3_1_VCA_TOKEN    = value;
          "REG_P10_P2_0_VCA_TOKEN"        : u_nps_reg.REG_P10_P2_0_VCA_TOKEN    = value;
          "REG_P10_P2_1_VCA_TOKEN"        : u_nps_reg.REG_P10_P2_1_VCA_TOKEN    = value;
          "REG_P11_P3_0_VCA_TOKEN"        : u_nps_reg.REG_P11_P3_0_VCA_TOKEN    = value;
          "REG_P11_P3_1_VCA_TOKEN"        : u_nps_reg.REG_P11_P3_1_VCA_TOKEN    = value;
          "REG_P12_P0_0_VCA_TOKEN"        : u_nps_reg.REG_P12_P0_0_VCA_TOKEN    = value;
          "REG_P12_P0_1_VCA_TOKEN"        : u_nps_reg.REG_P12_P0_1_VCA_TOKEN    = value;
          "REG_P20_P3_0_VCA_TOKEN"        : u_nps_reg.REG_P20_P3_0_VCA_TOKEN    = value;
          "REG_P20_P3_1_VCA_TOKEN"        : u_nps_reg.REG_P20_P3_1_VCA_TOKEN    = value;
          "REG_P21_P0_0_VCA_TOKEN"        : u_nps_reg.REG_P21_P0_0_VCA_TOKEN    = value;
          "REG_P21_P0_1_VCA_TOKEN"        : u_nps_reg.REG_P21_P0_1_VCA_TOKEN    = value;
          "REG_P22_P1_0_VCA_TOKEN"        : u_nps_reg.REG_P22_P1_0_VCA_TOKEN    = value;
          "REG_P22_P1_1_VCA_TOKEN"        : u_nps_reg.REG_P22_P1_1_VCA_TOKEN    = value;
          "REG_P30_P0_0_VCA_TOKEN"        : u_nps_reg.REG_P30_P0_0_VCA_TOKEN    = value;
          "REG_P30_P0_1_VCA_TOKEN"        : u_nps_reg.REG_P30_P0_1_VCA_TOKEN    = value;
          "REG_P31_P1_0_VCA_TOKEN"        : u_nps_reg.REG_P31_P1_0_VCA_TOKEN    = value;
          "REG_P31_P1_1_VCA_TOKEN"        : u_nps_reg.REG_P31_P1_1_VCA_TOKEN    = value;
          "REG_P32_P2_0_VCA_TOKEN"        : u_nps_reg.REG_P32_P2_0_VCA_TOKEN    = value;
          "REG_P32_P2_1_VCA_TOKEN"        : u_nps_reg.REG_P32_P2_1_VCA_TOKEN    = value;
          "REG_CLOCK_MUX"   : u_nps_reg.REG_CLOCK_MUX     = value;
