    .INIT_00(256'h022bfc205362f032022bfc2053801001022bfc250002d010022bfc204f20101c),
    .INIT_01(256'h022bfc09c0c204f4022bfc2b03c204f8022bfc2b80c20518022bfc204f420582),
    .INIT_02(256'h022bfc204cc204f2022bfc09c0c20526022bfc2b02c2052e022bfc204cc2200a),
    .INIT_03(256'h022bfc2b00c20512022bfc204cc20516022bfc09c0c20522022bfc2b01c25000),
    .INIT_04(256'h022bfc2500020522022bfc204f225000022bfc204cc204f4022bfc09c0c20530),
    .INIT_05(256'h022bfc20540204f4022bfc2054020538022bfc2054020522022bfc205402052c),
    .INIT_06(256'h022bfc2054020514022bfc2054020518022bfc2054020534022bfc2054025000),
    .INIT_07(256'h022bfc366242051c022bfc1d00025000022bfc0b032204f4022bfc2500020526),
    .INIT_08(256'h022bfc204f20300f022bfc2053409001022bfc2052e204f4022bfc2051620536),
    .INIT_09(256'h022bfc2051220512022bfc2052825000022bfc20516204f2022bfc25000204cb),
    .INIT_0A(256'h022bfc1d00003008022bfc0b03209002022bfc25000204f4022bfc204f22051c),
    .INIT_0B(256'h022bfc20518204cb022bfc2052c1400e022bfc2051a1400e022bfc366311400e),
    .INIT_0C(256'h022bfc2051601100022bfc2051a010c0022bfc2500025000022bfc204f2204f2),
    .INIT_0D(256'h022bfc2053001d00022bfc2060201e02022bfc204f201f00022bfc20516207c4),
    .INIT_0E(256'h022bfc1410601000022bfc0b11325000022bfc204f4207f2022bfc2051201c00),
    .INIT_0F(256'h022bfc0b00f01e00022bfc1410601f00022bfc14106207c4022bfc1410601103),
    .INIT_10(256'h022bfc204cb25000022bfc0b00e207f2022bfc204cb01c00022bfc0401001d00),
    .INIT_11(256'h022bfc204cb01f00022bfc0b00c207c4022bfc204cb01100022bfc0b00d010c0),
    .INIT_12(256'h022bfc204f4207f2022bfc2051201c00022bfc2052801d01022bfc204f201e00),
    .INIT_13(256'h022bfc14106207c4022bfc0b11301100022bfc204cb010a0022bfc0100025000),
    .INIT_14(256'h022bfc204cb01c00022bfc0401001d00022bfc0b01201e00022bfc1410601f00),
    .INIT_15(256'h022bfc204cb03f81022bfc0b010207e2022bfc204cb25000022bfc0b011207f2),
    .INIT_16(256'h022bfc1dcff05f00022bfc0bc1703c3f022bfc2500003d7c022bfc204f203e3c),
    .INIT_17(256'h022bfc3469e207f2022bfc1dcff05c00022bfc0bc1605d02022bfc3469805e40),
    .INIT_18(256'h022bfc0bc1803e7f022bfc3469803fff022bfc1dcff207e2022bfc0bc1925000),
    .INIT_19(256'h022bfc1dcff05e80022bfc0bc1b05f00022bfc3469e03cff022bfc1dcff03dfd),
    .INIT_1A(256'h022bfc3469e25000022bfc1dcff207f2022bfc0bc1a05c00022bfc3469805d00),
    .INIT_1B(256'h022bfc0bc1c25000022bfc34698207c4022bfc1dcff01101022bfc0bc1d010c0),
    .INIT_1C(256'h022bfc0bd2003dfe022bfc2500003eff022bfc3469e03fff022bfc1dcff207e2),
    .INIT_1D(256'h022bfc20698206b0022bfc0bc1725000022bfc3267c207f2022bfc1dd0003cff),
    .INIT_1E(256'h022bfc206aa20270022bfc0bc2001100022bfc206a401010022bfc0bc162026c),
    .INIT_1F(256'h022bfc0bc1925000022bfc32685207db022bfc1dd0001010022bfc0bd2101100),
    .INIT_20(256'h022bfc0bc2101100022bfc206a401014022bfc0bc182026c022bfc20698207a6),
    .INIT_21(256'h022bfc3268e207db022bfc1dd0001014022bfc0bd2201100022bfc206aa20270),
    .INIT_22(256'h022bfc206a401018022bfc0bc1a2026c022bfc20698207ac022bfc0bc1b25000),
    .INIT_23(256'h022bfc1dd0001018022bfc0bd2301100022bfc206aa20270022bfc0bc2201100),
    .INIT_24(256'h022bfc0bc1c2026c022bfc20698207b6022bfc0bc1d25000022bfc32697207db),
    .INIT_25(256'h022bfc250000101c022bfc206aa20270022bfc0bc2301100022bfc206a40101c),
    .INIT_26(256'h022bfc204cc207e2022bfc204f425000022bfc20518207db022bfc2053e01100),
    .INIT_27(256'h022bfc2053803cff022bfc2051403dfe022bfc2500003eff022bfc204f403fff),
    .INIT_28(256'h022bfc2500005c00022bfc204f205d01022bfc204cc05e00022bfc204f405f00),
    .INIT_29(256'h022bfc204cc2026c022bfc204f4206b0022bfc2053825000022bfc20514207f2),
    .INIT_2A(256'h022bfc2053c01100022bfc205282029b022bfc2500001100022bfc204f401010),
    .INIT_2B(256'h022bfc25000207a6022bfc204f225000022bfc204cc207db022bfc204f401010),
    .INIT_2C(256'h022bfc2b08e2029b022bfc2b1bb01100022bfc2b21a01014022bfc2bec92026c),
    .INIT_2D(256'h022bfc01c0025000022bfc25000207db022bfc2007301014022bfc2083501100),
    .INIT_2E(256'h022bfc206c901100022bfc01c1001018022bfc250002026c022bfc206c9207ac),
    .INIT_2F(256'h022bfc25000207db022bfc206c901018022bfc01c0701100022bfc250002029b),
    .INIT_30(256'h022bfc01c010101c022bfc250002026c022bfc206c9207b6022bfc01c0d25000),
    .INIT_31(256'h022bfc206c901100022bfc01c040101c022bfc250002029b022bfc206c901100),
    .INIT_32(256'h022bfc01f001d001022bfc01e000b01e022bfc01d0025000022bfc25000207db),
    .INIT_33(256'h022bfc207c40b517022bfc011000b416022bfc0108001200022bfc207cd36333),
    .INIT_34(256'h022bfc2b00a04210022bfc2b3892f917022bfc250002f816022bfc206d820849),
    .INIT_35(256'h022bfc250002f818022bfc2083520849022bfc2b08e0b519022bfc2b63b0b418),
    .INIT_36(256'h022bfc2b08e0b51b022bfc2b37b0b41a022bfc2b00a04210022bfc2b2092f919),
    .INIT_37(256'h022bfc2b64904210022bfc206c62f91b022bfc250002f81a022bfc2083520849),
    .INIT_38(256'h022bfc208352f81c022bfc2b08e20849022bfc2b5bb0b51d022bfc2b62a0b41c),
    .INIT_39(256'h022bfc206b0322f5022bfc207660d202022bfc206b004210022bfc250002f91d),
    .INIT_3A(256'h022bfc2b5bb2061d022bfc2b62a20632022bfc2b6492f21e022bfc206c601202),
    .INIT_3B(256'h022bfc206b032378022bfc250001d001022bfc208350b032022bfc2b08e2062a),
    .INIT_3C(256'h022bfc206b005020022bfc2076620551022bfc206b03239e022bfc207661d002),
    .INIT_3D(256'h022bfc2b5bb208ab022bfc2b62a2f21e022bfc2b64901204022bfc206c622374),
    .INIT_3E(256'h022bfc206b02f115022bfc250002f014022bfc208350b117022bfc2b08e0b016),
    .INIT_3F(256'h022bfc206b00b018022bfc2076634496022bfc206b01f1ff022bfc207661d0ff),
    .INIT_40(256'h022bfc2b6491d0ff022bfc206c62f115022bfc206b02f014022bfc207660b119),
    .INIT_41(256'h022bfc208350b11b022bfc2b08e0b01a022bfc2b5bb34496022bfc2b62a1f1ff),
    .INIT_42(256'h022bfc2b10a1f1ff022bfc2b6491d0ff022bfc206c32f115022bfc250002f014),
    .INIT_43(256'h022bfc2b6c92f014022bfc208350b11d022bfc2b08e0b01c022bfc2bdfb34496),
    .INIT_44(256'h022bfc2083534496022bfc2b08e1f1ff022bfc2bebb1d0ff022bfc2b10a2f115),
    .INIT_45(256'h022bfc207e90b013022bfc01ccc36327022bfc206b01d000022bfc250000b032),
    .INIT_46(256'h022bfc2b64932322022bfc206c31d001022bfc206b032320022bfc2075a1d000),
    .INIT_47(256'h022bfc2083532326022bfc2b08e1d003022bfc2bdfb32324022bfc2b10a1d002),
    .INIT_48(256'h022bfc2b08e22327022bfc2bebb20814022bfc2b10a22327022bfc2b6c92080a),
    .INIT_49(256'h022bfc01cd820632022bfc206b02082a022bfc2500022327022bfc208352081f),
    .INIT_4A(256'h022bfc01ccc0b032022bfc206b02062a022bfc2075a2065a022bfc207e92061d),
    .INIT_4B(256'h022bfc206c33239e022bfc206b01d002022bfc2075a32378022bfc207e91d001),
    .INIT_4C(256'h022bfc2b08e1d008022bfc2bdfb22374022bfc2b10a030df022bfc2b64920551),
    .INIT_4D(256'h022bfc2bebb20516022bfc2b10a20534022bfc2b6c920516022bfc2083536340),
    .INIT_4E(256'h022bfc206b01d001022bfc250000b032022bfc2083520602022bfc2b08e204f2),
    .INIT_4F(256'h022bfc206b022374022bfc2075a05020022bfc207e920551022bfc01ce432378),
    .INIT_50(256'h022bfc206b02053a022bfc2075a20512022bfc207e93634d022bfc01cd81d010),
    .INIT_51(256'h022bfc206b00b032022bfc2075a20602022bfc207e9204f2022bfc01ccc20540),
    .INIT_52(256'h022bfc2bdfb05020022bfc2b10a20551022bfc2b64932378022bfc206c31d001),
    .INIT_53(256'h022bfc2b10a20512022bfc2b6c93635a022bfc208351d020022bfc2b08e22374),
    .INIT_54(256'h022bfc2500020602022bfc20835204f2022bfc2b08e20540022bfc2bebb2053a),
    .INIT_55(256'h022bfc2b08e20551022bfc2b47b32378022bfc2b22a1d001022bfc2b1c90b032),
    .INIT_56(256'h022bfc2b22a36367022bfc2b4891d040022bfc2500022374022bfc20835030df),
    .INIT_57(256'h022bfc25000204f2022bfc2083520540022bfc2b08e2053a022bfc2b57b20512),
    .INIT_58(256'h022bfc2b08e32378022bfc2b6bb1d001022bfc2b66a0b032022bfc2b5c920602),
    .INIT_59(256'h022bfc2b66a1d080022bfc2b6c922374022bfc25000030df022bfc2083520551),
    .INIT_5A(256'h022bfc250002052a022bfc208352052e022bfc2b08e20534022bfc2b7bb3602a),
    .INIT_5B(256'h022bfc010801d001022bfc206b00b032022bfc2076620602022bfc206b0204f2),
    .INIT_5C(256'h022bfc2500022374022bfc206d2030df022bfc207c420551022bfc0110132378),
    .INIT_5D(256'h022bfc2075a2200a022bfc207e920566022bfc01c0e01008022bfc206b02055a),
    .INIT_5E(256'h022bfc206b01d002022bfc250000b002022bfc206b720280022bfc206b020277),
    .INIT_5F(256'h022bfc206b01d003022bfc2075a0b002022bfc207e920289022bfc01c1e32382),
    .INIT_60(256'h022bfc2075a01060022bfc207e92076c022bfc01c0e20292022bfc206b732382),
    .INIT_61(256'h022bfc206b02d003022bfc250002f032022bfc206b701000022bfc206b02055a),
    .INIT_62(256'h022bfc206b02b04f022bfc2075a2b08f022bfc207e92b20f022bfc01c2e2b40f),
    .INIT_63(256'h022bfc2075a2d010022bfc207e901020022bfc01c1e2d010022bfc206b701040),
    .INIT_64(256'h022bfc207e92d010022bfc01c0e01004022bfc206b72d010022bfc206b001008),
    .INIT_65(256'h022bfc250002d010022bfc206b701080022bfc206b02b10f022bfc2075a2b80f),
    .INIT_66(256'h022bfc1d00320566022bfc3279f01000022bfc1d0022d010022bfc0b00201010),
    .INIT_67(256'h022bfc207742d003022bfc327a301002022bfc1d0042200a022bfc327a120594),
    .INIT_68(256'h022bfc2078736412022bfc227a41d004022bfc2077b0b01e022bfc227a42200a),
    .INIT_69(256'h022bfc01c0e2045f022bfc206b0323f6022bfc250000d004022bfc0b00209002),
    .INIT_6A(256'h022bfc25000011b3022bfc206b001e40022bfc2075a01f0a022bfc207e920485),
    .INIT_6B(256'h022bfc2075a2df0a022bfc207e909d07022bfc01c1a2043f022bfc206b00120b),
    .INIT_6C(256'h022bfc2075a363b7022bfc207e91ce10022bfc01c0e2dd08022bfc206b02de09),
    .INIT_6D(256'h022bfc01c2611e01022bfc206b0223ba022bfc25000363b7022bfc206b01cf20),
    .INIT_6E(256'h022bfc01c1a0b117022bfc206b00b016022bfc2075a223ad022bfc207e913f00),
    .INIT_6F(256'h022bfc01c0e1f1ff022bfc206b01d0ff022bfc2075a2f115022bfc207e92f014),
    .INIT_70(256'h022bfc250000d0ff022bfc206b001200022bfc2075a20447022bfc207e9323c6),
    .INIT_71(256'h022bfc2d1080b119022bfc2d0080b018022bfc2b4192f220022bfc2b00a14200),
    .INIT_72(256'h022bfc2d1081f1ff022bfc2d0081d0ff022bfc2b2592f115022bfc2b00a2f014),
    .INIT_73(256'h022bfc2dc080d0ff022bfc2b28901200022bfc2b00a20447022bfc25000323d2),
    .INIT_74(256'h022bfc250000b11b022bfc2df080b01a022bfc2de082f221022bfc2dd0814200),
    .INIT_75(256'h022bfc09d081f1ff022bfc09c081d0ff022bfc2b2892f115022bfc2b00a2f014),
    .INIT_76(256'h022bfc2d10a0d0ff022bfc2500001200022bfc09f0820447022bfc09e08323de),
    .INIT_77(256'h022bfc2de080b11d022bfc2dd080b01c022bfc2dc082f222022bfc2d00914200),
    .INIT_78(256'h022bfc2d0091d0ff022bfc2d10a2f115022bfc250002f014022bfc2df0801200),
    .INIT_79(256'h022bfc09f0801200022bfc09e0820447022bfc09d08323eb022bfc09c081f1ff),
    .INIT_7A(256'h022bfc2d10a20625022bfc011022f223022bfc0105014200022bfc250000d0ff),
    .INIT_7B(256'h022bfc206d20b121022bfc250000b020022bfc2dc082062a022bfc2d00920673),
    .INIT_7C(256'h022bfc206d80b123022bfc207cd04010022bfc250000b122022bfc207d404010),
    .INIT_7D(256'h022bfc2500005040022bfc2080120551022bfc206b0323f9022bfc2500004010),
    .INIT_7E(256'h022bfc207ac2055a022bfc25000030bf022bfc2080120551022bfc207a6223fb),
    .INIT_7F(256'h022bfc208011900102d003207b60b01f0010ff250002f03b02bff0208010b00e),
    .INITP_00(256'hd6d16a71de5f5455ded5dedaf7cede56de5b5ac8dddc43c25add7ac47268e0c5),
    .INITP_01(256'he8e673f0fbc7c2ec657ed066e3e87c46f87d7bd5c672f7427976657359fc7a69),
    .INITP_02(256'h5cd9e0dcda71f64cca67c8f4d579ede673c9cd79c2ece5ddd6f1c6e4c86ad579),
    .INITP_03(256'he1517bd0c8e958e9dafb5afc477fd952e7dbdd79d7dbe9d45bf0dad5745e52e1),
    .INITP_04(256'he5f57f475749726177c868d9efd4fd547c4bc8725f68df7a4dfd51c8f3def35d),
    .INITP_05(256'hf97ae970f96974fa7af95f5d63c5e7fcf3ced0c3fa7a72c35d41e8fdf5c9d2c3),
    .INITP_06(256'hf2e5e04b60ed5363654be5cf53e6616bc15ad659ea5659f9f96d70f96b74f1e1),
    .INITP_07(256'hdb64d9fed77552e07ecafb6f4dec51785f6bd0e0e24ef57fdc60d26dcc77e2cd),
    .INITP_08(256'hdafd65e37fe6dafd4166c4ff5ee6d875dbd062647be77675d361e3c6e770596c),
    .INITP_09(256'hc8744e7547ff51e741f3dcccfcf16bf5f04166dc7bdfeec77bcf60ca73d7eec7),
    .INITP_0A(256'hf4dc6a65ff48e4caeac17df37edbe04a7a464df774777fe6d36b437755e15667),
    .INITP_0B(256'hc2e9cbf741fc49d0fecd64d4e4ecca4fccd36bd8f0596ed5f64ae5d6607e6d57),
    .INITP_0C(256'h7fe95af3566cd6eae04248ed57e55154f54262c54ef0d0e543fcced4eb41e8c4),
    .INITP_0D(256'he9c7eec2e3df7bd0644be7c1f25461d1e34eef5cfb48f5cbecd778f37b4be4ce),
    .INITP_0E(256'hefe6cfccf2714863675ad1d8fc416df6495bd3f7615c4cd8ed4069ccfd5d6b4f),
    .INITP_0F(256'h4dd61470e8644bf9e04b50f0f7447b5d74f347587b455bfd476be24446f47542),
